magic
tech sky130B
magscale 1 2
timestamp 1666464484
<< nwell >>
rect 2372 -270 14193 34
<< pwell >>
rect 699 -220 2257 4351
<< obsli1 >>
rect 122 0 14571 39532
rect 122 -194 2231 0
rect 2407 -23 2609 0
rect 13946 -23 14136 0
rect 2407 -213 14136 -23
<< obsm1 >>
rect 37 0 14583 39538
rect 725 -181 1771 0
rect 2407 -23 2670 0
tri 2670 -23 2693 0 sw
tri 13885 -23 13908 0 se
rect 13908 -23 14136 0
rect 2407 -213 14136 -23
<< metal2 >>
rect 99 -407 4879 4
rect 10078 -407 14858 4725
<< obsm2 >>
rect 53 4781 14858 38608
rect 53 60 10022 4781
rect 4935 0 10022 60
rect 5179 -407 5579 -23
<< metal3 >>
rect 99 -407 4879 2985
rect 5179 -407 7379 138
rect 7578 -407 9778 1859
rect 10078 -407 14858 2985
<< obsm3 >>
rect 48 3065 14858 39593
rect 4959 1939 9998 3065
rect 4959 218 7498 1939
rect 4959 138 5099 218
rect 7459 138 7498 218
rect 9858 138 9998 1939
<< metal4 >>
rect 0 39593 241 39993
rect 14845 39593 15000 39993
rect 0 34750 254 39593
rect 14746 34750 15000 39593
rect 0 13600 254 18593
rect 14746 13600 15000 18593
rect 0 12410 254 13300
rect 14746 12410 15000 13300
rect 0 11240 254 12130
rect 14746 11240 15000 12130
rect 0 10814 15000 11214
rect 0 10218 254 10814
rect 14746 10218 15000 10814
rect 0 9922 254 10158
rect 14746 9922 15000 10158
rect 0 9266 15000 9922
rect 0 9140 254 9206
rect 14746 9140 15000 9206
rect 0 7910 254 8840
rect 14746 7910 15000 8840
rect 0 6940 254 7630
rect 14746 6940 15000 7630
rect 0 5970 254 6660
rect 14746 5970 15000 6660
rect 0 4760 254 5690
rect 14746 4760 15000 5690
rect 0 3550 254 4480
rect 14746 3550 15000 4480
rect 0 2580 193 3270
rect 14807 2580 15000 3270
rect 0 1370 254 2300
rect 14746 1370 15000 2300
rect 0 0 254 1090
rect 14746 0 15000 1090
<< obsm4 >>
rect 241 39593 14845 39993
rect 334 34670 14666 39593
rect 0 18629 15000 34670
rect 0 18593 143 18629
rect 0 13520 143 13600
rect 334 13520 14666 18629
rect 0 13300 15000 13520
rect 0 12330 143 12410
rect 334 12330 14666 13300
rect 0 12130 15000 12330
rect 334 11294 14666 12130
rect 334 10218 14666 10734
rect 0 10158 15000 10218
rect 334 10002 14666 10158
rect 0 9206 15000 9240
rect 0 9060 143 9140
rect 334 9060 14666 9186
rect 0 8840 15000 9060
rect 0 7830 143 7910
rect 334 7830 14666 8840
rect 0 7630 15000 7830
rect 0 6860 143 6940
rect 334 6860 14666 7630
rect 0 6660 15000 6860
rect 0 5890 143 5970
rect 334 5890 14666 6660
rect 0 5690 15000 5890
rect 0 4680 143 4760
rect 334 4680 14666 5690
rect 0 4480 15000 4680
rect 0 3513 105 3550
rect 0 3489 143 3513
rect 0 3470 105 3489
rect 334 3470 14666 4480
rect 0 3350 15000 3470
rect 0 3337 105 3350
rect 273 3337 14727 3350
rect 0 3313 15000 3337
rect 0 3270 105 3313
rect 0 2500 143 2580
rect 273 2500 14727 3313
rect 0 2300 15000 2500
rect 0 1290 143 1370
rect 334 1290 14666 2300
rect 0 1090 15000 1290
rect 334 0 14666 1090
<< metal5 >>
rect 1410 20617 13578 32782
rect 0 13600 254 18590
rect 14746 13600 15000 18590
rect 0 12430 254 13280
rect 14746 12430 15000 13280
rect 0 11260 254 12110
rect 14746 11260 15000 12110
rect 0 9140 254 10940
rect 14746 9140 15000 10940
rect 0 7930 254 8820
rect 14746 7930 15000 8820
rect 0 6961 254 7610
rect 14746 6961 15000 7610
rect 0 5990 254 6640
rect 14746 5990 15000 6640
rect 0 4780 254 5670
rect 14746 4780 15000 5670
rect 0 3570 254 4460
rect 14746 3570 15000 4460
rect 0 2600 193 3250
rect 14807 2600 15000 3250
rect 0 1390 254 2280
rect 14746 1390 15000 2280
rect 0 20 254 1070
rect 14746 20 15000 1070
<< obsm5 >>
rect 0 33102 15000 39993
rect 0 20297 1090 33102
rect 13898 20297 15000 33102
rect 0 18910 15000 20297
rect 0 18729 143 18910
rect 574 18729 14426 18910
rect 0 18629 15000 18729
rect 0 18590 143 18629
rect 0 13420 143 13600
rect 574 13420 14426 18629
rect 0 13280 15000 13420
rect 0 12250 143 12430
rect 574 12250 14426 13280
rect 0 12110 15000 12250
rect 574 11260 14426 12110
rect 0 10940 15000 11260
rect 0 8960 143 9140
rect 574 8960 14426 10940
rect 0 8820 15000 8960
rect 0 7750 143 7930
rect 574 7750 14426 8820
rect 0 7620 15000 7750
rect 0 7610 143 7620
rect 0 6780 143 6961
rect 574 6780 14426 7620
rect 0 6650 15000 6780
rect 0 6640 143 6650
rect 0 5810 143 5990
rect 574 5810 14426 6650
rect 0 5670 15000 5810
rect 0 4600 143 4780
rect 574 4600 14426 5670
rect 0 4460 15000 4600
rect 0 3390 143 3570
rect 574 3390 14426 4460
rect 0 3260 15000 3390
rect 0 3250 143 3260
rect 574 3250 14426 3260
rect 513 2600 14487 3250
rect 0 2420 143 2600
rect 574 2420 14426 2600
rect 0 2280 15000 2420
rect 0 1209 143 1390
rect 574 1209 14426 2280
rect 0 1070 15000 1209
rect 574 20 14426 1070
<< labels >>
rlabel metal4 s 14746 10218 15000 10814 6 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel metal4 s 0 10218 254 10814 6 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel metal4 s 0 9266 15000 9922 6 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel metal4 s 0 9266 254 9862 6 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel metal2 s 10078 -407 14858 4725 6 DRN_HVC
port 3 nsew power bidirectional
rlabel metal3 s 7578 -407 9778 1859 6 DRN_HVC
port 3 nsew power bidirectional
rlabel metal2 s 99 -407 4879 4 8 SRC_BDY_HVC
port 4 nsew ground bidirectional
rlabel metal3 s 5179 -407 7379 138 8 SRC_BDY_HVC
port 4 nsew ground bidirectional
rlabel metal5 s 1410 20617 13578 32782 6 VDDA_PAD
port 5 nsew power bidirectional
rlabel metal5 s 14746 9140 15000 10940 6 VSSA
port 6 nsew ground bidirectional
rlabel metal5 s 14746 6961 15000 7610 6 VSSA
port 6 nsew ground bidirectional
rlabel metal5 s 0 9140 254 10940 6 VSSA
port 6 nsew ground bidirectional
rlabel metal5 s 0 6961 254 7610 6 VSSA
port 6 nsew ground bidirectional
rlabel metal4 s 14746 9922 15000 10158 6 VSSA
port 6 nsew ground bidirectional
rlabel metal4 s 0 10814 15000 11214 6 VSSA
port 6 nsew ground bidirectional
rlabel metal4 s 14746 9140 15000 9206 6 VSSA
port 6 nsew ground bidirectional
rlabel metal4 s 14746 6940 15000 7630 6 VSSA
port 6 nsew ground bidirectional
rlabel metal4 s 0 9140 254 9206 6 VSSA
port 6 nsew ground bidirectional
rlabel metal4 s 0 9922 254 10158 6 VSSA
port 6 nsew ground bidirectional
rlabel metal4 s 0 10874 254 10940 6 VSSA
port 6 nsew ground bidirectional
rlabel metal4 s 0 6940 254 7630 6 VSSA
port 6 nsew ground bidirectional
rlabel metal3 s 10078 -407 14858 2985 6 VDDA
port 7 nsew power bidirectional
rlabel metal3 s 99 -407 4879 2985 6 VDDA
port 7 nsew power bidirectional
rlabel metal5 s 14807 2600 15000 3250 6 VDDA
port 7 nsew power bidirectional
rlabel metal5 s 0 2600 193 3250 6 VDDA
port 7 nsew power bidirectional
rlabel metal4 s 14807 2580 15000 3270 6 VDDA
port 7 nsew power bidirectional
rlabel metal4 s 0 2580 193 3270 6 VDDA
port 7 nsew power bidirectional
rlabel metal5 s 14746 5990 15000 6640 6 VSWITCH
port 8 nsew power bidirectional
rlabel metal5 s 0 5990 254 6640 6 VSWITCH
port 8 nsew power bidirectional
rlabel metal4 s 14746 5970 15000 6660 6 VSWITCH
port 8 nsew power bidirectional
rlabel metal4 s 0 5970 254 6660 6 VSWITCH
port 8 nsew power bidirectional
rlabel metal5 s 14746 12430 15000 13280 6 VDDIO_Q
port 9 nsew power bidirectional
rlabel metal5 s 0 12430 254 13280 6 VDDIO_Q
port 9 nsew power bidirectional
rlabel metal4 s 14746 12410 15000 13300 6 VDDIO_Q
port 9 nsew power bidirectional
rlabel metal4 s 0 12410 254 13300 6 VDDIO_Q
port 9 nsew power bidirectional
rlabel metal5 s 14746 20 15000 1070 6 VCCHIB
port 10 nsew power bidirectional
rlabel metal5 s 0 20 254 1070 6 VCCHIB
port 10 nsew power bidirectional
rlabel metal4 s 14746 0 15000 1090 6 VCCHIB
port 10 nsew power bidirectional
rlabel metal4 s 0 0 254 1090 6 VCCHIB
port 10 nsew power bidirectional
rlabel metal5 s 14746 13600 15000 18590 6 VDDIO
port 11 nsew power bidirectional
rlabel metal5 s 14746 3570 15000 4460 6 VDDIO
port 11 nsew power bidirectional
rlabel metal5 s 0 13600 254 18590 6 VDDIO
port 11 nsew power bidirectional
rlabel metal5 s 0 3570 254 4460 6 VDDIO
port 11 nsew power bidirectional
rlabel metal4 s 14746 3550 15000 4480 6 VDDIO
port 11 nsew power bidirectional
rlabel metal4 s 14746 13600 15000 18593 6 VDDIO
port 11 nsew power bidirectional
rlabel metal4 s 0 3550 254 4480 6 VDDIO
port 11 nsew power bidirectional
rlabel metal4 s 0 13600 254 18593 6 VDDIO
port 11 nsew power bidirectional
rlabel metal5 s 14746 1390 15000 2280 6 VCCD
port 12 nsew power bidirectional
rlabel metal5 s 0 1390 254 2280 6 VCCD
port 12 nsew power bidirectional
rlabel metal4 s 14746 1370 15000 2300 6 VCCD
port 12 nsew power bidirectional
rlabel metal4 s 0 1370 254 2300 6 VCCD
port 12 nsew power bidirectional
rlabel metal4 s 14845 34750 15000 39993 6 VSSIO
port 13 nsew ground bidirectional
rlabel metal4 s 0 34750 241 39993 6 VSSIO
port 13 nsew ground bidirectional
rlabel metal4 s 126 37913 128 37915 6 VSSIO
port 13 nsew ground bidirectional
rlabel metal4 s 14872 37913 14874 37915 6 VSSIO
port 13 nsew ground bidirectional
rlabel metal5 s 14746 4780 15000 5670 6 VSSIO
port 13 nsew ground bidirectional
rlabel metal5 s 0 4780 254 5670 6 VSSIO
port 13 nsew ground bidirectional
rlabel metal4 s 14746 4760 15000 5690 6 VSSIO
port 13 nsew ground bidirectional
rlabel metal4 s 14746 34750 15000 39593 6 VSSIO
port 13 nsew ground bidirectional
rlabel metal4 s 0 34750 254 39593 6 VSSIO
port 13 nsew ground bidirectional
rlabel metal4 s 0 4760 254 5690 6 VSSIO
port 13 nsew ground bidirectional
rlabel metal5 s 14746 7930 15000 8820 6 VSSD
port 14 nsew ground bidirectional
rlabel metal5 s 0 7930 254 8820 6 VSSD
port 14 nsew ground bidirectional
rlabel metal4 s 14746 7910 15000 8840 6 VSSD
port 14 nsew ground bidirectional
rlabel metal4 s 0 7910 254 8840 6 VSSD
port 14 nsew ground bidirectional
rlabel metal5 s 14746 11260 15000 12110 6 VSSIO_Q
port 15 nsew ground bidirectional
rlabel metal5 s 0 11260 254 12110 6 VSSIO_Q
port 15 nsew ground bidirectional
rlabel metal4 s 14746 11240 15000 12130 6 VSSIO_Q
port 15 nsew ground bidirectional
rlabel metal4 s 0 11240 254 12130 6 VSSIO_Q
port 15 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 15000 39593
string LEFclass PAD POWER
string LEFview TRUE
string GDS_END 2458880
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io.gds
string GDS_START 2445208
<< end >>
