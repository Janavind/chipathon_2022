magic
tech sky130A
timestamp 1666199351
<< properties >>
string GDS_END 3228654
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 3225706
<< end >>
