magic
tech sky130A
magscale 1 2
timestamp 1666199351
<< nwell >>
rect -36 679 8508 1471
<< locali >>
rect 0 1397 8472 1431
rect 64 636 98 702
rect 196 652 449 686
rect 547 653 817 687
rect 919 674 1293 708
rect 1609 690 2093 724
rect 2860 690 3865 724
rect 6125 690 6159 724
rect 919 670 953 674
rect 0 -17 8472 17
use sky130_sram_2kbyte_1rw1r_32x512_8_pinv_0  sky130_sram_2kbyte_1rw1r_32x512_8_pinv_0_0
timestamp 1666199351
transform 1 0 368 0 1 0
box -36 -17 404 1471
use sky130_sram_2kbyte_1rw1r_32x512_8_pinv_0  sky130_sram_2kbyte_1rw1r_32x512_8_pinv_0_1
timestamp 1666199351
transform 1 0 0 0 1 0
box -36 -17 404 1471
use sky130_sram_2kbyte_1rw1r_32x512_8_pinv_7  sky130_sram_2kbyte_1rw1r_32x512_8_pinv_7_0
timestamp 1666199351
transform 1 0 736 0 1 0
box -36 -17 512 1471
use sky130_sram_2kbyte_1rw1r_32x512_8_pinv_18  sky130_sram_2kbyte_1rw1r_32x512_8_pinv_18_0
timestamp 1666199351
transform 1 0 1212 0 1 0
box -36 -17 836 1471
use sky130_sram_2kbyte_1rw1r_32x512_8_pinv_19  sky130_sram_2kbyte_1rw1r_32x512_8_pinv_19_0
timestamp 1666199351
transform 1 0 2012 0 1 0
box -36 -17 1808 1471
use sky130_sram_2kbyte_1rw1r_32x512_8_pinv_20  sky130_sram_2kbyte_1rw1r_32x512_8_pinv_20_0
timestamp 1666199351
transform 1 0 3784 0 1 0
box -36 -17 4724 1471
<< labels >>
rlabel locali s 6142 707 6142 707 4 Z
port 1 nsew
rlabel locali s 81 669 81 669 4 A
port 2 nsew
rlabel locali s 4236 0 4236 0 4 gnd
port 3 nsew
rlabel locali s 4236 1414 4236 1414 4 vdd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 8472 1414
string GDS_END 10923926
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_2kbyte_1rw1r_32x512_8.gds
string GDS_START 10922036
<< end >>
