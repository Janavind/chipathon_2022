magic
tech sky130B
magscale 1 2
timestamp 1666464484
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 1 21 827 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 289 47 319 177
rect 387 47 417 177
rect 491 47 521 177
rect 603 47 633 177
rect 719 47 749 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 289 297 319 497
rect 387 297 417 497
rect 491 297 521 497
rect 605 297 635 497
rect 719 297 749 497
<< ndiff >>
rect 27 161 79 177
rect 27 127 35 161
rect 69 127 79 161
rect 27 93 79 127
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 161 163 177
rect 109 127 119 161
rect 153 127 163 161
rect 109 93 163 127
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 93 289 177
rect 193 59 219 93
rect 253 59 289 93
rect 193 47 289 59
rect 319 47 387 177
rect 417 47 491 177
rect 521 131 603 177
rect 521 97 558 131
rect 592 97 603 131
rect 521 47 603 97
rect 633 97 719 177
rect 633 63 660 97
rect 694 63 719 97
rect 633 47 719 63
rect 749 101 801 177
rect 749 67 759 101
rect 793 67 801 101
rect 749 47 801 67
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 349 79 383
rect 27 315 35 349
rect 69 315 79 349
rect 27 297 79 315
rect 109 485 163 497
rect 109 451 119 485
rect 153 451 163 485
rect 109 417 163 451
rect 109 383 119 417
rect 153 383 163 417
rect 109 349 163 383
rect 109 315 119 349
rect 153 315 163 349
rect 109 297 163 315
rect 193 485 289 497
rect 193 451 232 485
rect 266 451 289 485
rect 193 417 289 451
rect 193 383 232 417
rect 266 383 289 417
rect 193 297 289 383
rect 319 477 387 497
rect 319 443 334 477
rect 368 443 387 477
rect 319 401 387 443
rect 319 367 334 401
rect 368 367 387 401
rect 319 297 387 367
rect 417 485 491 497
rect 417 451 441 485
rect 475 451 491 485
rect 417 297 491 451
rect 521 477 605 497
rect 521 443 555 477
rect 589 443 605 477
rect 521 401 605 443
rect 521 367 555 401
rect 589 367 605 401
rect 521 297 605 367
rect 635 297 719 497
rect 749 477 801 497
rect 749 443 759 477
rect 793 443 801 477
rect 749 409 801 443
rect 749 375 759 409
rect 793 375 801 409
rect 749 297 801 375
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 119 127 153 161
rect 119 59 153 93
rect 219 59 253 93
rect 558 97 592 131
rect 660 63 694 97
rect 759 67 793 101
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 119 451 153 485
rect 119 383 153 417
rect 119 315 153 349
rect 232 451 266 485
rect 232 383 266 417
rect 334 443 368 477
rect 334 367 368 401
rect 441 451 475 485
rect 555 443 589 477
rect 555 367 589 401
rect 759 443 793 477
rect 759 375 793 409
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 289 497 319 523
rect 387 497 417 523
rect 491 497 521 523
rect 605 497 635 523
rect 719 497 749 523
rect 79 265 109 297
rect 163 265 193 297
rect 289 265 319 297
rect 387 265 417 297
rect 491 265 521 297
rect 605 265 635 297
rect 719 265 749 297
rect 79 249 247 265
rect 79 215 203 249
rect 237 215 247 249
rect 79 199 247 215
rect 289 249 343 265
rect 289 215 299 249
rect 333 215 343 249
rect 289 199 343 215
rect 387 249 441 265
rect 387 215 397 249
rect 431 215 441 249
rect 387 199 441 215
rect 491 249 545 265
rect 491 215 501 249
rect 535 215 545 249
rect 491 199 545 215
rect 603 249 657 265
rect 603 215 613 249
rect 647 215 657 249
rect 603 199 657 215
rect 719 249 783 265
rect 719 215 739 249
rect 773 215 783 249
rect 719 199 783 215
rect 79 177 109 199
rect 163 177 193 199
rect 289 177 319 199
rect 387 177 417 199
rect 491 177 521 199
rect 603 177 633 199
rect 719 177 749 199
rect 79 21 109 47
rect 163 21 193 47
rect 289 21 319 47
rect 387 21 417 47
rect 491 21 521 47
rect 603 21 633 47
rect 719 21 749 47
<< polycont >>
rect 203 215 237 249
rect 299 215 333 249
rect 397 215 431 249
rect 501 215 535 249
rect 613 215 647 249
rect 739 215 773 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 18 485 69 527
rect 232 485 276 527
rect 18 451 35 485
rect 18 417 69 451
rect 18 383 35 417
rect 18 349 69 383
rect 18 315 35 349
rect 18 299 69 315
rect 103 451 119 485
rect 153 451 169 485
rect 103 417 169 451
rect 103 383 119 417
rect 153 383 169 417
rect 103 349 169 383
rect 266 451 276 485
rect 232 417 276 451
rect 266 383 276 417
rect 232 367 276 383
rect 318 477 368 493
rect 318 443 334 477
rect 425 485 491 527
rect 425 451 441 485
rect 475 451 491 485
rect 543 477 605 493
rect 318 401 368 443
rect 543 443 555 477
rect 589 443 605 477
rect 543 401 605 443
rect 318 367 334 401
rect 368 367 555 401
rect 589 367 605 401
rect 759 477 793 493
rect 759 409 793 443
rect 103 315 119 349
rect 153 315 169 349
rect 759 333 793 375
rect 18 161 69 177
rect 18 127 35 161
rect 18 93 69 127
rect 18 59 35 93
rect 103 161 169 315
rect 103 127 119 161
rect 153 127 169 161
rect 203 299 793 333
rect 203 249 237 299
rect 203 165 237 215
rect 299 249 342 265
rect 333 215 342 249
rect 299 199 342 215
rect 379 249 433 265
rect 379 215 397 249
rect 431 215 433 249
rect 203 131 339 165
rect 103 93 169 127
rect 103 59 119 93
rect 153 59 169 93
rect 203 59 219 93
rect 253 59 269 93
rect 18 17 69 59
rect 203 17 269 59
rect 305 85 339 131
rect 379 121 433 215
rect 488 249 535 265
rect 488 215 501 249
rect 488 199 535 215
rect 579 249 647 265
rect 579 215 613 249
rect 579 199 647 215
rect 739 249 801 265
rect 773 215 801 249
rect 739 199 801 215
rect 488 121 524 199
rect 558 131 793 165
rect 759 101 793 131
rect 558 85 592 97
rect 305 51 592 85
rect 644 63 660 97
rect 694 63 710 97
rect 644 17 710 63
rect 759 51 793 67
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
flabel locali s 122 425 156 459 0 FreeSans 200 0 0 0 X
port 10 nsew signal output
flabel locali s 764 221 798 255 0 FreeSans 200 0 0 0 C1
port 5 nsew signal input
flabel locali s 582 221 616 255 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 490 221 524 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 398 221 432 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 306 221 340 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 122 85 156 119 0 FreeSans 200 0 0 0 X
port 10 nsew signal output
flabel locali s 122 153 156 187 0 FreeSans 200 0 0 0 X
port 10 nsew signal output
flabel locali s 122 221 156 255 0 FreeSans 200 0 0 0 X
port 10 nsew signal output
flabel locali s 122 289 156 323 0 FreeSans 200 0 0 0 X
port 10 nsew signal output
flabel locali s 122 357 156 391 0 FreeSans 200 0 0 0 X
port 10 nsew signal output
rlabel comment s 0 0 0 0 4 a311o_2
rlabel metal1 s 0 -48 828 48 1 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 828 592 1 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 828 544
string GDS_END 3708814
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3701494
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 20.700 0.000 
<< end >>
