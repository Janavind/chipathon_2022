magic
tech sky130B
magscale 1 2
timestamp 1666199351
<< locali >>
rect 12028 18138 12590 18733
rect 1835 1730 2397 2325
rect 1835 -41064 2397 -40469
<< obsli1 >>
rect 20504 20659 21046 20675
rect 20504 20625 20506 20659
rect 20540 20625 20578 20659
rect 20612 20625 20650 20659
rect 20684 20625 20722 20659
rect 20756 20625 20794 20659
rect 20828 20625 20866 20659
rect 20900 20625 20938 20659
rect 20972 20625 21010 20659
rect 21044 20625 21046 20659
rect 20504 20609 21046 20625
rect 20414 20547 20448 20563
rect 20414 20475 20448 20513
rect 20414 20403 20448 20441
rect 20414 20331 20448 20369
rect 20414 20259 20448 20297
rect 20414 20187 20448 20225
rect 13851 20143 13985 20159
rect 13851 20109 13865 20143
rect 13899 20109 13937 20143
rect 13971 20109 13985 20143
rect 13851 20093 13985 20109
rect 20414 20115 20448 20153
rect 13815 20043 13849 20059
rect 13815 19993 13849 20009
rect 13901 19993 13935 20059
rect 13987 20043 14021 20059
rect 13987 19993 14021 20009
rect 20414 20043 20448 20081
rect 20414 19993 20448 20009
rect 20500 19993 20534 20563
rect 20586 20547 20620 20563
rect 20586 20475 20620 20513
rect 20586 20403 20620 20441
rect 20586 20331 20620 20369
rect 20586 20259 20620 20297
rect 20586 20187 20620 20225
rect 20586 20115 20620 20153
rect 20586 20043 20620 20081
rect 20586 19993 20620 20009
rect 20672 19993 20706 20563
rect 20758 20547 20792 20563
rect 20758 20475 20792 20513
rect 20758 20403 20792 20441
rect 20758 20331 20792 20369
rect 20758 20259 20792 20297
rect 20758 20187 20792 20225
rect 20758 20115 20792 20153
rect 20758 20043 20792 20081
rect 20758 19993 20792 20009
rect 20844 19993 20878 20563
rect 20930 20547 20964 20563
rect 20930 20475 20964 20513
rect 20930 20403 20964 20441
rect 20930 20331 20964 20369
rect 20930 20259 20964 20297
rect 20930 20187 20964 20225
rect 20930 20115 20964 20153
rect 20930 20043 20964 20081
rect 20930 19993 20964 20009
rect 21016 19993 21050 20563
rect 21102 20547 21136 20563
rect 21102 20475 21136 20513
rect 21102 20403 21136 20441
rect 21102 20331 21136 20369
rect 21102 20259 21136 20297
rect 21102 20187 21136 20225
rect 21102 20115 21136 20153
rect 21102 20043 21136 20081
rect 21102 19993 21136 20009
rect 20591 -24383 20725 -24367
rect 20591 -24417 20605 -24383
rect 20639 -24417 20677 -24383
rect 20711 -24417 20725 -24383
rect 20591 -24435 20725 -24417
rect 20555 -24497 20589 -24481
rect 20555 -24569 20589 -24531
rect 20555 -24641 20589 -24603
rect 20555 -24713 20589 -24675
rect 20555 -24785 20589 -24747
rect 13653 -24815 13787 -24799
rect 13653 -24849 13667 -24815
rect 13701 -24849 13739 -24815
rect 13773 -24849 13787 -24815
rect 13653 -24867 13787 -24849
rect 20555 -24857 20589 -24819
rect 13617 -24929 13651 -24913
rect 13617 -25001 13651 -24963
rect 13617 -25051 13651 -25035
rect 13703 -25051 13737 -24913
rect 13789 -24929 13823 -24913
rect 13789 -25001 13823 -24963
rect 13789 -25051 13823 -25035
rect 20555 -24929 20589 -24891
rect 20555 -25001 20589 -24963
rect 20555 -25055 20589 -25035
rect 20641 -25051 20675 -24481
rect 20727 -24497 20761 -24481
rect 20727 -24569 20761 -24531
rect 20727 -24641 20761 -24603
rect 20727 -24713 20761 -24675
rect 20727 -24785 20761 -24747
rect 20727 -24857 20761 -24819
rect 20727 -24929 20761 -24891
rect 20727 -25001 20761 -24963
rect 20727 -25051 20761 -25035
<< obsli1c >>
rect 20506 20625 20540 20659
rect 20578 20625 20612 20659
rect 20650 20625 20684 20659
rect 20722 20625 20756 20659
rect 20794 20625 20828 20659
rect 20866 20625 20900 20659
rect 20938 20625 20972 20659
rect 21010 20625 21044 20659
rect 20414 20513 20448 20547
rect 20414 20441 20448 20475
rect 20414 20369 20448 20403
rect 20414 20297 20448 20331
rect 20414 20225 20448 20259
rect 13865 20109 13899 20143
rect 13937 20109 13971 20143
rect 20414 20153 20448 20187
rect 20414 20081 20448 20115
rect 13815 20009 13849 20043
rect 13987 20009 14021 20043
rect 20414 20009 20448 20043
rect 20586 20513 20620 20547
rect 20586 20441 20620 20475
rect 20586 20369 20620 20403
rect 20586 20297 20620 20331
rect 20586 20225 20620 20259
rect 20586 20153 20620 20187
rect 20586 20081 20620 20115
rect 20586 20009 20620 20043
rect 20758 20513 20792 20547
rect 20758 20441 20792 20475
rect 20758 20369 20792 20403
rect 20758 20297 20792 20331
rect 20758 20225 20792 20259
rect 20758 20153 20792 20187
rect 20758 20081 20792 20115
rect 20758 20009 20792 20043
rect 20930 20513 20964 20547
rect 20930 20441 20964 20475
rect 20930 20369 20964 20403
rect 20930 20297 20964 20331
rect 20930 20225 20964 20259
rect 20930 20153 20964 20187
rect 20930 20081 20964 20115
rect 20930 20009 20964 20043
rect 21102 20513 21136 20547
rect 21102 20441 21136 20475
rect 21102 20369 21136 20403
rect 21102 20297 21136 20331
rect 21102 20225 21136 20259
rect 21102 20153 21136 20187
rect 21102 20081 21136 20115
rect 21102 20009 21136 20043
rect 20605 -24417 20639 -24383
rect 20677 -24417 20711 -24383
rect 20555 -24531 20589 -24497
rect 20555 -24603 20589 -24569
rect 20555 -24675 20589 -24641
rect 20555 -24747 20589 -24713
rect 13667 -24849 13701 -24815
rect 13739 -24849 13773 -24815
rect 20555 -24819 20589 -24785
rect 20555 -24891 20589 -24857
rect 13617 -24963 13651 -24929
rect 13617 -25035 13651 -25001
rect 13789 -24963 13823 -24929
rect 13789 -25035 13823 -25001
rect 20555 -24963 20589 -24929
rect 20555 -25035 20589 -25001
rect 20727 -24531 20761 -24497
rect 20727 -24603 20761 -24569
rect 20727 -24675 20761 -24641
rect 20727 -24747 20761 -24713
rect 20727 -24819 20761 -24785
rect 20727 -24891 20761 -24857
rect 20727 -24963 20761 -24929
rect 20727 -25035 20761 -25001
<< metal1 >>
rect 20494 20659 21056 22366
rect 20494 20625 20506 20659
rect 20540 20625 20578 20659
rect 20612 20625 20650 20659
rect 20684 20625 20722 20659
rect 20756 20625 20794 20659
rect 20828 20625 20866 20659
rect 20900 20625 20938 20659
rect 20972 20625 21010 20659
rect 21044 20625 21056 20659
rect 20494 20613 21056 20625
rect 20408 20547 20454 20563
rect 20408 20513 20414 20547
rect 20448 20513 20454 20547
rect 20408 20475 20454 20513
rect 20408 20441 20414 20475
rect 20448 20441 20454 20475
rect 20408 20403 20454 20441
rect 20408 20369 20414 20403
rect 20448 20369 20454 20403
rect 20408 20331 20454 20369
rect 20408 20297 20414 20331
rect 20448 20297 20454 20331
rect 20408 20259 20454 20297
rect 20408 20225 20414 20259
rect 20448 20225 20454 20259
rect 20408 20187 20454 20225
rect 13853 20143 13983 20155
rect 13853 20109 13865 20143
rect 13899 20109 13937 20143
rect 13971 20109 13983 20143
rect 13853 20097 13983 20109
rect 20408 20153 20414 20187
rect 20448 20153 20454 20187
rect 20408 20115 20454 20153
rect 20408 20081 20414 20115
rect 20448 20081 20454 20115
rect 13809 20043 13855 20062
rect 13809 20009 13815 20043
rect 13849 20009 13855 20043
rect 13809 19913 13855 20009
rect 13981 20043 14027 20062
rect 13981 20009 13987 20043
rect 14021 20009 14027 20043
rect 13981 19913 14027 20009
rect 13809 19853 14027 19913
rect 20408 20043 20454 20081
rect 20408 20009 20414 20043
rect 20448 20009 20454 20043
rect 20408 19913 20454 20009
rect 20580 20547 20626 20563
rect 20580 20513 20586 20547
rect 20620 20513 20626 20547
rect 20580 20475 20626 20513
rect 20580 20441 20586 20475
rect 20620 20441 20626 20475
rect 20580 20403 20626 20441
rect 20580 20369 20586 20403
rect 20620 20369 20626 20403
rect 20580 20331 20626 20369
rect 20580 20297 20586 20331
rect 20620 20297 20626 20331
rect 20580 20259 20626 20297
rect 20580 20225 20586 20259
rect 20620 20225 20626 20259
rect 20580 20187 20626 20225
rect 20580 20153 20586 20187
rect 20620 20153 20626 20187
rect 20580 20115 20626 20153
rect 20580 20081 20586 20115
rect 20620 20081 20626 20115
rect 20580 20043 20626 20081
rect 20580 20009 20586 20043
rect 20620 20009 20626 20043
rect 20580 19913 20626 20009
rect 20752 20547 20798 20563
rect 20752 20513 20758 20547
rect 20792 20513 20798 20547
rect 20752 20475 20798 20513
rect 20752 20441 20758 20475
rect 20792 20441 20798 20475
rect 20752 20403 20798 20441
rect 20752 20369 20758 20403
rect 20792 20369 20798 20403
rect 20752 20331 20798 20369
rect 20752 20297 20758 20331
rect 20792 20297 20798 20331
rect 20752 20259 20798 20297
rect 20752 20225 20758 20259
rect 20792 20225 20798 20259
rect 20752 20187 20798 20225
rect 20752 20153 20758 20187
rect 20792 20153 20798 20187
rect 20752 20115 20798 20153
rect 20752 20081 20758 20115
rect 20792 20081 20798 20115
rect 20752 20043 20798 20081
rect 20752 20009 20758 20043
rect 20792 20009 20798 20043
rect 20752 19913 20798 20009
rect 20924 20547 20970 20563
rect 20924 20513 20930 20547
rect 20964 20513 20970 20547
rect 20924 20475 20970 20513
rect 20924 20441 20930 20475
rect 20964 20441 20970 20475
rect 20924 20403 20970 20441
rect 20924 20369 20930 20403
rect 20964 20369 20970 20403
rect 20924 20331 20970 20369
rect 20924 20297 20930 20331
rect 20964 20297 20970 20331
rect 20924 20259 20970 20297
rect 20924 20225 20930 20259
rect 20964 20225 20970 20259
rect 20924 20187 20970 20225
rect 20924 20153 20930 20187
rect 20964 20153 20970 20187
rect 20924 20115 20970 20153
rect 20924 20081 20930 20115
rect 20964 20081 20970 20115
rect 20924 20043 20970 20081
rect 20924 20009 20930 20043
rect 20964 20009 20970 20043
rect 20924 19913 20970 20009
rect 21096 20547 21142 20563
rect 21096 20513 21102 20547
rect 21136 20513 21142 20547
rect 21096 20475 21142 20513
rect 21096 20441 21102 20475
rect 21136 20441 21142 20475
rect 21096 20403 21142 20441
rect 21096 20369 21102 20403
rect 21136 20369 21142 20403
rect 21096 20331 21142 20369
rect 21096 20297 21102 20331
rect 21136 20297 21142 20331
rect 21096 20259 21142 20297
rect 21096 20225 21102 20259
rect 21136 20225 21142 20259
rect 21096 20187 21142 20225
rect 21096 20153 21102 20187
rect 21136 20153 21142 20187
rect 21096 20115 21142 20153
rect 21096 20081 21102 20115
rect 21136 20081 21142 20115
rect 21096 20043 21142 20081
rect 21096 20009 21102 20043
rect 21136 20009 21142 20043
rect 21096 19913 21142 20009
rect 20408 17651 21142 19913
rect 20593 -24383 20723 -24111
rect 20593 -24417 20605 -24383
rect 20639 -24417 20677 -24383
rect 20711 -24417 20723 -24383
rect 20593 -24429 20723 -24417
rect 20549 -24497 20595 -24481
rect 20549 -24531 20555 -24497
rect 20589 -24531 20595 -24497
rect 20549 -24569 20595 -24531
rect 20549 -24603 20555 -24569
rect 20589 -24603 20595 -24569
rect 20549 -24641 20595 -24603
rect 20549 -24675 20555 -24641
rect 20589 -24675 20595 -24641
rect 20549 -24713 20595 -24675
rect 20549 -24747 20555 -24713
rect 20589 -24747 20595 -24713
rect 20549 -24785 20595 -24747
rect 13655 -24815 13785 -24803
rect 13655 -24849 13667 -24815
rect 13701 -24849 13739 -24815
rect 13773 -24849 13785 -24815
rect 13655 -24861 13785 -24849
rect 20549 -24819 20555 -24785
rect 20589 -24819 20595 -24785
rect 20549 -24857 20595 -24819
rect 20549 -24891 20555 -24857
rect 20589 -24891 20595 -24857
rect 13611 -24929 13657 -24913
rect 13611 -24963 13617 -24929
rect 13651 -24963 13657 -24929
rect 13611 -25001 13657 -24963
rect 13611 -25035 13617 -25001
rect 13651 -25035 13657 -25001
rect 13611 -25131 13657 -25035
rect 13783 -24929 13829 -24913
rect 13783 -24963 13789 -24929
rect 13823 -24963 13829 -24929
rect 13783 -25001 13829 -24963
rect 13783 -25035 13789 -25001
rect 13823 -25035 13829 -25001
rect 13783 -25131 13829 -25035
rect 13611 -25191 13829 -25131
rect 20549 -24929 20595 -24891
rect 20549 -24963 20555 -24929
rect 20589 -24963 20595 -24929
rect 20549 -25001 20595 -24963
rect 20549 -25035 20555 -25001
rect 20589 -25035 20595 -25001
rect 20549 -25131 20595 -25035
rect 20721 -24497 20767 -24481
rect 20721 -24531 20727 -24497
rect 20761 -24531 20767 -24497
rect 20721 -24569 20767 -24531
rect 20721 -24603 20727 -24569
rect 20761 -24603 20767 -24569
rect 20721 -24641 20767 -24603
rect 20721 -24675 20727 -24641
rect 20761 -24675 20767 -24641
rect 20721 -24713 20767 -24675
rect 20721 -24747 20727 -24713
rect 20761 -24747 20767 -24713
rect 20721 -24785 20767 -24747
rect 20721 -24819 20727 -24785
rect 20761 -24819 20767 -24785
rect 20721 -24857 20767 -24819
rect 20721 -24891 20727 -24857
rect 20761 -24891 20767 -24857
rect 20721 -24929 20767 -24891
rect 20721 -24963 20727 -24929
rect 20761 -24963 20767 -24929
rect 20721 -25001 20767 -24963
rect 20721 -25035 20727 -25001
rect 20761 -25035 20767 -25001
rect 20721 -25131 20767 -25035
rect 20549 -25409 20767 -25131
<< obsm1 >>
rect 13892 19993 13944 20062
rect 20491 19993 20543 20563
rect 20663 19993 20715 20563
rect 20835 19993 20887 20563
rect 21007 19993 21059 20563
rect 13694 -25051 13746 -24913
rect 20632 -25051 20684 -24481
<< metal2 >>
rect 13892 19993 13944 20062
rect 20120 -24614 20684 -24486
rect 13694 -25046 13746 -24918
<< obsm2 >>
rect 20484 20415 20550 20569
rect 20656 20415 20722 20569
rect 20828 20415 20894 20569
rect 21000 20415 21066 20569
<< metal3 >>
rect 20484 20503 21836 20569
rect 20484 20415 20550 20503
rect 20656 20415 20722 20503
rect 20828 20415 20894 20503
rect 21000 20415 21836 20503
<< labels >>
rlabel locali s 1835 -41064 2397 -40469 8 B_P
port 1 nsew
rlabel metal3 s 21000 20415 21836 20503 6 D_N2
port 2 nsew
rlabel metal3 s 20828 20415 20894 20503 6 D_N2
port 2 nsew
rlabel metal3 s 20656 20415 20722 20503 6 D_N2
port 2 nsew
rlabel metal3 s 20484 20503 21836 20569 6 D_N2
port 2 nsew
rlabel metal3 s 20484 20415 20550 20503 6 D_N2
port 2 nsew
rlabel metal2 s 13694 -25046 13746 -24918 8 D_P
port 3 nsew
rlabel metal2 s 20120 -24614 20684 -24486 8 D_P2
port 4 nsew
rlabel metal1 s 13853 20097 13983 20155 6 G
port 5 nsew
rlabel metal1 s 20494 20613 21056 22366 6 G_N2
port 6 nsew
rlabel metal1 s 13655 -24861 13785 -24803 8 G_P
port 7 nsew
rlabel metal1 s 20593 -24429 20723 -24111 8 G_P2
port 8 nsew
rlabel locali s 1835 1730 2397 2325 6 NWELL
port 9 nsew
rlabel metal1 s 13981 19913 14027 20062 6 S
port 10 nsew
rlabel metal1 s 13809 19913 13855 20062 6 S
port 10 nsew
rlabel metal1 s 13809 19853 14027 19913 6 S
port 10 nsew
rlabel metal1 s 21096 19913 21142 20563 6 S_N2
port 11 nsew
rlabel metal1 s 20924 19913 20970 20563 6 S_N2
port 11 nsew
rlabel metal1 s 20752 19913 20798 20563 6 S_N2
port 11 nsew
rlabel metal1 s 20580 19913 20626 20563 6 S_N2
port 11 nsew
rlabel metal1 s 20408 19913 20454 20563 6 S_N2
port 11 nsew
rlabel metal1 s 20408 17651 21142 19913 6 S_N2
port 11 nsew
rlabel metal1 s 13783 -25131 13829 -24913 8 S_P
port 12 nsew
rlabel metal1 s 13611 -25131 13657 -24913 8 S_P
port 12 nsew
rlabel metal1 s 13611 -25191 13829 -25131 8 S_P
port 12 nsew
rlabel metal1 s 20721 -25131 20767 -24481 8 S_P2
port 13 nsew
rlabel metal1 s 20549 -25131 20595 -24481 8 S_P2
port 13 nsew
rlabel metal1 s 20549 -25409 20767 -25131 8 S_P2
port 13 nsew
rlabel locali s 12028 18138 12590 18733 6 VGND
port 14 nsew ground default
rlabel metal2 s 13892 19993 13944 20062 6 VPWR
port 15 nsew power default
<< properties >>
string FIXED_BBOX 0 -42794 311106 39640
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 10480152
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 10476062
<< end >>
