magic
tech sky130B
magscale 1 2
timestamp 1666464484
<< nwell >>
rect 1326 758 1860 1138
<< pwell >>
rect 103 558 1265 910
rect 117 132 1823 384
rect 117 110 590 132
rect 64 24 590 110
<< mvnmos >>
rect 182 584 282 884
rect 338 584 438 884
rect 494 584 594 884
rect 650 584 750 884
rect 930 584 1030 884
rect 1086 584 1186 884
<< mvpmos >>
rect 1445 824 1565 964
rect 1621 824 1741 964
<< mvnnmos >>
rect 738 158 918 358
rect 974 158 1154 358
rect 1328 158 1508 358
rect 1564 158 1744 358
<< nmoslvt >>
rect 196 158 226 358
rect 282 158 312 358
rect 368 158 398 358
rect 454 158 484 358
<< ndiff >>
rect 143 340 196 358
rect 143 306 151 340
rect 185 306 196 340
rect 143 272 196 306
rect 143 238 151 272
rect 185 238 196 272
rect 143 204 196 238
rect 143 170 151 204
rect 185 170 196 204
rect 143 158 196 170
rect 226 340 282 358
rect 226 306 237 340
rect 271 306 282 340
rect 226 272 282 306
rect 226 238 237 272
rect 271 238 282 272
rect 226 204 282 238
rect 226 170 237 204
rect 271 170 282 204
rect 226 158 282 170
rect 312 340 368 358
rect 312 306 323 340
rect 357 306 368 340
rect 312 272 368 306
rect 312 238 323 272
rect 357 238 368 272
rect 312 204 368 238
rect 312 170 323 204
rect 357 170 368 204
rect 312 158 368 170
rect 398 340 454 358
rect 398 306 409 340
rect 443 306 454 340
rect 398 272 454 306
rect 398 238 409 272
rect 443 238 454 272
rect 398 204 454 238
rect 398 170 409 204
rect 443 170 454 204
rect 398 158 454 170
rect 484 340 537 358
rect 484 306 495 340
rect 529 306 537 340
rect 484 272 537 306
rect 484 238 495 272
rect 529 238 537 272
rect 484 204 537 238
rect 484 170 495 204
rect 529 170 537 204
rect 484 158 537 170
<< mvndiff >>
rect 129 872 182 884
rect 129 838 137 872
rect 171 838 182 872
rect 129 804 182 838
rect 129 770 137 804
rect 171 770 182 804
rect 129 736 182 770
rect 129 702 137 736
rect 171 702 182 736
rect 129 668 182 702
rect 129 634 137 668
rect 171 634 182 668
rect 129 584 182 634
rect 282 872 338 884
rect 282 838 293 872
rect 327 838 338 872
rect 282 804 338 838
rect 282 770 293 804
rect 327 770 338 804
rect 282 736 338 770
rect 282 702 293 736
rect 327 702 338 736
rect 282 668 338 702
rect 282 634 293 668
rect 327 634 338 668
rect 282 584 338 634
rect 438 872 494 884
rect 438 838 449 872
rect 483 838 494 872
rect 438 804 494 838
rect 438 770 449 804
rect 483 770 494 804
rect 438 736 494 770
rect 438 702 449 736
rect 483 702 494 736
rect 438 668 494 702
rect 438 634 449 668
rect 483 634 494 668
rect 438 584 494 634
rect 594 872 650 884
rect 594 838 605 872
rect 639 838 650 872
rect 594 804 650 838
rect 594 770 605 804
rect 639 770 650 804
rect 594 736 650 770
rect 594 702 605 736
rect 639 702 650 736
rect 594 668 650 702
rect 594 634 605 668
rect 639 634 650 668
rect 594 584 650 634
rect 750 872 803 884
rect 750 838 761 872
rect 795 838 803 872
rect 750 804 803 838
rect 750 770 761 804
rect 795 770 803 804
rect 750 736 803 770
rect 750 702 761 736
rect 795 702 803 736
rect 750 668 803 702
rect 750 634 761 668
rect 795 634 803 668
rect 750 584 803 634
rect 877 872 930 884
rect 877 838 885 872
rect 919 838 930 872
rect 877 804 930 838
rect 877 770 885 804
rect 919 770 930 804
rect 877 736 930 770
rect 877 702 885 736
rect 919 702 930 736
rect 877 668 930 702
rect 877 634 885 668
rect 919 634 930 668
rect 877 584 930 634
rect 1030 872 1086 884
rect 1030 838 1041 872
rect 1075 838 1086 872
rect 1030 804 1086 838
rect 1030 770 1041 804
rect 1075 770 1086 804
rect 1030 736 1086 770
rect 1030 702 1041 736
rect 1075 702 1086 736
rect 1030 668 1086 702
rect 1030 634 1041 668
rect 1075 634 1086 668
rect 1030 584 1086 634
rect 1186 872 1239 884
rect 1186 838 1197 872
rect 1231 838 1239 872
rect 1186 804 1239 838
rect 1186 770 1197 804
rect 1231 770 1239 804
rect 1186 736 1239 770
rect 1186 702 1197 736
rect 1231 702 1239 736
rect 1186 668 1239 702
rect 1186 634 1197 668
rect 1231 634 1239 668
rect 1186 584 1239 634
rect 685 340 738 358
rect 685 306 693 340
rect 727 306 738 340
rect 685 272 738 306
rect 685 238 693 272
rect 727 238 738 272
rect 685 204 738 238
rect 685 170 693 204
rect 727 170 738 204
rect 685 158 738 170
rect 918 340 974 358
rect 918 306 929 340
rect 963 306 974 340
rect 918 272 974 306
rect 918 238 929 272
rect 963 238 974 272
rect 918 204 974 238
rect 918 170 929 204
rect 963 170 974 204
rect 918 158 974 170
rect 1154 340 1207 358
rect 1154 306 1165 340
rect 1199 306 1207 340
rect 1154 272 1207 306
rect 1154 238 1165 272
rect 1199 238 1207 272
rect 1154 204 1207 238
rect 1154 170 1165 204
rect 1199 170 1207 204
rect 1154 158 1207 170
rect 1275 346 1328 358
rect 1275 312 1283 346
rect 1317 312 1328 346
rect 1275 278 1328 312
rect 1275 244 1283 278
rect 1317 244 1328 278
rect 1275 210 1328 244
rect 1275 176 1283 210
rect 1317 176 1328 210
rect 1275 158 1328 176
rect 1508 346 1564 358
rect 1508 312 1519 346
rect 1553 312 1564 346
rect 1508 278 1564 312
rect 1508 244 1519 278
rect 1553 244 1564 278
rect 1508 210 1564 244
rect 1508 176 1519 210
rect 1553 176 1564 210
rect 1508 158 1564 176
rect 1744 346 1797 358
rect 1744 312 1755 346
rect 1789 312 1797 346
rect 1744 278 1797 312
rect 1744 244 1755 278
rect 1789 244 1797 278
rect 1744 210 1797 244
rect 1744 176 1755 210
rect 1789 176 1797 210
rect 1744 158 1797 176
<< mvpdiff >>
rect 1392 952 1445 964
rect 1392 918 1400 952
rect 1434 918 1445 952
rect 1392 884 1445 918
rect 1392 850 1400 884
rect 1434 850 1445 884
rect 1392 824 1445 850
rect 1565 952 1621 964
rect 1565 918 1576 952
rect 1610 918 1621 952
rect 1565 884 1621 918
rect 1565 850 1576 884
rect 1610 850 1621 884
rect 1565 824 1621 850
rect 1741 952 1794 964
rect 1741 918 1752 952
rect 1786 918 1794 952
rect 1741 884 1794 918
rect 1741 850 1752 884
rect 1786 850 1794 884
rect 1741 824 1794 850
<< ndiffc >>
rect 151 306 185 340
rect 151 238 185 272
rect 151 170 185 204
rect 237 306 271 340
rect 237 238 271 272
rect 237 170 271 204
rect 323 306 357 340
rect 323 238 357 272
rect 323 170 357 204
rect 409 306 443 340
rect 409 238 443 272
rect 409 170 443 204
rect 495 306 529 340
rect 495 238 529 272
rect 495 170 529 204
<< mvndiffc >>
rect 137 838 171 872
rect 137 770 171 804
rect 137 702 171 736
rect 137 634 171 668
rect 293 838 327 872
rect 293 770 327 804
rect 293 702 327 736
rect 293 634 327 668
rect 449 838 483 872
rect 449 770 483 804
rect 449 702 483 736
rect 449 634 483 668
rect 605 838 639 872
rect 605 770 639 804
rect 605 702 639 736
rect 605 634 639 668
rect 761 838 795 872
rect 761 770 795 804
rect 761 702 795 736
rect 761 634 795 668
rect 885 838 919 872
rect 885 770 919 804
rect 885 702 919 736
rect 885 634 919 668
rect 1041 838 1075 872
rect 1041 770 1075 804
rect 1041 702 1075 736
rect 1041 634 1075 668
rect 1197 838 1231 872
rect 1197 770 1231 804
rect 1197 702 1231 736
rect 1197 634 1231 668
rect 693 306 727 340
rect 693 238 727 272
rect 693 170 727 204
rect 929 306 963 340
rect 929 238 963 272
rect 929 170 963 204
rect 1165 306 1199 340
rect 1165 238 1199 272
rect 1165 170 1199 204
rect 1283 312 1317 346
rect 1283 244 1317 278
rect 1283 176 1317 210
rect 1519 312 1553 346
rect 1519 244 1553 278
rect 1519 176 1553 210
rect 1755 312 1789 346
rect 1755 244 1789 278
rect 1755 176 1789 210
<< mvpdiffc >>
rect 1400 918 1434 952
rect 1400 850 1434 884
rect 1576 918 1610 952
rect 1576 850 1610 884
rect 1752 918 1786 952
rect 1752 850 1786 884
<< psubdiff >>
rect 90 50 114 84
rect 148 50 192 84
rect 226 50 270 84
rect 304 50 348 84
rect 382 50 427 84
rect 461 50 506 84
rect 540 50 564 84
<< mvnsubdiff >>
rect 1392 1038 1416 1072
rect 1450 1038 1496 1072
rect 1530 1038 1576 1072
rect 1610 1038 1656 1072
rect 1690 1038 1736 1072
rect 1770 1038 1794 1072
<< psubdiffcont >>
rect 114 50 148 84
rect 192 50 226 84
rect 270 50 304 84
rect 348 50 382 84
rect 427 50 461 84
rect 506 50 540 84
<< mvnsubdiffcont >>
rect 1416 1038 1450 1072
rect 1496 1038 1530 1072
rect 1576 1038 1610 1072
rect 1656 1038 1690 1072
rect 1736 1038 1770 1072
<< poly >>
rect 1445 964 1565 996
rect 1621 964 1741 996
rect 182 884 282 916
rect 338 884 438 916
rect 494 884 594 916
rect 650 884 750 916
rect 930 884 1030 916
rect 1086 884 1186 916
rect 1445 771 1565 824
rect 1445 737 1494 771
rect 1528 737 1565 771
rect 1445 703 1565 737
rect 1445 669 1494 703
rect 1528 669 1565 703
rect 1445 653 1565 669
rect 1621 771 1741 824
rect 1621 737 1669 771
rect 1703 737 1741 771
rect 1621 703 1741 737
rect 1621 669 1669 703
rect 1703 669 1741 703
rect 1621 653 1741 669
rect 182 558 282 584
rect 338 558 438 584
rect 182 542 438 558
rect 182 508 198 542
rect 232 508 293 542
rect 327 508 388 542
rect 422 508 438 542
rect 182 492 438 508
rect 494 558 594 584
rect 650 558 750 584
rect 930 558 1030 584
rect 1086 558 1186 584
rect 494 542 1186 558
rect 494 508 510 542
rect 544 508 579 542
rect 613 508 648 542
rect 682 508 717 542
rect 751 508 786 542
rect 820 508 856 542
rect 890 508 926 542
rect 960 508 996 542
rect 1030 508 1066 542
rect 1100 508 1136 542
rect 1170 508 1186 542
rect 494 492 1186 508
rect 178 434 312 450
rect 178 400 194 434
rect 228 400 262 434
rect 296 400 312 434
rect 178 384 312 400
rect 196 358 226 384
rect 282 358 312 384
rect 368 434 502 450
rect 368 400 384 434
rect 418 400 452 434
rect 486 400 502 434
rect 368 384 502 400
rect 738 434 1744 450
rect 738 400 932 434
rect 966 400 1002 434
rect 1036 400 1072 434
rect 1106 400 1142 434
rect 1176 400 1211 434
rect 1245 400 1280 434
rect 1314 400 1349 434
rect 1383 400 1418 434
rect 1452 400 1487 434
rect 1521 400 1556 434
rect 1590 400 1625 434
rect 1659 400 1694 434
rect 1728 400 1744 434
rect 738 384 1744 400
rect 368 358 398 384
rect 454 358 484 384
rect 738 358 918 384
rect 974 358 1154 384
rect 1328 358 1508 384
rect 1564 358 1744 384
rect 196 126 226 158
rect 282 126 312 158
rect 368 126 398 158
rect 454 126 484 158
rect 738 126 918 158
rect 974 126 1154 158
rect 1328 126 1508 158
rect 1564 126 1744 158
<< polycont >>
rect 1494 737 1528 771
rect 1494 669 1528 703
rect 1669 737 1703 771
rect 1669 669 1703 703
rect 198 508 232 542
rect 293 508 327 542
rect 388 508 422 542
rect 510 508 544 542
rect 579 508 613 542
rect 648 508 682 542
rect 717 508 751 542
rect 786 508 820 542
rect 856 508 890 542
rect 926 508 960 542
rect 996 508 1030 542
rect 1066 508 1100 542
rect 1136 508 1170 542
rect 194 400 228 434
rect 262 400 296 434
rect 384 400 418 434
rect 452 400 486 434
rect 932 400 966 434
rect 1002 400 1036 434
rect 1072 400 1106 434
rect 1142 400 1176 434
rect 1211 400 1245 434
rect 1280 400 1314 434
rect 1349 400 1383 434
rect 1418 400 1452 434
rect 1487 400 1521 434
rect 1556 400 1590 434
rect 1625 400 1659 434
rect 1694 400 1728 434
<< locali >>
rect 1392 1069 1416 1072
rect 1450 1069 1496 1072
rect 1530 1069 1576 1072
rect 1610 1069 1656 1072
rect 1690 1069 1736 1072
rect 1392 1038 1411 1069
rect 1450 1038 1492 1069
rect 1530 1038 1573 1069
rect 1610 1038 1654 1069
rect 1690 1038 1735 1069
rect 1770 1038 1794 1072
rect 1445 1035 1492 1038
rect 1526 1035 1573 1038
rect 1607 1035 1654 1038
rect 1688 1035 1735 1038
rect 1400 952 1434 968
rect 137 872 171 888
rect 137 826 171 838
rect 293 872 327 888
rect 136 804 174 826
rect 136 792 137 804
rect 171 792 174 804
rect 293 804 327 838
rect 449 872 483 888
rect 449 826 483 838
rect 605 872 639 888
rect 137 736 171 770
rect 137 668 171 702
rect 137 618 171 634
rect 448 804 486 826
rect 448 792 449 804
rect 293 746 327 770
rect 293 674 327 702
rect 293 618 327 634
rect 483 792 486 804
rect 605 804 639 838
rect 761 872 795 888
rect 761 826 795 838
rect 885 872 919 888
rect 449 736 483 770
rect 449 668 483 702
rect 449 618 483 634
rect 739 804 777 826
rect 739 792 761 804
rect 885 804 919 838
rect 1041 872 1075 888
rect 1041 834 1075 838
rect 1197 872 1231 888
rect 605 736 639 770
rect 605 668 639 702
rect 605 623 639 634
rect 761 736 795 770
rect 761 668 795 702
rect 596 589 634 623
rect 761 618 795 634
rect 1040 804 1078 834
rect 1040 800 1041 804
rect 885 736 919 770
rect 885 668 919 702
rect 885 610 919 634
rect 1075 800 1078 804
rect 1197 804 1231 838
rect 1400 884 1434 918
rect 1400 834 1434 850
rect 1576 896 1610 918
rect 1576 834 1610 850
rect 1751 952 1819 968
rect 1751 918 1752 952
rect 1786 918 1819 952
rect 1751 884 1819 918
rect 1751 850 1752 884
rect 1786 850 1819 884
rect 1041 736 1075 770
rect 1041 668 1075 702
rect 1041 618 1075 634
rect 1370 800 1408 834
rect 1197 736 1231 770
rect 1197 668 1231 702
rect 1197 610 1231 634
rect 1477 771 1563 787
rect 1477 737 1494 771
rect 1528 737 1563 771
rect 1669 771 1703 787
rect 1477 703 1563 737
rect 1638 737 1669 747
rect 1638 713 1676 737
rect 1477 669 1494 703
rect 1528 669 1563 703
rect 1477 648 1563 669
rect 1669 703 1703 713
rect 1669 653 1703 669
rect 1477 614 1481 648
rect 1515 614 1553 648
rect 1751 619 1819 850
rect 1587 614 1819 619
rect 908 576 946 610
rect 1167 576 1205 610
rect 1477 576 1819 614
rect 182 508 198 542
rect 243 527 281 561
rect 232 508 293 527
rect 327 508 388 542
rect 422 508 438 542
rect 494 508 510 542
rect 544 508 579 542
rect 613 508 648 542
rect 682 508 717 542
rect 751 530 786 542
rect 820 530 856 542
rect 890 530 926 542
rect 960 530 996 542
rect 1030 530 1066 542
rect 751 508 769 530
rect 820 508 842 530
rect 890 508 915 530
rect 960 508 988 530
rect 1030 508 1062 530
rect 1100 508 1136 542
rect 1170 508 1186 542
rect 803 496 842 508
rect 876 496 915 508
rect 949 496 988 508
rect 1022 496 1062 508
rect 1096 496 1136 508
rect 178 440 199 474
rect 233 440 271 474
rect 305 440 312 474
rect 178 434 312 440
rect 178 400 194 434
rect 228 400 262 434
rect 296 400 312 434
rect 368 456 502 462
rect 368 434 432 456
rect 466 434 504 456
rect 368 400 384 434
rect 418 422 432 434
rect 486 422 504 434
rect 1471 434 1518 446
rect 1552 434 1598 446
rect 1632 434 1678 446
rect 418 400 452 422
rect 486 400 502 422
rect 810 377 848 411
rect 916 400 932 434
rect 966 400 1002 434
rect 1036 400 1072 434
rect 1106 400 1142 434
rect 1176 400 1211 434
rect 1245 400 1280 434
rect 1314 400 1349 434
rect 1383 400 1418 434
rect 1471 412 1487 434
rect 1552 412 1556 434
rect 1452 400 1487 412
rect 1521 400 1556 412
rect 1590 412 1598 434
rect 1659 412 1678 434
rect 1590 400 1625 412
rect 1659 400 1694 412
rect 1728 400 1744 434
rect 151 340 185 356
rect 151 272 185 306
rect 151 228 185 238
rect 151 156 185 170
rect 237 294 271 306
rect 237 204 271 238
rect 237 154 271 170
rect 323 340 357 356
rect 323 272 357 306
rect 323 228 357 238
rect 323 156 357 170
rect 776 358 882 377
rect 776 356 960 358
rect 409 294 443 306
rect 409 204 443 238
rect 409 154 443 170
rect 477 340 581 356
rect 693 355 727 356
rect 477 306 495 340
rect 529 306 581 340
rect 650 321 688 355
rect 722 340 727 355
rect 477 272 581 306
rect 477 238 495 272
rect 529 238 581 272
rect 477 209 581 238
rect 693 272 727 306
rect 511 204 549 209
rect 529 175 549 204
rect 693 204 727 238
rect 477 170 495 175
rect 529 170 581 175
rect 477 154 581 170
rect 693 154 727 170
rect 776 340 963 356
rect 1165 355 1199 356
rect 776 306 929 340
rect 1134 340 1172 355
rect 1134 321 1165 340
rect 1307 346 1345 366
rect 1317 332 1345 346
rect 1519 346 1553 362
rect 776 272 963 306
rect 776 238 929 272
rect 776 204 963 238
rect 776 170 929 204
rect 776 154 963 170
rect 1165 272 1199 306
rect 1165 204 1199 238
rect 1165 154 1199 170
rect 1283 278 1317 312
rect 1717 332 1755 366
rect 1519 292 1553 312
rect 1497 278 1535 292
rect 1497 258 1519 278
rect 1755 278 1789 312
rect 1283 210 1317 244
rect 1283 160 1317 176
rect 1519 210 1553 244
rect 1519 160 1553 176
rect 1755 210 1789 244
rect 1755 160 1789 176
rect 776 153 960 154
rect 109 50 114 84
rect 148 50 150 84
rect 184 50 192 84
rect 259 50 270 84
rect 334 50 348 84
rect 409 50 427 84
rect 484 50 506 84
rect 559 50 600 84
rect 634 50 675 84
rect 709 50 750 84
rect 784 50 825 84
rect 859 50 900 84
rect 934 50 975 84
rect 1009 50 1049 84
rect 1083 50 1123 84
rect 1157 50 1197 84
rect 1231 50 1271 84
rect 1305 50 1345 84
rect 1379 50 1419 84
rect 1453 50 1493 84
rect 1527 50 1567 84
rect 1601 50 1641 84
<< viali >>
rect 1411 1038 1416 1069
rect 1416 1038 1445 1069
rect 1492 1038 1496 1069
rect 1496 1038 1526 1069
rect 1573 1038 1576 1069
rect 1576 1038 1607 1069
rect 1654 1038 1656 1069
rect 1656 1038 1688 1069
rect 1735 1038 1736 1069
rect 1736 1038 1769 1069
rect 1411 1035 1445 1038
rect 1492 1035 1526 1038
rect 1573 1035 1607 1038
rect 1654 1035 1688 1038
rect 1735 1035 1769 1038
rect 102 792 136 826
rect 174 792 208 826
rect 414 792 448 826
rect 293 736 327 746
rect 293 712 327 736
rect 293 668 327 674
rect 293 640 327 668
rect 486 792 520 826
rect 705 792 739 826
rect 777 804 811 826
rect 777 792 795 804
rect 795 792 811 804
rect 562 589 596 623
rect 634 589 668 623
rect 1006 800 1040 834
rect 1078 800 1112 834
rect 1576 952 1610 968
rect 1576 934 1610 952
rect 1576 884 1610 896
rect 1576 862 1610 884
rect 1336 800 1370 834
rect 1408 800 1442 834
rect 1604 713 1638 747
rect 1676 737 1703 747
rect 1703 737 1710 747
rect 1676 713 1710 737
rect 1481 614 1515 648
rect 1553 614 1587 648
rect 874 576 908 610
rect 946 576 980 610
rect 1133 576 1167 610
rect 1205 576 1239 610
rect 209 542 243 561
rect 209 527 232 542
rect 232 527 243 542
rect 281 542 315 561
rect 281 527 293 542
rect 293 527 315 542
rect 769 508 786 530
rect 786 508 803 530
rect 842 508 856 530
rect 856 508 876 530
rect 915 508 926 530
rect 926 508 949 530
rect 988 508 996 530
rect 996 508 1022 530
rect 1062 508 1066 530
rect 1066 508 1096 530
rect 1136 508 1170 530
rect 769 496 803 508
rect 842 496 876 508
rect 915 496 949 508
rect 988 496 1022 508
rect 1062 496 1096 508
rect 1136 496 1170 508
rect 199 440 233 474
rect 271 440 305 474
rect 432 434 466 456
rect 432 422 452 434
rect 452 422 466 434
rect 504 422 538 456
rect 1437 434 1471 446
rect 1518 434 1552 446
rect 1598 434 1632 446
rect 1678 434 1712 446
rect 776 377 810 411
rect 848 377 882 411
rect 1437 412 1452 434
rect 1452 412 1471 434
rect 1518 412 1521 434
rect 1521 412 1552 434
rect 1598 412 1625 434
rect 1625 412 1632 434
rect 1678 412 1694 434
rect 1694 412 1712 434
rect 151 204 185 228
rect 151 194 185 204
rect 151 122 185 156
rect 237 340 271 366
rect 237 332 271 340
rect 237 272 271 294
rect 237 260 271 272
rect 323 204 357 228
rect 323 194 357 204
rect 323 122 357 156
rect 409 340 443 366
rect 409 332 443 340
rect 409 272 443 294
rect 409 260 443 272
rect 616 321 650 355
rect 688 340 722 355
rect 688 321 693 340
rect 693 321 722 340
rect 477 204 511 209
rect 477 175 495 204
rect 495 175 511 204
rect 549 175 583 209
rect 1100 321 1134 355
rect 1172 340 1206 355
rect 1172 321 1199 340
rect 1199 321 1206 340
rect 1273 346 1307 366
rect 1273 332 1283 346
rect 1283 332 1307 346
rect 1345 332 1379 366
rect 1683 332 1717 366
rect 1755 346 1789 366
rect 1755 332 1789 346
rect 1463 258 1497 292
rect 1535 278 1569 292
rect 1535 258 1553 278
rect 1553 258 1569 278
rect 75 50 109 84
rect 150 50 184 84
rect 225 50 226 84
rect 226 50 259 84
rect 300 50 304 84
rect 304 50 334 84
rect 375 50 382 84
rect 382 50 409 84
rect 450 50 461 84
rect 461 50 484 84
rect 525 50 540 84
rect 540 50 559 84
rect 600 50 634 84
rect 675 50 709 84
rect 750 50 784 84
rect 825 50 859 84
rect 900 50 934 84
rect 975 50 1009 84
rect 1049 50 1083 84
rect 1123 50 1157 84
rect 1197 50 1231 84
rect 1271 50 1305 84
rect 1345 50 1379 84
rect 1419 50 1453 84
rect 1493 50 1527 84
rect 1567 50 1601 84
rect 1641 50 1675 84
<< metal1 >>
rect 58 1069 1824 1076
rect 58 1035 1411 1069
rect 1445 1035 1492 1069
rect 1526 1035 1573 1069
rect 1607 1035 1654 1069
rect 1688 1035 1735 1069
rect 1769 1035 1824 1069
rect 58 968 1824 1035
rect 58 934 1576 968
rect 1610 934 1824 968
rect 58 896 1824 934
rect 58 874 1576 896
tri 1546 862 1558 874 ne
rect 1558 862 1576 874
rect 1610 874 1824 896
rect 1610 862 1616 874
tri 1558 850 1570 862 ne
rect 1570 850 1616 862
tri 1616 850 1640 874 nw
rect 994 834 1454 840
rect 90 826 899 832
rect 90 792 102 826
rect 136 792 174 826
rect 208 792 414 826
rect 448 792 486 826
rect 520 792 705 826
rect 739 792 777 826
rect 811 800 899 826
tri 899 800 931 832 sw
rect 994 800 1006 834
rect 1040 800 1078 834
rect 1112 800 1336 834
rect 1370 800 1408 834
rect 1442 800 1454 834
rect 811 792 931 800
tri 931 792 939 800 sw
rect 994 794 1454 800
tri 1454 794 1463 803 sw
tri 1325 792 1327 794 ne
rect 1327 792 1463 794
tri 1463 792 1465 794 sw
rect 90 786 939 792
tri 879 758 907 786 ne
rect 907 758 939 786
rect 77 746 333 758
tri 907 747 918 758 ne
rect 918 747 939 758
tri 939 747 984 792 sw
tri 1327 753 1366 792 ne
rect 1366 753 1465 792
tri 1465 753 1504 792 sw
tri 1366 747 1372 753 ne
rect 1372 747 1722 753
rect 77 712 293 746
rect 327 712 333 746
tri 918 726 939 747 ne
rect 939 726 984 747
tri 984 726 1005 747 sw
tri 1372 726 1393 747 ne
rect 1393 726 1604 747
tri 939 713 952 726 ne
rect 952 713 1301 726
tri 1301 713 1314 726 sw
tri 1393 713 1406 726 ne
rect 1406 713 1604 726
rect 1638 713 1676 747
rect 1710 713 1722 747
rect 77 674 333 712
tri 952 684 981 713 ne
rect 981 707 1314 713
tri 1314 707 1320 713 sw
tri 1406 707 1412 713 ne
rect 1412 707 1722 713
rect 981 684 1320 707
rect 77 640 293 674
rect 327 640 333 674
tri 1263 654 1293 684 ne
rect 1293 654 1320 684
tri 1320 654 1373 707 sw
tri 1293 648 1299 654 ne
rect 1299 648 1599 654
tri 1299 646 1301 648 ne
rect 1301 646 1481 648
rect 77 628 333 640
tri 1301 629 1318 646 ne
rect 1318 629 1481 646
tri 62 277 77 292 se
rect 77 277 154 628
rect 550 623 684 629
rect 550 589 562 623
rect 596 589 634 623
rect 668 614 684 623
tri 684 614 699 629 sw
tri 1318 616 1331 629 ne
rect 1331 616 1481 629
rect 668 610 699 614
tri 699 610 703 614 sw
rect 862 610 1251 616
tri 1331 614 1333 616 ne
rect 1333 614 1481 616
rect 1515 614 1553 648
rect 1587 614 1599 648
rect 668 608 703 610
tri 703 608 705 610 sw
rect 668 589 705 608
rect 550 587 705 589
tri 705 587 726 608 sw
rect 550 583 726 587
tri 666 576 673 583 ne
rect 673 576 726 583
tri 673 567 682 576 ne
rect 682 567 726 576
rect 862 576 874 610
rect 908 576 946 610
rect 980 576 1133 610
rect 1167 576 1205 610
rect 1239 576 1251 610
tri 1333 608 1339 614 ne
rect 1339 608 1599 614
rect 862 570 1251 576
tri 1251 570 1258 577 sw
rect 197 561 329 567
rect 197 527 209 561
rect 243 527 281 561
rect 315 527 329 561
tri 682 551 698 567 ne
tri 397 530 398 531 se
rect 398 530 652 531
rect 197 521 329 527
tri 388 521 397 530 se
rect 397 521 652 530
tri 363 496 388 521 se
rect 388 503 652 521
rect 388 496 406 503
tri 406 496 413 503 nw
tri 355 488 363 496 se
rect 363 488 398 496
tri 398 488 406 496 nw
tri 351 484 355 488 se
rect 355 484 394 488
tri 394 484 398 488 nw
rect 187 474 317 480
rect 187 440 199 474
rect 233 440 271 474
rect 305 440 317 474
rect 187 434 317 440
tri 340 395 351 406 se
rect 351 395 379 484
tri 379 469 394 484 nw
rect 420 456 550 462
rect 420 422 432 456
rect 466 422 504 456
rect 538 422 550 456
rect 420 416 550 422
tri 323 378 340 395 se
rect 340 394 379 395
rect 340 378 363 394
tri 363 378 379 394 nw
rect 624 389 652 503
rect 698 446 726 567
tri 1218 536 1252 570 ne
rect 1252 536 1258 570
rect 757 530 1182 536
tri 1252 530 1258 536 ne
tri 1258 530 1298 570 sw
rect 757 496 769 530
rect 803 496 842 530
rect 876 496 915 530
rect 949 496 988 530
rect 1022 496 1062 530
rect 1096 496 1136 530
rect 1170 496 1182 530
tri 1258 527 1261 530 ne
rect 757 490 1182 496
tri 726 446 731 451 sw
rect 698 417 731 446
tri 731 417 760 446 sw
rect 698 411 894 417
tri 652 389 658 395 sw
rect 698 389 776 411
tri 621 378 624 381 se
rect 624 378 658 389
rect 231 377 362 378
tri 362 377 363 378 nw
rect 231 373 358 377
tri 358 373 362 377 nw
rect 231 366 351 373
tri 351 366 358 373 nw
rect 403 366 449 378
tri 620 377 621 378 se
rect 621 377 658 378
tri 658 377 670 389 sw
tri 746 377 758 389 ne
rect 758 377 776 389
rect 810 377 848 411
rect 882 377 894 411
tri 616 373 620 377 se
rect 620 373 670 377
tri 670 373 674 377 sw
tri 758 373 762 377 ne
rect 762 373 894 377
tri 449 366 456 373 sw
tri 609 366 616 373 se
rect 616 371 674 373
tri 674 371 676 373 sw
tri 762 371 764 373 ne
rect 764 371 894 373
rect 1261 372 1298 530
rect 1425 446 1724 452
rect 1425 412 1437 446
rect 1471 412 1518 446
rect 1552 412 1598 446
rect 1632 412 1678 446
rect 1712 412 1724 446
rect 1425 406 1724 412
tri 1298 372 1332 406 sw
rect 616 366 676 371
tri 676 366 681 371 sw
rect 1261 366 1801 372
rect 231 332 237 366
rect 271 339 324 366
tri 324 339 351 366 nw
rect 271 332 317 339
tri 317 332 324 339 nw
rect 403 332 409 366
rect 443 355 456 366
tri 456 355 467 366 sw
tri 604 361 609 366 se
rect 609 361 681 366
tri 681 361 686 366 sw
rect 604 355 734 361
tri 734 355 740 361 sw
tri 1082 355 1088 361 se
rect 1088 355 1218 361
rect 443 339 467 355
tri 467 339 483 355 sw
rect 443 332 533 339
rect 231 326 311 332
tri 311 326 317 332 nw
rect 403 326 533 332
tri 533 326 546 339 sw
rect 231 321 306 326
tri 306 321 311 326 nw
rect 403 321 546 326
tri 546 321 551 326 sw
rect 604 321 616 355
rect 650 321 688 355
rect 722 343 740 355
tri 740 343 752 355 sw
tri 1070 343 1082 355 se
rect 1082 343 1100 355
rect 722 321 1100 343
rect 1134 321 1172 355
rect 1206 321 1218 355
rect 1261 332 1273 366
rect 1307 332 1345 366
rect 1379 332 1683 366
rect 1717 332 1755 366
rect 1789 332 1801 366
rect 1261 326 1801 332
rect 231 294 279 321
tri 279 294 306 321 nw
rect 403 315 551 321
tri 551 315 557 321 sw
rect 604 315 1218 321
rect 403 298 557 315
tri 557 298 574 315 sw
rect 403 294 574 298
tri 45 260 62 277 se
rect 62 260 154 277
tri 154 260 171 277 sw
rect 231 260 237 294
rect 271 260 277 294
tri 277 292 279 294 nw
tri 43 258 45 260 se
rect 45 258 171 260
tri 171 258 173 260 sw
tri 38 253 43 258 se
rect 43 253 173 258
tri 173 253 178 258 sw
rect 38 240 178 253
tri 178 240 191 253 sw
rect 231 248 277 260
rect 403 260 409 294
rect 443 293 574 294
rect 443 292 482 293
tri 482 292 483 293 nw
tri 523 292 524 293 ne
rect 524 292 574 293
tri 574 292 580 298 sw
tri 1445 292 1451 298 se
rect 1451 292 1581 298
rect 443 287 477 292
tri 477 287 482 292 nw
tri 524 287 529 292 ne
rect 529 287 580 292
tri 580 287 585 292 sw
tri 1440 287 1445 292 se
rect 1445 287 1463 292
rect 443 283 473 287
tri 473 283 477 287 nw
tri 529 283 533 287 ne
rect 533 283 1463 287
rect 443 277 467 283
tri 467 277 473 283 nw
tri 533 277 539 283 ne
rect 539 277 1463 283
rect 443 260 449 277
rect 403 248 449 260
tri 449 259 467 277 nw
tri 539 259 557 277 ne
rect 557 259 1463 277
tri 1444 258 1445 259 ne
rect 1445 258 1463 259
rect 1497 258 1535 292
rect 1569 258 1581 292
tri 1445 253 1450 258 ne
rect 1450 253 1581 258
tri 1450 252 1451 253 ne
rect 1451 252 1581 253
tri 1699 252 1700 253 se
rect 1700 252 1829 253
tri 1695 248 1699 252 se
rect 1699 248 1829 252
tri 1687 240 1695 248 se
rect 1695 240 1829 248
rect 38 228 191 240
tri 191 228 203 240 sw
tri 305 228 317 240 se
rect 317 228 363 240
rect 38 194 151 228
rect 185 220 203 228
tri 203 220 211 228 sw
tri 297 220 305 228 se
rect 305 220 323 228
rect 185 194 323 220
rect 357 220 363 228
tri 363 220 383 240 sw
tri 1667 220 1687 240 se
rect 1687 220 1829 240
rect 357 209 1829 220
rect 357 194 477 209
rect 38 175 477 194
rect 511 175 549 209
rect 583 175 1829 209
rect 38 156 1829 175
rect 38 122 151 156
rect 185 122 323 156
rect 357 122 1829 156
rect 38 84 1829 122
rect 38 50 75 84
rect 109 50 150 84
rect 184 50 225 84
rect 259 50 300 84
rect 334 50 375 84
rect 409 50 450 84
rect 484 50 525 84
rect 559 50 600 84
rect 634 50 675 84
rect 709 50 750 84
rect 784 50 825 84
rect 859 50 900 84
rect 934 50 975 84
rect 1009 50 1049 84
rect 1083 50 1123 84
rect 1157 50 1197 84
rect 1231 50 1271 84
rect 1305 50 1345 84
rect 1379 50 1419 84
rect 1453 50 1493 84
rect 1527 50 1567 84
rect 1601 50 1641 84
rect 1675 50 1829 84
rect 38 39 1829 50
use sky130_fd_pr__nfet_01v8__example_55959141808496  sky130_fd_pr__nfet_01v8__example_55959141808496_0
timestamp 1666464484
transform -1 0 1744 0 -1 358
box -1 0 417 1
use sky130_fd_pr__nfet_01v8__example_55959141808497  sky130_fd_pr__nfet_01v8__example_55959141808497_0
timestamp 1666464484
transform -1 0 1154 0 1 158
box -1 0 417 1
use sky130_fd_pr__nfet_01v8__example_55959141808498  sky130_fd_pr__nfet_01v8__example_55959141808498_0
timestamp 1666464484
transform -1 0 484 0 1 158
box -1 0 117 1
use sky130_fd_pr__nfet_01v8__example_55959141808498  sky130_fd_pr__nfet_01v8__example_55959141808498_1
timestamp 1666464484
transform -1 0 312 0 1 158
box -1 0 117 1
use sky130_fd_pr__nfet_01v8__example_55959141808582  sky130_fd_pr__nfet_01v8__example_55959141808582_0
timestamp 1666464484
transform -1 0 1186 0 -1 884
box -1 0 257 1
use sky130_fd_pr__nfet_01v8__example_55959141808583  sky130_fd_pr__nfet_01v8__example_55959141808583_0
timestamp 1666464484
transform -1 0 438 0 -1 884
box -1 0 257 1
use sky130_fd_pr__nfet_01v8__example_55959141808583  sky130_fd_pr__nfet_01v8__example_55959141808583_1
timestamp 1666464484
transform -1 0 750 0 -1 884
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_55959141808580  sky130_fd_pr__pfet_01v8__example_55959141808580_0
timestamp 1666464484
transform -1 0 1565 0 -1 964
box -1 0 121 1
use sky130_fd_pr__pfet_01v8__example_55959141808580  sky130_fd_pr__pfet_01v8__example_55959141808580_1
timestamp 1666464484
transform 1 0 1621 0 -1 964
box -1 0 121 1
<< labels >>
flabel metal1 s 1626 414 1654 442 3 FreeSans 280 0 0 0 VPWR_LV
port 1 nsew
flabel metal1 s 245 529 273 557 3 FreeSans 280 0 0 0 RST_H
port 2 nsew
flabel metal1 s 1372 805 1400 833 3 FreeSans 280 0 0 0 OUT_H_N
port 3 nsew
flabel metal1 s 455 425 483 453 3 FreeSans 280 0 0 0 IN
port 4 nsew
flabel metal1 s 240 445 268 473 3 FreeSans 280 0 0 0 IN_B
port 5 nsew
flabel metal1 s 1108 498 1136 526 3 FreeSans 280 0 0 0 HLD_H_N
port 6 nsew
flabel metal1 s 1541 619 1569 647 3 FreeSans 280 270 0 0 OUT_H
port 7 nsew
flabel metal1 s 73 174 101 202 3 FreeSans 280 0 0 0 VGND
port 8 nsew
flabel metal1 s 1491 984 1519 1012 3 FreeSans 280 0 0 0 VPWR_HV
port 9 nsew
<< properties >>
string GDS_END 43537918
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 43518734
<< end >>
