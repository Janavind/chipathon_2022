magic
tech sky130A
magscale 1 2
timestamp 1666199351
<< nwell >>
rect -38 261 590 582
<< pwell >>
rect 1 21 419 183
rect 29 -17 63 21
<< locali >>
rect 17 149 85 265
rect 119 259 191 493
rect 337 259 403 493
rect 119 203 403 259
rect 119 136 191 203
rect 119 51 243 136
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 19 299 85 527
rect 231 293 297 527
rect 443 293 509 527
rect 19 17 85 115
rect 335 17 401 155
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
<< metal1 >>
rect 0 561 552 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 0 496 552 527
rect 0 17 552 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
rect 0 -48 552 -17
<< labels >>
rlabel locali s 17 149 85 265 6 A
port 1 nsew signal input
rlabel metal1 s 0 -48 552 48 8 VGND
port 2 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 3 nsew ground bidirectional
rlabel pwell s 1 21 419 183 6 VNB
port 3 nsew ground bidirectional
rlabel nwell s -38 261 590 582 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 496 552 592 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 119 51 243 136 6 Y
port 6 nsew signal output
rlabel locali s 119 136 191 203 6 Y
port 6 nsew signal output
rlabel locali s 119 203 403 259 6 Y
port 6 nsew signal output
rlabel locali s 337 259 403 493 6 Y
port 6 nsew signal output
rlabel locali s 119 259 191 493 6 Y
port 6 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 552 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3333294
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3328254
<< end >>
