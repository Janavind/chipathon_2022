magic
tech sky130A
magscale 1 2
timestamp 1666464484
<< pwell >>
rect -10 2190 2276 2276
rect -10 76 76 2190
rect 1551 1747 1572 1796
rect 2190 76 2276 2190
rect -10 -10 2276 76
<< locali >>
rect 16 2216 2250 2250
rect 16 50 50 2216
rect 2216 50 2250 2216
rect 16 16 2250 50
<< metal1 >>
rect 0 2259 2266 2266
rect 0 2207 56 2259
rect 108 2207 136 2259
rect 188 2207 216 2259
rect 268 2207 296 2259
rect 348 2207 376 2259
rect 428 2207 456 2259
rect 508 2207 536 2259
rect 588 2207 616 2259
rect 668 2207 696 2259
rect 748 2207 776 2259
rect 828 2207 856 2259
rect 908 2207 936 2259
rect 988 2207 1016 2259
rect 1068 2207 1198 2259
rect 1250 2207 1278 2259
rect 1330 2207 1358 2259
rect 1410 2207 1438 2259
rect 1490 2207 1518 2259
rect 1570 2207 1598 2259
rect 1650 2207 1678 2259
rect 1730 2207 1758 2259
rect 1810 2207 1838 2259
rect 1890 2207 1918 2259
rect 1970 2207 1998 2259
rect 2050 2207 2078 2259
rect 2130 2207 2158 2259
rect 2210 2207 2266 2259
rect 0 2200 2266 2207
rect 0 2130 66 2200
rect 0 2078 7 2130
rect 59 2078 66 2130
rect 0 2050 66 2078
rect 0 1998 7 2050
rect 59 1998 66 2050
rect 0 1970 66 1998
rect 0 1918 7 1970
rect 59 1918 66 1970
rect 0 1890 66 1918
rect 0 1838 7 1890
rect 59 1838 66 1890
rect 0 1810 66 1838
rect 0 1758 7 1810
rect 59 1758 66 1810
rect 0 1730 66 1758
rect 0 1678 7 1730
rect 59 1678 66 1730
rect 0 1650 66 1678
rect 0 1598 7 1650
rect 59 1598 66 1650
rect 0 1570 66 1598
rect 0 1518 7 1570
rect 59 1518 66 1570
rect 0 1490 66 1518
rect 0 1438 7 1490
rect 59 1438 66 1490
rect 0 1410 66 1438
rect 0 1358 7 1410
rect 59 1358 66 1410
rect 0 1330 66 1358
rect 0 1278 7 1330
rect 59 1278 66 1330
rect 0 1250 66 1278
rect 0 1198 7 1250
rect 59 1198 66 1250
rect 0 1068 66 1198
rect 0 1016 7 1068
rect 59 1016 66 1068
rect 0 988 66 1016
rect 0 936 7 988
rect 59 936 66 988
rect 0 908 66 936
rect 0 856 7 908
rect 59 856 66 908
rect 0 828 66 856
rect 0 776 7 828
rect 59 776 66 828
rect 0 748 66 776
rect 0 696 7 748
rect 59 696 66 748
rect 0 668 66 696
rect 0 616 7 668
rect 59 616 66 668
rect 0 588 66 616
rect 0 536 7 588
rect 59 536 66 588
rect 0 508 66 536
rect 0 456 7 508
rect 59 456 66 508
rect 0 428 66 456
rect 0 376 7 428
rect 59 376 66 428
rect 0 348 66 376
rect 0 296 7 348
rect 59 296 66 348
rect 0 268 66 296
rect 0 216 7 268
rect 59 216 66 268
rect 0 188 66 216
rect 0 136 7 188
rect 59 136 66 188
rect 0 66 66 136
rect 94 1164 122 2172
rect 150 1192 178 2200
rect 206 1164 234 2172
rect 262 1192 290 2200
rect 318 1164 346 2172
rect 374 1192 402 2200
rect 430 1164 458 2172
rect 486 1192 514 2200
rect 542 1164 570 2172
rect 598 1192 626 2200
rect 654 1164 682 2172
rect 710 1192 738 2200
rect 766 1164 794 2172
rect 822 1192 850 2200
rect 878 1164 906 2172
rect 934 1192 962 2200
rect 990 1164 1018 2172
rect 1046 1192 1074 2200
rect 1102 2119 1164 2172
rect 1102 2067 1107 2119
rect 1159 2067 1164 2119
rect 1102 2039 1164 2067
rect 1102 1987 1107 2039
rect 1159 1987 1164 2039
rect 1102 1959 1164 1987
rect 1102 1907 1107 1959
rect 1159 1907 1164 1959
rect 1102 1879 1164 1907
rect 1102 1827 1107 1879
rect 1159 1827 1164 1879
rect 1102 1799 1164 1827
rect 1102 1747 1107 1799
rect 1159 1747 1164 1799
rect 1102 1719 1164 1747
rect 1102 1667 1107 1719
rect 1159 1667 1164 1719
rect 1102 1639 1164 1667
rect 1102 1587 1107 1639
rect 1159 1587 1164 1639
rect 1102 1559 1164 1587
rect 1102 1507 1107 1559
rect 1159 1507 1164 1559
rect 1102 1479 1164 1507
rect 1102 1427 1107 1479
rect 1159 1427 1164 1479
rect 1102 1399 1164 1427
rect 1102 1347 1107 1399
rect 1159 1347 1164 1399
rect 1102 1319 1164 1347
rect 1102 1267 1107 1319
rect 1159 1267 1164 1319
rect 1102 1239 1164 1267
rect 1102 1187 1107 1239
rect 1159 1187 1164 1239
rect 1192 1192 1220 2200
rect 1102 1164 1164 1187
rect 1248 1164 1276 2172
rect 1304 1192 1332 2200
rect 1360 1164 1388 2172
rect 1416 1192 1444 2200
rect 1472 1164 1500 2172
rect 1528 1192 1556 2200
rect 1584 1164 1612 2172
rect 1640 1192 1668 2200
rect 1696 1164 1724 2172
rect 1752 1192 1780 2200
rect 1808 1164 1836 2172
rect 1864 1192 1892 2200
rect 1920 1164 1948 2172
rect 1976 1192 2004 2200
rect 2032 1164 2060 2172
rect 2088 1192 2116 2200
rect 2144 1164 2172 2172
rect 94 1159 2172 1164
rect 94 1107 147 1159
rect 199 1107 227 1159
rect 279 1107 307 1159
rect 359 1107 387 1159
rect 439 1107 467 1159
rect 519 1107 547 1159
rect 599 1107 627 1159
rect 679 1107 707 1159
rect 759 1107 787 1159
rect 839 1107 867 1159
rect 919 1107 947 1159
rect 999 1107 1027 1159
rect 1079 1107 1107 1159
rect 1159 1107 1187 1159
rect 1239 1107 1267 1159
rect 1319 1107 1347 1159
rect 1399 1107 1427 1159
rect 1479 1107 1507 1159
rect 1559 1107 1587 1159
rect 1639 1107 1667 1159
rect 1719 1107 1747 1159
rect 1799 1107 1827 1159
rect 1879 1107 1907 1159
rect 1959 1107 1987 1159
rect 2039 1107 2067 1159
rect 2119 1107 2172 1159
rect 94 1102 2172 1107
rect 94 94 122 1102
rect 150 66 178 1074
rect 206 94 234 1102
rect 262 66 290 1074
rect 318 94 346 1102
rect 374 66 402 1074
rect 430 94 458 1102
rect 486 66 514 1074
rect 542 94 570 1102
rect 598 66 626 1074
rect 654 94 682 1102
rect 710 66 738 1074
rect 766 94 794 1102
rect 822 66 850 1074
rect 878 94 906 1102
rect 934 66 962 1074
rect 990 94 1018 1102
rect 1102 1079 1164 1102
rect 1046 66 1074 1074
rect 1102 1027 1107 1079
rect 1159 1027 1164 1079
rect 1102 999 1164 1027
rect 1102 947 1107 999
rect 1159 947 1164 999
rect 1102 919 1164 947
rect 1102 867 1107 919
rect 1159 867 1164 919
rect 1102 839 1164 867
rect 1102 787 1107 839
rect 1159 787 1164 839
rect 1102 759 1164 787
rect 1102 707 1107 759
rect 1159 707 1164 759
rect 1102 679 1164 707
rect 1102 627 1107 679
rect 1159 627 1164 679
rect 1102 599 1164 627
rect 1102 547 1107 599
rect 1159 547 1164 599
rect 1102 519 1164 547
rect 1102 467 1107 519
rect 1159 467 1164 519
rect 1102 439 1164 467
rect 1102 387 1107 439
rect 1159 387 1164 439
rect 1102 359 1164 387
rect 1102 307 1107 359
rect 1159 307 1164 359
rect 1102 279 1164 307
rect 1102 227 1107 279
rect 1159 227 1164 279
rect 1102 199 1164 227
rect 1102 147 1107 199
rect 1159 147 1164 199
rect 1102 94 1164 147
rect 1192 66 1220 1074
rect 1248 94 1276 1102
rect 1304 66 1332 1074
rect 1360 94 1388 1102
rect 1416 66 1444 1074
rect 1472 94 1500 1102
rect 1528 66 1556 1074
rect 1584 94 1612 1102
rect 1640 66 1668 1074
rect 1696 94 1724 1102
rect 1752 66 1780 1074
rect 1808 94 1836 1102
rect 1864 66 1892 1074
rect 1920 94 1948 1102
rect 1976 66 2004 1074
rect 2032 94 2060 1102
rect 2088 66 2116 1074
rect 2144 94 2172 1102
rect 2200 2130 2266 2200
rect 2200 2078 2207 2130
rect 2259 2078 2266 2130
rect 2200 2050 2266 2078
rect 2200 1998 2207 2050
rect 2259 1998 2266 2050
rect 2200 1970 2266 1998
rect 2200 1918 2207 1970
rect 2259 1918 2266 1970
rect 2200 1890 2266 1918
rect 2200 1838 2207 1890
rect 2259 1838 2266 1890
rect 2200 1810 2266 1838
rect 2200 1758 2207 1810
rect 2259 1758 2266 1810
rect 2200 1730 2266 1758
rect 2200 1678 2207 1730
rect 2259 1678 2266 1730
rect 2200 1650 2266 1678
rect 2200 1598 2207 1650
rect 2259 1598 2266 1650
rect 2200 1570 2266 1598
rect 2200 1518 2207 1570
rect 2259 1518 2266 1570
rect 2200 1490 2266 1518
rect 2200 1438 2207 1490
rect 2259 1438 2266 1490
rect 2200 1410 2266 1438
rect 2200 1358 2207 1410
rect 2259 1358 2266 1410
rect 2200 1330 2266 1358
rect 2200 1278 2207 1330
rect 2259 1278 2266 1330
rect 2200 1250 2266 1278
rect 2200 1198 2207 1250
rect 2259 1198 2266 1250
rect 2200 1068 2266 1198
rect 2200 1016 2207 1068
rect 2259 1016 2266 1068
rect 2200 988 2266 1016
rect 2200 936 2207 988
rect 2259 936 2266 988
rect 2200 908 2266 936
rect 2200 856 2207 908
rect 2259 856 2266 908
rect 2200 828 2266 856
rect 2200 776 2207 828
rect 2259 776 2266 828
rect 2200 748 2266 776
rect 2200 696 2207 748
rect 2259 696 2266 748
rect 2200 668 2266 696
rect 2200 616 2207 668
rect 2259 616 2266 668
rect 2200 588 2266 616
rect 2200 536 2207 588
rect 2259 536 2266 588
rect 2200 508 2266 536
rect 2200 456 2207 508
rect 2259 456 2266 508
rect 2200 428 2266 456
rect 2200 376 2207 428
rect 2259 376 2266 428
rect 2200 348 2266 376
rect 2200 296 2207 348
rect 2259 296 2266 348
rect 2200 268 2266 296
rect 2200 216 2207 268
rect 2259 216 2266 268
rect 2200 188 2266 216
rect 2200 136 2207 188
rect 2259 136 2266 188
rect 2200 66 2266 136
rect 0 59 2266 66
rect 0 7 56 59
rect 108 7 136 59
rect 188 7 216 59
rect 268 7 296 59
rect 348 7 376 59
rect 428 7 456 59
rect 508 7 536 59
rect 588 7 616 59
rect 668 7 696 59
rect 748 7 776 59
rect 828 7 856 59
rect 908 7 936 59
rect 988 7 1016 59
rect 1068 7 1198 59
rect 1250 7 1278 59
rect 1330 7 1358 59
rect 1410 7 1438 59
rect 1490 7 1518 59
rect 1570 7 1598 59
rect 1650 7 1678 59
rect 1730 7 1758 59
rect 1810 7 1838 59
rect 1890 7 1918 59
rect 1970 7 1998 59
rect 2050 7 2078 59
rect 2130 7 2158 59
rect 2210 7 2266 59
rect 0 0 2266 7
<< via1 >>
rect 56 2207 108 2259
rect 136 2207 188 2259
rect 216 2207 268 2259
rect 296 2207 348 2259
rect 376 2207 428 2259
rect 456 2207 508 2259
rect 536 2207 588 2259
rect 616 2207 668 2259
rect 696 2207 748 2259
rect 776 2207 828 2259
rect 856 2207 908 2259
rect 936 2207 988 2259
rect 1016 2207 1068 2259
rect 1198 2207 1250 2259
rect 1278 2207 1330 2259
rect 1358 2207 1410 2259
rect 1438 2207 1490 2259
rect 1518 2207 1570 2259
rect 1598 2207 1650 2259
rect 1678 2207 1730 2259
rect 1758 2207 1810 2259
rect 1838 2207 1890 2259
rect 1918 2207 1970 2259
rect 1998 2207 2050 2259
rect 2078 2207 2130 2259
rect 2158 2207 2210 2259
rect 7 2078 59 2130
rect 7 1998 59 2050
rect 7 1918 59 1970
rect 7 1838 59 1890
rect 7 1758 59 1810
rect 7 1678 59 1730
rect 7 1598 59 1650
rect 7 1518 59 1570
rect 7 1438 59 1490
rect 7 1358 59 1410
rect 7 1278 59 1330
rect 7 1198 59 1250
rect 7 1016 59 1068
rect 7 936 59 988
rect 7 856 59 908
rect 7 776 59 828
rect 7 696 59 748
rect 7 616 59 668
rect 7 536 59 588
rect 7 456 59 508
rect 7 376 59 428
rect 7 296 59 348
rect 7 216 59 268
rect 7 136 59 188
rect 1107 2067 1159 2119
rect 1107 1987 1159 2039
rect 1107 1907 1159 1959
rect 1107 1827 1159 1879
rect 1107 1747 1159 1799
rect 1107 1667 1159 1719
rect 1107 1587 1159 1639
rect 1107 1507 1159 1559
rect 1107 1427 1159 1479
rect 1107 1347 1159 1399
rect 1107 1267 1159 1319
rect 1107 1187 1159 1239
rect 147 1107 199 1159
rect 227 1107 279 1159
rect 307 1107 359 1159
rect 387 1107 439 1159
rect 467 1107 519 1159
rect 547 1107 599 1159
rect 627 1107 679 1159
rect 707 1107 759 1159
rect 787 1107 839 1159
rect 867 1107 919 1159
rect 947 1107 999 1159
rect 1027 1107 1079 1159
rect 1107 1107 1159 1159
rect 1187 1107 1239 1159
rect 1267 1107 1319 1159
rect 1347 1107 1399 1159
rect 1427 1107 1479 1159
rect 1507 1107 1559 1159
rect 1587 1107 1639 1159
rect 1667 1107 1719 1159
rect 1747 1107 1799 1159
rect 1827 1107 1879 1159
rect 1907 1107 1959 1159
rect 1987 1107 2039 1159
rect 2067 1107 2119 1159
rect 1107 1027 1159 1079
rect 1107 947 1159 999
rect 1107 867 1159 919
rect 1107 787 1159 839
rect 1107 707 1159 759
rect 1107 627 1159 679
rect 1107 547 1159 599
rect 1107 467 1159 519
rect 1107 387 1159 439
rect 1107 307 1159 359
rect 1107 227 1159 279
rect 1107 147 1159 199
rect 2207 2078 2259 2130
rect 2207 1998 2259 2050
rect 2207 1918 2259 1970
rect 2207 1838 2259 1890
rect 2207 1758 2259 1810
rect 2207 1678 2259 1730
rect 2207 1598 2259 1650
rect 2207 1518 2259 1570
rect 2207 1438 2259 1490
rect 2207 1358 2259 1410
rect 2207 1278 2259 1330
rect 2207 1198 2259 1250
rect 2207 1016 2259 1068
rect 2207 936 2259 988
rect 2207 856 2259 908
rect 2207 776 2259 828
rect 2207 696 2259 748
rect 2207 616 2259 668
rect 2207 536 2259 588
rect 2207 456 2259 508
rect 2207 376 2259 428
rect 2207 296 2259 348
rect 2207 216 2259 268
rect 2207 136 2259 188
rect 56 7 108 59
rect 136 7 188 59
rect 216 7 268 59
rect 296 7 348 59
rect 376 7 428 59
rect 456 7 508 59
rect 536 7 588 59
rect 616 7 668 59
rect 696 7 748 59
rect 776 7 828 59
rect 856 7 908 59
rect 936 7 988 59
rect 1016 7 1068 59
rect 1198 7 1250 59
rect 1278 7 1330 59
rect 1358 7 1410 59
rect 1438 7 1490 59
rect 1518 7 1570 59
rect 1598 7 1650 59
rect 1678 7 1730 59
rect 1758 7 1810 59
rect 1838 7 1890 59
rect 1918 7 1970 59
rect 1998 7 2050 59
rect 2078 7 2130 59
rect 2158 7 2210 59
<< metal2 >>
rect 0 2261 1074 2266
rect 0 2259 78 2261
rect 134 2259 204 2261
rect 260 2259 330 2261
rect 386 2259 456 2261
rect 512 2259 582 2261
rect 638 2259 708 2261
rect 764 2259 834 2261
rect 890 2259 960 2261
rect 1016 2259 1074 2261
rect 0 2207 56 2259
rect 134 2207 136 2259
rect 188 2207 204 2259
rect 268 2207 296 2259
rect 428 2207 456 2259
rect 512 2207 536 2259
rect 668 2207 696 2259
rect 764 2207 776 2259
rect 828 2207 834 2259
rect 908 2207 936 2259
rect 1068 2207 1074 2259
rect 0 2205 78 2207
rect 134 2205 204 2207
rect 260 2205 330 2207
rect 386 2205 456 2207
rect 512 2205 582 2207
rect 638 2205 708 2207
rect 764 2205 834 2207
rect 890 2205 960 2207
rect 1016 2205 1074 2207
rect 0 2200 1074 2205
rect 1192 2261 2266 2266
rect 1192 2259 1250 2261
rect 1306 2259 1376 2261
rect 1432 2259 1502 2261
rect 1558 2259 1628 2261
rect 1684 2259 1754 2261
rect 1810 2259 1880 2261
rect 1936 2259 2006 2261
rect 2062 2259 2132 2261
rect 2188 2259 2266 2261
rect 1192 2207 1198 2259
rect 1330 2207 1358 2259
rect 1432 2207 1438 2259
rect 1490 2207 1502 2259
rect 1570 2207 1598 2259
rect 1730 2207 1754 2259
rect 1810 2207 1838 2259
rect 1970 2207 1998 2259
rect 2062 2207 2078 2259
rect 2130 2207 2132 2259
rect 2210 2207 2266 2259
rect 1192 2205 1250 2207
rect 1306 2205 1376 2207
rect 1432 2205 1502 2207
rect 1558 2205 1628 2207
rect 1684 2205 1754 2207
rect 1810 2205 1880 2207
rect 1936 2205 2006 2207
rect 2062 2205 2132 2207
rect 2188 2205 2266 2207
rect 1192 2200 2266 2205
rect 0 2188 66 2200
rect 0 2132 5 2188
rect 61 2132 66 2188
rect 1102 2172 1164 2200
rect 2200 2188 2266 2200
rect 94 2169 2172 2172
rect 94 2144 1105 2169
rect 0 2130 66 2132
rect 0 2078 7 2130
rect 59 2116 66 2130
rect 59 2088 1074 2116
rect 1102 2113 1105 2144
rect 1161 2144 2172 2169
rect 1161 2113 1164 2144
rect 2200 2132 2205 2188
rect 2261 2132 2266 2188
rect 2200 2130 2266 2132
rect 2200 2116 2207 2130
rect 59 2078 66 2088
rect 0 2062 66 2078
rect 0 2006 5 2062
rect 61 2006 66 2062
rect 1102 2067 1107 2113
rect 1159 2067 1164 2113
rect 1192 2088 2207 2116
rect 1102 2060 1164 2067
rect 2200 2078 2207 2088
rect 2259 2078 2266 2130
rect 2200 2062 2266 2078
rect 94 2043 2172 2060
rect 94 2032 1105 2043
rect 0 1998 7 2006
rect 59 2004 66 2006
rect 59 1998 1074 2004
rect 0 1976 1074 1998
rect 1102 1987 1105 2032
rect 1161 2032 2172 2043
rect 1161 1987 1164 2032
rect 2200 2006 2205 2062
rect 2261 2006 2266 2062
rect 2200 2004 2207 2006
rect 0 1970 66 1976
rect 0 1936 7 1970
rect 59 1936 66 1970
rect 1102 1959 1164 1987
rect 1192 1998 2207 2004
rect 2259 1998 2266 2006
rect 1192 1976 2266 1998
rect 1102 1948 1107 1959
rect 0 1880 5 1936
rect 61 1892 66 1936
rect 94 1920 1107 1948
rect 1102 1917 1107 1920
rect 1159 1948 1164 1959
rect 2200 1970 2266 1976
rect 1159 1920 2172 1948
rect 2200 1936 2207 1970
rect 2259 1936 2266 1970
rect 1159 1917 1164 1920
rect 61 1880 1074 1892
rect 0 1838 7 1880
rect 59 1864 1074 1880
rect 59 1838 66 1864
rect 0 1810 66 1838
rect 1102 1861 1105 1917
rect 1161 1861 1164 1917
rect 2200 1892 2205 1936
rect 1192 1880 2205 1892
rect 2261 1880 2266 1936
rect 1192 1864 2207 1880
rect 1102 1836 1107 1861
rect 0 1754 5 1810
rect 61 1780 66 1810
rect 94 1827 1107 1836
rect 1159 1836 1164 1861
rect 2200 1838 2207 1864
rect 2259 1838 2266 1880
rect 1159 1827 2172 1836
rect 94 1808 2172 1827
rect 2200 1810 2266 1838
rect 1102 1799 1164 1808
rect 1102 1791 1107 1799
rect 1159 1791 1164 1799
rect 61 1754 1074 1780
rect 0 1752 1074 1754
rect 0 1730 66 1752
rect 0 1684 7 1730
rect 59 1684 66 1730
rect 1102 1735 1105 1791
rect 1161 1735 1164 1791
rect 2200 1780 2205 1810
rect 1192 1754 2205 1780
rect 2261 1754 2266 1810
rect 1192 1752 2266 1754
rect 1102 1724 1164 1735
rect 2200 1730 2266 1752
rect 94 1719 2172 1724
rect 94 1696 1107 1719
rect 0 1628 5 1684
rect 61 1668 66 1684
rect 61 1640 1074 1668
rect 1102 1667 1107 1696
rect 1159 1696 2172 1719
rect 1159 1667 1164 1696
rect 2200 1684 2207 1730
rect 2259 1684 2266 1730
rect 2200 1668 2205 1684
rect 1102 1665 1164 1667
rect 61 1628 66 1640
rect 0 1598 7 1628
rect 59 1598 66 1628
rect 1102 1612 1105 1665
rect 0 1570 66 1598
rect 94 1609 1105 1612
rect 1161 1612 1164 1665
rect 1192 1640 2205 1668
rect 2200 1628 2205 1640
rect 2261 1628 2266 1684
rect 1161 1609 2172 1612
rect 94 1587 1107 1609
rect 1159 1587 2172 1609
rect 94 1584 2172 1587
rect 2200 1598 2207 1628
rect 2259 1598 2266 1628
rect 0 1558 7 1570
rect 59 1558 66 1570
rect 0 1502 5 1558
rect 61 1556 66 1558
rect 1102 1559 1164 1584
rect 61 1528 1074 1556
rect 1102 1539 1107 1559
rect 1159 1539 1164 1559
rect 2200 1570 2266 1598
rect 2200 1558 2207 1570
rect 2259 1558 2266 1570
rect 2200 1556 2205 1558
rect 61 1502 66 1528
rect 0 1490 66 1502
rect 1102 1500 1105 1539
rect 0 1438 7 1490
rect 59 1444 66 1490
rect 94 1483 1105 1500
rect 1161 1500 1164 1539
rect 1192 1528 2205 1556
rect 2200 1502 2205 1528
rect 2261 1502 2266 1558
rect 1161 1483 2172 1500
rect 94 1479 2172 1483
rect 94 1472 1107 1479
rect 59 1438 1074 1444
rect 0 1432 1074 1438
rect 0 1376 5 1432
rect 61 1416 1074 1432
rect 1102 1427 1107 1472
rect 1159 1472 2172 1479
rect 2200 1490 2266 1502
rect 1159 1427 1164 1472
rect 2200 1444 2207 1490
rect 61 1376 66 1416
rect 1102 1413 1164 1427
rect 1192 1438 2207 1444
rect 2259 1438 2266 1490
rect 1192 1432 2266 1438
rect 1192 1416 2205 1432
rect 1102 1388 1105 1413
rect 0 1358 7 1376
rect 59 1358 66 1376
rect 94 1360 1105 1388
rect 0 1332 66 1358
rect 1102 1357 1105 1360
rect 1161 1388 1164 1413
rect 1161 1360 2172 1388
rect 2200 1376 2205 1416
rect 2261 1376 2266 1432
rect 1161 1357 1164 1360
rect 1102 1347 1107 1357
rect 1159 1347 1164 1357
rect 0 1330 1074 1332
rect 0 1306 7 1330
rect 59 1306 1074 1330
rect 0 1250 5 1306
rect 61 1304 1074 1306
rect 1102 1319 1164 1347
rect 2200 1358 2207 1376
rect 2259 1358 2266 1376
rect 2200 1332 2266 1358
rect 61 1250 66 1304
rect 1102 1287 1107 1319
rect 1159 1287 1164 1319
rect 1192 1330 2266 1332
rect 1192 1306 2207 1330
rect 2259 1306 2266 1330
rect 1192 1304 2205 1306
rect 1102 1276 1105 1287
rect 0 1198 7 1250
rect 59 1220 66 1250
rect 94 1248 1105 1276
rect 1161 1276 1164 1287
rect 1102 1231 1105 1248
rect 1161 1248 2172 1276
rect 2200 1250 2205 1304
rect 2261 1250 2266 1306
rect 1161 1231 1164 1248
rect 59 1198 1074 1220
rect 0 1192 1074 1198
rect 1102 1187 1107 1231
rect 1159 1187 1164 1231
rect 2200 1220 2207 1250
rect 1192 1198 2207 1220
rect 2259 1198 2266 1250
rect 1192 1192 2266 1198
rect 1102 1164 1164 1187
rect 66 1161 2200 1164
rect 66 1105 97 1161
rect 153 1159 223 1161
rect 279 1159 349 1161
rect 405 1159 475 1161
rect 531 1159 601 1161
rect 657 1159 727 1161
rect 783 1159 853 1161
rect 909 1159 979 1161
rect 1035 1159 1105 1161
rect 1161 1159 1231 1161
rect 1287 1159 1357 1161
rect 1413 1159 1483 1161
rect 1539 1159 1609 1161
rect 1665 1159 1735 1161
rect 1791 1159 1861 1161
rect 1917 1159 1987 1161
rect 2043 1159 2113 1161
rect 199 1107 223 1159
rect 279 1107 307 1159
rect 439 1107 467 1159
rect 531 1107 547 1159
rect 599 1107 601 1159
rect 679 1107 707 1159
rect 783 1107 787 1159
rect 839 1107 853 1159
rect 919 1107 947 1159
rect 1079 1107 1105 1159
rect 1161 1107 1187 1159
rect 1319 1107 1347 1159
rect 1413 1107 1427 1159
rect 1479 1107 1483 1159
rect 1559 1107 1587 1159
rect 1665 1107 1667 1159
rect 1719 1107 1735 1159
rect 1799 1107 1827 1159
rect 1959 1107 1987 1159
rect 2043 1107 2067 1159
rect 153 1105 223 1107
rect 279 1105 349 1107
rect 405 1105 475 1107
rect 531 1105 601 1107
rect 657 1105 727 1107
rect 783 1105 853 1107
rect 909 1105 979 1107
rect 1035 1105 1105 1107
rect 1161 1105 1231 1107
rect 1287 1105 1357 1107
rect 1413 1105 1483 1107
rect 1539 1105 1609 1107
rect 1665 1105 1735 1107
rect 1791 1105 1861 1107
rect 1917 1105 1987 1107
rect 2043 1105 2113 1107
rect 2169 1105 2200 1161
rect 66 1102 2200 1105
rect 1102 1079 1164 1102
rect 0 1068 1074 1074
rect 0 1016 7 1068
rect 59 1046 1074 1068
rect 59 1016 66 1046
rect 1102 1035 1107 1079
rect 1159 1035 1164 1079
rect 1192 1068 2266 1074
rect 1192 1046 2207 1068
rect 1102 1018 1105 1035
rect 0 960 5 1016
rect 61 962 66 1016
rect 94 990 1105 1018
rect 1161 1018 1164 1035
rect 1102 979 1105 990
rect 1161 990 2172 1018
rect 2200 1016 2207 1046
rect 2259 1016 2266 1068
rect 1161 979 1164 990
rect 61 960 1074 962
rect 0 936 7 960
rect 59 936 1074 960
rect 0 934 1074 936
rect 1102 947 1107 979
rect 1159 947 1164 979
rect 2200 962 2205 1016
rect 0 908 66 934
rect 0 890 7 908
rect 59 890 66 908
rect 1102 919 1164 947
rect 1192 960 2205 962
rect 2261 960 2266 1016
rect 1192 936 2207 960
rect 2259 936 2266 960
rect 1192 934 2266 936
rect 1102 909 1107 919
rect 1159 909 1164 919
rect 1102 906 1105 909
rect 0 834 5 890
rect 61 850 66 890
rect 94 878 1105 906
rect 1102 853 1105 878
rect 1161 906 1164 909
rect 2200 908 2266 934
rect 1161 878 2172 906
rect 2200 890 2207 908
rect 2259 890 2266 908
rect 1161 853 1164 878
rect 61 834 1074 850
rect 0 828 1074 834
rect 0 776 7 828
rect 59 822 1074 828
rect 1102 839 1164 853
rect 2200 850 2205 890
rect 59 776 66 822
rect 1102 794 1107 839
rect 0 764 66 776
rect 94 787 1107 794
rect 1159 794 1164 839
rect 1192 834 2205 850
rect 2261 834 2266 890
rect 1192 828 2266 834
rect 1192 822 2207 828
rect 1159 787 2172 794
rect 94 783 2172 787
rect 94 766 1105 783
rect 0 708 5 764
rect 61 738 66 764
rect 61 710 1074 738
rect 1102 727 1105 766
rect 1161 766 2172 783
rect 2200 776 2207 822
rect 2259 776 2266 828
rect 1161 727 1164 766
rect 2200 764 2266 776
rect 2200 738 2205 764
rect 61 708 66 710
rect 0 696 7 708
rect 59 696 66 708
rect 0 668 66 696
rect 1102 707 1107 727
rect 1159 707 1164 727
rect 1192 710 2205 738
rect 1102 682 1164 707
rect 2200 708 2205 710
rect 2261 708 2266 764
rect 2200 696 2207 708
rect 2259 696 2266 708
rect 0 638 7 668
rect 59 638 66 668
rect 94 679 2172 682
rect 94 657 1107 679
rect 1159 657 2172 679
rect 94 654 1105 657
rect 0 582 5 638
rect 61 626 66 638
rect 61 598 1074 626
rect 1102 601 1105 654
rect 1161 654 2172 657
rect 2200 668 2266 696
rect 1161 601 1164 654
rect 2200 638 2207 668
rect 2259 638 2266 668
rect 2200 626 2205 638
rect 1102 599 1164 601
rect 61 582 66 598
rect 0 536 7 582
rect 59 536 66 582
rect 1102 570 1107 599
rect 94 547 1107 570
rect 1159 570 1164 599
rect 1192 598 2205 626
rect 2200 582 2205 598
rect 2261 582 2266 638
rect 1159 547 2172 570
rect 94 542 2172 547
rect 0 514 66 536
rect 1102 531 1164 542
rect 0 512 1074 514
rect 0 456 5 512
rect 61 486 1074 512
rect 61 456 66 486
rect 1102 475 1105 531
rect 1161 475 1164 531
rect 2200 536 2207 582
rect 2259 536 2266 582
rect 2200 514 2266 536
rect 1192 512 2266 514
rect 1192 486 2205 512
rect 1102 467 1107 475
rect 1159 467 1164 475
rect 1102 458 1164 467
rect 0 428 66 456
rect 94 439 2172 458
rect 94 430 1107 439
rect 0 386 7 428
rect 59 402 66 428
rect 1102 405 1107 430
rect 1159 430 2172 439
rect 2200 456 2205 486
rect 2261 456 2266 512
rect 1159 405 1164 430
rect 59 386 1074 402
rect 0 330 5 386
rect 61 374 1074 386
rect 61 330 66 374
rect 1102 349 1105 405
rect 1161 349 1164 405
rect 2200 428 2266 456
rect 2200 402 2207 428
rect 1192 386 2207 402
rect 2259 386 2266 428
rect 1192 374 2205 386
rect 1102 346 1107 349
rect 0 296 7 330
rect 59 296 66 330
rect 94 318 1107 346
rect 0 290 66 296
rect 1102 307 1107 318
rect 1159 346 1164 349
rect 1159 318 2172 346
rect 2200 330 2205 374
rect 2261 330 2266 386
rect 1159 307 1164 318
rect 0 268 1074 290
rect 0 260 7 268
rect 59 262 1074 268
rect 1102 279 1164 307
rect 2200 296 2207 330
rect 2259 296 2266 330
rect 2200 290 2266 296
rect 59 260 66 262
rect 0 204 5 260
rect 61 204 66 260
rect 1102 234 1105 279
rect 94 223 1105 234
rect 1161 234 1164 279
rect 1192 268 2266 290
rect 1192 262 2207 268
rect 2200 260 2207 262
rect 2259 260 2266 268
rect 1161 223 2172 234
rect 94 206 2172 223
rect 0 188 66 204
rect 0 136 7 188
rect 59 178 66 188
rect 1102 199 1164 206
rect 59 150 1074 178
rect 1102 153 1107 199
rect 1159 153 1164 199
rect 2200 204 2205 260
rect 2261 204 2266 260
rect 2200 188 2266 204
rect 2200 178 2207 188
rect 59 136 66 150
rect 0 134 66 136
rect 0 78 5 134
rect 61 78 66 134
rect 1102 122 1105 153
rect 94 97 1105 122
rect 1161 122 1164 153
rect 1192 150 2207 178
rect 2200 136 2207 150
rect 2259 136 2266 188
rect 2200 134 2266 136
rect 1161 97 2172 122
rect 94 94 2172 97
rect 0 66 66 78
rect 1102 66 1164 94
rect 2200 78 2205 134
rect 2261 78 2266 134
rect 2200 66 2266 78
rect 0 61 1074 66
rect 0 59 78 61
rect 134 59 204 61
rect 260 59 330 61
rect 386 59 456 61
rect 512 59 582 61
rect 638 59 708 61
rect 764 59 834 61
rect 890 59 960 61
rect 1016 59 1074 61
rect 0 7 56 59
rect 134 7 136 59
rect 188 7 204 59
rect 268 7 296 59
rect 428 7 456 59
rect 512 7 536 59
rect 668 7 696 59
rect 764 7 776 59
rect 828 7 834 59
rect 908 7 936 59
rect 1068 7 1074 59
rect 0 5 78 7
rect 134 5 204 7
rect 260 5 330 7
rect 386 5 456 7
rect 512 5 582 7
rect 638 5 708 7
rect 764 5 834 7
rect 890 5 960 7
rect 1016 5 1074 7
rect 0 0 1074 5
rect 1192 61 2266 66
rect 1192 59 1250 61
rect 1306 59 1376 61
rect 1432 59 1502 61
rect 1558 59 1628 61
rect 1684 59 1754 61
rect 1810 59 1880 61
rect 1936 59 2006 61
rect 2062 59 2132 61
rect 2188 59 2266 61
rect 1192 7 1198 59
rect 1330 7 1358 59
rect 1432 7 1438 59
rect 1490 7 1502 59
rect 1570 7 1598 59
rect 1730 7 1754 59
rect 1810 7 1838 59
rect 1970 7 1998 59
rect 2062 7 2078 59
rect 2130 7 2132 59
rect 2210 7 2266 59
rect 1192 5 1250 7
rect 1306 5 1376 7
rect 1432 5 1502 7
rect 1558 5 1628 7
rect 1684 5 1754 7
rect 1810 5 1880 7
rect 1936 5 2006 7
rect 2062 5 2132 7
rect 2188 5 2266 7
rect 1192 0 2266 5
<< via2 >>
rect 78 2259 134 2261
rect 204 2259 260 2261
rect 330 2259 386 2261
rect 456 2259 512 2261
rect 582 2259 638 2261
rect 708 2259 764 2261
rect 834 2259 890 2261
rect 960 2259 1016 2261
rect 78 2207 108 2259
rect 108 2207 134 2259
rect 204 2207 216 2259
rect 216 2207 260 2259
rect 330 2207 348 2259
rect 348 2207 376 2259
rect 376 2207 386 2259
rect 456 2207 508 2259
rect 508 2207 512 2259
rect 582 2207 588 2259
rect 588 2207 616 2259
rect 616 2207 638 2259
rect 708 2207 748 2259
rect 748 2207 764 2259
rect 834 2207 856 2259
rect 856 2207 890 2259
rect 960 2207 988 2259
rect 988 2207 1016 2259
rect 78 2205 134 2207
rect 204 2205 260 2207
rect 330 2205 386 2207
rect 456 2205 512 2207
rect 582 2205 638 2207
rect 708 2205 764 2207
rect 834 2205 890 2207
rect 960 2205 1016 2207
rect 1250 2259 1306 2261
rect 1376 2259 1432 2261
rect 1502 2259 1558 2261
rect 1628 2259 1684 2261
rect 1754 2259 1810 2261
rect 1880 2259 1936 2261
rect 2006 2259 2062 2261
rect 2132 2259 2188 2261
rect 1250 2207 1278 2259
rect 1278 2207 1306 2259
rect 1376 2207 1410 2259
rect 1410 2207 1432 2259
rect 1502 2207 1518 2259
rect 1518 2207 1558 2259
rect 1628 2207 1650 2259
rect 1650 2207 1678 2259
rect 1678 2207 1684 2259
rect 1754 2207 1758 2259
rect 1758 2207 1810 2259
rect 1880 2207 1890 2259
rect 1890 2207 1918 2259
rect 1918 2207 1936 2259
rect 2006 2207 2050 2259
rect 2050 2207 2062 2259
rect 2132 2207 2158 2259
rect 2158 2207 2188 2259
rect 1250 2205 1306 2207
rect 1376 2205 1432 2207
rect 1502 2205 1558 2207
rect 1628 2205 1684 2207
rect 1754 2205 1810 2207
rect 1880 2205 1936 2207
rect 2006 2205 2062 2207
rect 2132 2205 2188 2207
rect 5 2132 61 2188
rect 1105 2119 1161 2169
rect 1105 2113 1107 2119
rect 1107 2113 1159 2119
rect 1159 2113 1161 2119
rect 2205 2132 2261 2188
rect 5 2050 61 2062
rect 5 2006 7 2050
rect 7 2006 59 2050
rect 59 2006 61 2050
rect 1105 2039 1161 2043
rect 1105 1987 1107 2039
rect 1107 1987 1159 2039
rect 1159 1987 1161 2039
rect 2205 2050 2261 2062
rect 2205 2006 2207 2050
rect 2207 2006 2259 2050
rect 2259 2006 2261 2050
rect 5 1918 7 1936
rect 7 1918 59 1936
rect 59 1918 61 1936
rect 5 1890 61 1918
rect 5 1880 7 1890
rect 7 1880 59 1890
rect 59 1880 61 1890
rect 1105 1907 1107 1917
rect 1107 1907 1159 1917
rect 1159 1907 1161 1917
rect 1105 1879 1161 1907
rect 1105 1861 1107 1879
rect 1107 1861 1159 1879
rect 1159 1861 1161 1879
rect 2205 1918 2207 1936
rect 2207 1918 2259 1936
rect 2259 1918 2261 1936
rect 2205 1890 2261 1918
rect 2205 1880 2207 1890
rect 2207 1880 2259 1890
rect 2259 1880 2261 1890
rect 5 1758 7 1810
rect 7 1758 59 1810
rect 59 1758 61 1810
rect 5 1754 61 1758
rect 1105 1747 1107 1791
rect 1107 1747 1159 1791
rect 1159 1747 1161 1791
rect 1105 1735 1161 1747
rect 2205 1758 2207 1810
rect 2207 1758 2259 1810
rect 2259 1758 2261 1810
rect 2205 1754 2261 1758
rect 5 1678 7 1684
rect 7 1678 59 1684
rect 59 1678 61 1684
rect 5 1650 61 1678
rect 5 1628 7 1650
rect 7 1628 59 1650
rect 59 1628 61 1650
rect 2205 1678 2207 1684
rect 2207 1678 2259 1684
rect 2259 1678 2261 1684
rect 1105 1639 1161 1665
rect 1105 1609 1107 1639
rect 1107 1609 1159 1639
rect 1159 1609 1161 1639
rect 2205 1650 2261 1678
rect 2205 1628 2207 1650
rect 2207 1628 2259 1650
rect 2259 1628 2261 1650
rect 5 1518 7 1558
rect 7 1518 59 1558
rect 59 1518 61 1558
rect 5 1502 61 1518
rect 1105 1507 1107 1539
rect 1107 1507 1159 1539
rect 1159 1507 1161 1539
rect 1105 1483 1161 1507
rect 2205 1518 2207 1558
rect 2207 1518 2259 1558
rect 2259 1518 2261 1558
rect 2205 1502 2261 1518
rect 5 1410 61 1432
rect 5 1376 7 1410
rect 7 1376 59 1410
rect 59 1376 61 1410
rect 1105 1399 1161 1413
rect 1105 1357 1107 1399
rect 1107 1357 1159 1399
rect 1159 1357 1161 1399
rect 2205 1410 2261 1432
rect 2205 1376 2207 1410
rect 2207 1376 2259 1410
rect 2259 1376 2261 1410
rect 5 1278 7 1306
rect 7 1278 59 1306
rect 59 1278 61 1306
rect 5 1250 61 1278
rect 1105 1267 1107 1287
rect 1107 1267 1159 1287
rect 1159 1267 1161 1287
rect 1105 1239 1161 1267
rect 2205 1278 2207 1306
rect 2207 1278 2259 1306
rect 2259 1278 2261 1306
rect 2205 1250 2261 1278
rect 1105 1231 1107 1239
rect 1107 1231 1159 1239
rect 1159 1231 1161 1239
rect 97 1159 153 1161
rect 223 1159 279 1161
rect 349 1159 405 1161
rect 475 1159 531 1161
rect 601 1159 657 1161
rect 727 1159 783 1161
rect 853 1159 909 1161
rect 979 1159 1035 1161
rect 1105 1159 1161 1161
rect 1231 1159 1287 1161
rect 1357 1159 1413 1161
rect 1483 1159 1539 1161
rect 1609 1159 1665 1161
rect 1735 1159 1791 1161
rect 1861 1159 1917 1161
rect 1987 1159 2043 1161
rect 2113 1159 2169 1161
rect 97 1107 147 1159
rect 147 1107 153 1159
rect 223 1107 227 1159
rect 227 1107 279 1159
rect 349 1107 359 1159
rect 359 1107 387 1159
rect 387 1107 405 1159
rect 475 1107 519 1159
rect 519 1107 531 1159
rect 601 1107 627 1159
rect 627 1107 657 1159
rect 727 1107 759 1159
rect 759 1107 783 1159
rect 853 1107 867 1159
rect 867 1107 909 1159
rect 979 1107 999 1159
rect 999 1107 1027 1159
rect 1027 1107 1035 1159
rect 1105 1107 1107 1159
rect 1107 1107 1159 1159
rect 1159 1107 1161 1159
rect 1231 1107 1239 1159
rect 1239 1107 1267 1159
rect 1267 1107 1287 1159
rect 1357 1107 1399 1159
rect 1399 1107 1413 1159
rect 1483 1107 1507 1159
rect 1507 1107 1539 1159
rect 1609 1107 1639 1159
rect 1639 1107 1665 1159
rect 1735 1107 1747 1159
rect 1747 1107 1791 1159
rect 1861 1107 1879 1159
rect 1879 1107 1907 1159
rect 1907 1107 1917 1159
rect 1987 1107 2039 1159
rect 2039 1107 2043 1159
rect 2113 1107 2119 1159
rect 2119 1107 2169 1159
rect 97 1105 153 1107
rect 223 1105 279 1107
rect 349 1105 405 1107
rect 475 1105 531 1107
rect 601 1105 657 1107
rect 727 1105 783 1107
rect 853 1105 909 1107
rect 979 1105 1035 1107
rect 1105 1105 1161 1107
rect 1231 1105 1287 1107
rect 1357 1105 1413 1107
rect 1483 1105 1539 1107
rect 1609 1105 1665 1107
rect 1735 1105 1791 1107
rect 1861 1105 1917 1107
rect 1987 1105 2043 1107
rect 2113 1105 2169 1107
rect 1105 1027 1107 1035
rect 1107 1027 1159 1035
rect 1159 1027 1161 1035
rect 5 988 61 1016
rect 5 960 7 988
rect 7 960 59 988
rect 59 960 61 988
rect 1105 999 1161 1027
rect 1105 979 1107 999
rect 1107 979 1159 999
rect 1159 979 1161 999
rect 2205 988 2261 1016
rect 2205 960 2207 988
rect 2207 960 2259 988
rect 2259 960 2261 988
rect 5 856 7 890
rect 7 856 59 890
rect 59 856 61 890
rect 5 834 61 856
rect 1105 867 1107 909
rect 1107 867 1159 909
rect 1159 867 1161 909
rect 1105 853 1161 867
rect 2205 856 2207 890
rect 2207 856 2259 890
rect 2259 856 2261 890
rect 2205 834 2261 856
rect 5 748 61 764
rect 5 708 7 748
rect 7 708 59 748
rect 59 708 61 748
rect 1105 759 1161 783
rect 1105 727 1107 759
rect 1107 727 1159 759
rect 1159 727 1161 759
rect 2205 748 2261 764
rect 2205 708 2207 748
rect 2207 708 2259 748
rect 2259 708 2261 748
rect 5 616 7 638
rect 7 616 59 638
rect 59 616 61 638
rect 5 588 61 616
rect 1105 627 1107 657
rect 1107 627 1159 657
rect 1159 627 1161 657
rect 1105 601 1161 627
rect 5 582 7 588
rect 7 582 59 588
rect 59 582 61 588
rect 2205 616 2207 638
rect 2207 616 2259 638
rect 2259 616 2261 638
rect 2205 588 2261 616
rect 2205 582 2207 588
rect 2207 582 2259 588
rect 2259 582 2261 588
rect 5 508 61 512
rect 5 456 7 508
rect 7 456 59 508
rect 59 456 61 508
rect 1105 519 1161 531
rect 1105 475 1107 519
rect 1107 475 1159 519
rect 1159 475 1161 519
rect 2205 508 2261 512
rect 2205 456 2207 508
rect 2207 456 2259 508
rect 2259 456 2261 508
rect 5 376 7 386
rect 7 376 59 386
rect 59 376 61 386
rect 5 348 61 376
rect 5 330 7 348
rect 7 330 59 348
rect 59 330 61 348
rect 1105 387 1107 405
rect 1107 387 1159 405
rect 1159 387 1161 405
rect 1105 359 1161 387
rect 1105 349 1107 359
rect 1107 349 1159 359
rect 1159 349 1161 359
rect 2205 376 2207 386
rect 2207 376 2259 386
rect 2259 376 2261 386
rect 2205 348 2261 376
rect 2205 330 2207 348
rect 2207 330 2259 348
rect 2259 330 2261 348
rect 5 216 7 260
rect 7 216 59 260
rect 59 216 61 260
rect 5 204 61 216
rect 1105 227 1107 279
rect 1107 227 1159 279
rect 1159 227 1161 279
rect 1105 223 1161 227
rect 2205 216 2207 260
rect 2207 216 2259 260
rect 2259 216 2261 260
rect 2205 204 2261 216
rect 5 78 61 134
rect 1105 147 1107 153
rect 1107 147 1159 153
rect 1159 147 1161 153
rect 1105 97 1161 147
rect 2205 78 2261 134
rect 78 59 134 61
rect 204 59 260 61
rect 330 59 386 61
rect 456 59 512 61
rect 582 59 638 61
rect 708 59 764 61
rect 834 59 890 61
rect 960 59 1016 61
rect 78 7 108 59
rect 108 7 134 59
rect 204 7 216 59
rect 216 7 260 59
rect 330 7 348 59
rect 348 7 376 59
rect 376 7 386 59
rect 456 7 508 59
rect 508 7 512 59
rect 582 7 588 59
rect 588 7 616 59
rect 616 7 638 59
rect 708 7 748 59
rect 748 7 764 59
rect 834 7 856 59
rect 856 7 890 59
rect 960 7 988 59
rect 988 7 1016 59
rect 78 5 134 7
rect 204 5 260 7
rect 330 5 386 7
rect 456 5 512 7
rect 582 5 638 7
rect 708 5 764 7
rect 834 5 890 7
rect 960 5 1016 7
rect 1250 59 1306 61
rect 1376 59 1432 61
rect 1502 59 1558 61
rect 1628 59 1684 61
rect 1754 59 1810 61
rect 1880 59 1936 61
rect 2006 59 2062 61
rect 2132 59 2188 61
rect 1250 7 1278 59
rect 1278 7 1306 59
rect 1376 7 1410 59
rect 1410 7 1432 59
rect 1502 7 1518 59
rect 1518 7 1558 59
rect 1628 7 1650 59
rect 1650 7 1678 59
rect 1678 7 1684 59
rect 1754 7 1758 59
rect 1758 7 1810 59
rect 1880 7 1890 59
rect 1890 7 1918 59
rect 1918 7 1936 59
rect 2006 7 2050 59
rect 2050 7 2062 59
rect 2132 7 2158 59
rect 2158 7 2188 59
rect 1250 5 1306 7
rect 1376 5 1432 7
rect 1502 5 1558 7
rect 1628 5 1684 7
rect 1754 5 1810 7
rect 1880 5 1936 7
rect 2006 5 2062 7
rect 2132 5 2188 7
<< metal3 >>
rect 0 2265 1026 2266
rect 0 2201 74 2265
rect 138 2201 200 2265
rect 264 2201 326 2265
rect 390 2201 452 2265
rect 516 2201 578 2265
rect 642 2201 704 2265
rect 768 2201 830 2265
rect 894 2201 956 2265
rect 1020 2201 1026 2265
rect 0 2200 1026 2201
rect 1240 2265 2266 2266
rect 1240 2201 1246 2265
rect 1310 2201 1372 2265
rect 1436 2201 1498 2265
rect 1562 2201 1624 2265
rect 1688 2201 1750 2265
rect 1814 2201 1876 2265
rect 1940 2201 2002 2265
rect 2066 2201 2128 2265
rect 2192 2201 2266 2265
rect 1240 2200 2266 2201
rect 0 2192 66 2200
rect 0 2128 1 2192
rect 65 2128 66 2192
rect 0 2066 66 2128
rect 0 2002 1 2066
rect 65 2002 66 2066
rect 0 1940 66 2002
rect 0 1876 1 1940
rect 65 1876 66 1940
rect 0 1814 66 1876
rect 0 1750 1 1814
rect 65 1750 66 1814
rect 0 1688 66 1750
rect 0 1624 1 1688
rect 65 1624 66 1688
rect 0 1562 66 1624
rect 0 1498 1 1562
rect 65 1498 66 1562
rect 0 1436 66 1498
rect 0 1372 1 1436
rect 65 1372 66 1436
rect 0 1310 66 1372
rect 0 1246 1 1310
rect 65 1246 66 1310
rect 0 1240 66 1246
rect 126 1180 186 2140
rect 246 1240 306 2200
rect 366 1180 426 2140
rect 486 1240 546 2200
rect 606 1180 666 2140
rect 726 1240 786 2200
rect 846 1180 906 2140
rect 966 1240 1026 2200
rect 1086 2169 1180 2200
rect 1086 2113 1105 2169
rect 1161 2113 1180 2169
rect 1086 2047 1180 2113
rect 1086 1983 1101 2047
rect 1165 1983 1180 2047
rect 1086 1921 1180 1983
rect 1086 1857 1101 1921
rect 1165 1857 1180 1921
rect 1086 1795 1180 1857
rect 1086 1731 1101 1795
rect 1165 1731 1180 1795
rect 1086 1669 1180 1731
rect 1086 1605 1101 1669
rect 1165 1605 1180 1669
rect 1086 1543 1180 1605
rect 1086 1479 1101 1543
rect 1165 1479 1180 1543
rect 1086 1417 1180 1479
rect 1086 1353 1101 1417
rect 1165 1353 1180 1417
rect 1086 1291 1180 1353
rect 1086 1227 1101 1291
rect 1165 1227 1180 1291
rect 1240 1240 1300 2200
rect 1086 1180 1180 1227
rect 1360 1180 1420 2140
rect 1480 1240 1540 2200
rect 1600 1180 1660 2140
rect 1720 1240 1780 2200
rect 1840 1180 1900 2140
rect 1960 1240 2020 2200
rect 2200 2192 2266 2200
rect 2080 1180 2140 2140
rect 2200 2128 2201 2192
rect 2265 2128 2266 2192
rect 2200 2066 2266 2128
rect 2200 2002 2201 2066
rect 2265 2002 2266 2066
rect 2200 1940 2266 2002
rect 2200 1876 2201 1940
rect 2265 1876 2266 1940
rect 2200 1814 2266 1876
rect 2200 1750 2201 1814
rect 2265 1750 2266 1814
rect 2200 1688 2266 1750
rect 2200 1624 2201 1688
rect 2265 1624 2266 1688
rect 2200 1562 2266 1624
rect 2200 1498 2201 1562
rect 2265 1498 2266 1562
rect 2200 1436 2266 1498
rect 2200 1372 2201 1436
rect 2265 1372 2266 1436
rect 2200 1310 2266 1372
rect 2200 1246 2201 1310
rect 2265 1246 2266 1310
rect 2200 1240 2266 1246
rect 66 1165 2200 1180
rect 66 1161 219 1165
rect 66 1105 97 1161
rect 153 1105 219 1161
rect 66 1101 219 1105
rect 283 1101 345 1165
rect 409 1101 471 1165
rect 535 1101 597 1165
rect 661 1101 723 1165
rect 787 1101 849 1165
rect 913 1101 975 1165
rect 1039 1101 1101 1165
rect 1165 1101 1227 1165
rect 1291 1101 1353 1165
rect 1417 1101 1479 1165
rect 1543 1101 1605 1165
rect 1669 1101 1731 1165
rect 1795 1101 1857 1165
rect 1921 1101 1983 1165
rect 2047 1161 2200 1165
rect 2047 1105 2113 1161
rect 2169 1105 2200 1161
rect 2047 1101 2200 1105
rect 66 1086 2200 1101
rect 0 1020 66 1026
rect 0 956 1 1020
rect 65 956 66 1020
rect 0 894 66 956
rect 0 830 1 894
rect 65 830 66 894
rect 0 768 66 830
rect 0 704 1 768
rect 65 704 66 768
rect 0 642 66 704
rect 0 578 1 642
rect 65 578 66 642
rect 0 516 66 578
rect 0 452 1 516
rect 65 452 66 516
rect 0 390 66 452
rect 0 326 1 390
rect 65 326 66 390
rect 0 264 66 326
rect 0 200 1 264
rect 65 200 66 264
rect 0 138 66 200
rect 0 74 1 138
rect 65 74 66 138
rect 126 126 186 1086
rect 0 66 66 74
rect 246 66 306 1026
rect 366 126 426 1086
rect 486 66 546 1026
rect 606 126 666 1086
rect 726 66 786 1026
rect 846 126 906 1086
rect 1086 1039 1180 1086
rect 966 66 1026 1026
rect 1086 975 1101 1039
rect 1165 975 1180 1039
rect 1086 913 1180 975
rect 1086 849 1101 913
rect 1165 849 1180 913
rect 1086 787 1180 849
rect 1086 723 1101 787
rect 1165 723 1180 787
rect 1086 661 1180 723
rect 1086 597 1101 661
rect 1165 597 1180 661
rect 1086 535 1180 597
rect 1086 471 1101 535
rect 1165 471 1180 535
rect 1086 409 1180 471
rect 1086 345 1101 409
rect 1165 345 1180 409
rect 1086 283 1180 345
rect 1086 219 1101 283
rect 1165 219 1180 283
rect 1086 153 1180 219
rect 1086 97 1105 153
rect 1161 97 1180 153
rect 1086 66 1180 97
rect 1240 66 1300 1026
rect 1360 126 1420 1086
rect 1480 66 1540 1026
rect 1600 126 1660 1086
rect 1720 66 1780 1026
rect 1840 126 1900 1086
rect 1960 66 2020 1026
rect 2080 126 2140 1086
rect 2200 1020 2266 1026
rect 2200 956 2201 1020
rect 2265 956 2266 1020
rect 2200 894 2266 956
rect 2200 830 2201 894
rect 2265 830 2266 894
rect 2200 768 2266 830
rect 2200 704 2201 768
rect 2265 704 2266 768
rect 2200 642 2266 704
rect 2200 578 2201 642
rect 2265 578 2266 642
rect 2200 516 2266 578
rect 2200 452 2201 516
rect 2265 452 2266 516
rect 2200 390 2266 452
rect 2200 326 2201 390
rect 2265 326 2266 390
rect 2200 264 2266 326
rect 2200 200 2201 264
rect 2265 200 2266 264
rect 2200 138 2266 200
rect 2200 74 2201 138
rect 2265 74 2266 138
rect 2200 66 2266 74
rect 0 65 1026 66
rect 0 1 74 65
rect 138 1 200 65
rect 264 1 326 65
rect 390 1 452 65
rect 516 1 578 65
rect 642 1 704 65
rect 768 1 830 65
rect 894 1 956 65
rect 1020 1 1026 65
rect 0 0 1026 1
rect 1240 65 2266 66
rect 1240 1 1246 65
rect 1310 1 1372 65
rect 1436 1 1498 65
rect 1562 1 1624 65
rect 1688 1 1750 65
rect 1814 1 1876 65
rect 1940 1 2002 65
rect 2066 1 2128 65
rect 2192 1 2266 65
rect 1240 0 2266 1
<< via3 >>
rect 74 2261 138 2265
rect 74 2205 78 2261
rect 78 2205 134 2261
rect 134 2205 138 2261
rect 74 2201 138 2205
rect 200 2261 264 2265
rect 200 2205 204 2261
rect 204 2205 260 2261
rect 260 2205 264 2261
rect 200 2201 264 2205
rect 326 2261 390 2265
rect 326 2205 330 2261
rect 330 2205 386 2261
rect 386 2205 390 2261
rect 326 2201 390 2205
rect 452 2261 516 2265
rect 452 2205 456 2261
rect 456 2205 512 2261
rect 512 2205 516 2261
rect 452 2201 516 2205
rect 578 2261 642 2265
rect 578 2205 582 2261
rect 582 2205 638 2261
rect 638 2205 642 2261
rect 578 2201 642 2205
rect 704 2261 768 2265
rect 704 2205 708 2261
rect 708 2205 764 2261
rect 764 2205 768 2261
rect 704 2201 768 2205
rect 830 2261 894 2265
rect 830 2205 834 2261
rect 834 2205 890 2261
rect 890 2205 894 2261
rect 830 2201 894 2205
rect 956 2261 1020 2265
rect 956 2205 960 2261
rect 960 2205 1016 2261
rect 1016 2205 1020 2261
rect 956 2201 1020 2205
rect 1246 2261 1310 2265
rect 1246 2205 1250 2261
rect 1250 2205 1306 2261
rect 1306 2205 1310 2261
rect 1246 2201 1310 2205
rect 1372 2261 1436 2265
rect 1372 2205 1376 2261
rect 1376 2205 1432 2261
rect 1432 2205 1436 2261
rect 1372 2201 1436 2205
rect 1498 2261 1562 2265
rect 1498 2205 1502 2261
rect 1502 2205 1558 2261
rect 1558 2205 1562 2261
rect 1498 2201 1562 2205
rect 1624 2261 1688 2265
rect 1624 2205 1628 2261
rect 1628 2205 1684 2261
rect 1684 2205 1688 2261
rect 1624 2201 1688 2205
rect 1750 2261 1814 2265
rect 1750 2205 1754 2261
rect 1754 2205 1810 2261
rect 1810 2205 1814 2261
rect 1750 2201 1814 2205
rect 1876 2261 1940 2265
rect 1876 2205 1880 2261
rect 1880 2205 1936 2261
rect 1936 2205 1940 2261
rect 1876 2201 1940 2205
rect 2002 2261 2066 2265
rect 2002 2205 2006 2261
rect 2006 2205 2062 2261
rect 2062 2205 2066 2261
rect 2002 2201 2066 2205
rect 2128 2261 2192 2265
rect 2128 2205 2132 2261
rect 2132 2205 2188 2261
rect 2188 2205 2192 2261
rect 2128 2201 2192 2205
rect 1 2188 65 2192
rect 1 2132 5 2188
rect 5 2132 61 2188
rect 61 2132 65 2188
rect 1 2128 65 2132
rect 1 2062 65 2066
rect 1 2006 5 2062
rect 5 2006 61 2062
rect 61 2006 65 2062
rect 1 2002 65 2006
rect 1 1936 65 1940
rect 1 1880 5 1936
rect 5 1880 61 1936
rect 61 1880 65 1936
rect 1 1876 65 1880
rect 1 1810 65 1814
rect 1 1754 5 1810
rect 5 1754 61 1810
rect 61 1754 65 1810
rect 1 1750 65 1754
rect 1 1684 65 1688
rect 1 1628 5 1684
rect 5 1628 61 1684
rect 61 1628 65 1684
rect 1 1624 65 1628
rect 1 1558 65 1562
rect 1 1502 5 1558
rect 5 1502 61 1558
rect 61 1502 65 1558
rect 1 1498 65 1502
rect 1 1432 65 1436
rect 1 1376 5 1432
rect 5 1376 61 1432
rect 61 1376 65 1432
rect 1 1372 65 1376
rect 1 1306 65 1310
rect 1 1250 5 1306
rect 5 1250 61 1306
rect 61 1250 65 1306
rect 1 1246 65 1250
rect 1101 2043 1165 2047
rect 1101 1987 1105 2043
rect 1105 1987 1161 2043
rect 1161 1987 1165 2043
rect 1101 1983 1165 1987
rect 1101 1917 1165 1921
rect 1101 1861 1105 1917
rect 1105 1861 1161 1917
rect 1161 1861 1165 1917
rect 1101 1857 1165 1861
rect 1101 1791 1165 1795
rect 1101 1735 1105 1791
rect 1105 1735 1161 1791
rect 1161 1735 1165 1791
rect 1101 1731 1165 1735
rect 1101 1665 1165 1669
rect 1101 1609 1105 1665
rect 1105 1609 1161 1665
rect 1161 1609 1165 1665
rect 1101 1605 1165 1609
rect 1101 1539 1165 1543
rect 1101 1483 1105 1539
rect 1105 1483 1161 1539
rect 1161 1483 1165 1539
rect 1101 1479 1165 1483
rect 1101 1413 1165 1417
rect 1101 1357 1105 1413
rect 1105 1357 1161 1413
rect 1161 1357 1165 1413
rect 1101 1353 1165 1357
rect 1101 1287 1165 1291
rect 1101 1231 1105 1287
rect 1105 1231 1161 1287
rect 1161 1231 1165 1287
rect 1101 1227 1165 1231
rect 2201 2188 2265 2192
rect 2201 2132 2205 2188
rect 2205 2132 2261 2188
rect 2261 2132 2265 2188
rect 2201 2128 2265 2132
rect 2201 2062 2265 2066
rect 2201 2006 2205 2062
rect 2205 2006 2261 2062
rect 2261 2006 2265 2062
rect 2201 2002 2265 2006
rect 2201 1936 2265 1940
rect 2201 1880 2205 1936
rect 2205 1880 2261 1936
rect 2261 1880 2265 1936
rect 2201 1876 2265 1880
rect 2201 1810 2265 1814
rect 2201 1754 2205 1810
rect 2205 1754 2261 1810
rect 2261 1754 2265 1810
rect 2201 1750 2265 1754
rect 2201 1684 2265 1688
rect 2201 1628 2205 1684
rect 2205 1628 2261 1684
rect 2261 1628 2265 1684
rect 2201 1624 2265 1628
rect 2201 1558 2265 1562
rect 2201 1502 2205 1558
rect 2205 1502 2261 1558
rect 2261 1502 2265 1558
rect 2201 1498 2265 1502
rect 2201 1432 2265 1436
rect 2201 1376 2205 1432
rect 2205 1376 2261 1432
rect 2261 1376 2265 1432
rect 2201 1372 2265 1376
rect 2201 1306 2265 1310
rect 2201 1250 2205 1306
rect 2205 1250 2261 1306
rect 2261 1250 2265 1306
rect 2201 1246 2265 1250
rect 219 1161 283 1165
rect 219 1105 223 1161
rect 223 1105 279 1161
rect 279 1105 283 1161
rect 219 1101 283 1105
rect 345 1161 409 1165
rect 345 1105 349 1161
rect 349 1105 405 1161
rect 405 1105 409 1161
rect 345 1101 409 1105
rect 471 1161 535 1165
rect 471 1105 475 1161
rect 475 1105 531 1161
rect 531 1105 535 1161
rect 471 1101 535 1105
rect 597 1161 661 1165
rect 597 1105 601 1161
rect 601 1105 657 1161
rect 657 1105 661 1161
rect 597 1101 661 1105
rect 723 1161 787 1165
rect 723 1105 727 1161
rect 727 1105 783 1161
rect 783 1105 787 1161
rect 723 1101 787 1105
rect 849 1161 913 1165
rect 849 1105 853 1161
rect 853 1105 909 1161
rect 909 1105 913 1161
rect 849 1101 913 1105
rect 975 1161 1039 1165
rect 975 1105 979 1161
rect 979 1105 1035 1161
rect 1035 1105 1039 1161
rect 975 1101 1039 1105
rect 1101 1161 1165 1165
rect 1101 1105 1105 1161
rect 1105 1105 1161 1161
rect 1161 1105 1165 1161
rect 1101 1101 1165 1105
rect 1227 1161 1291 1165
rect 1227 1105 1231 1161
rect 1231 1105 1287 1161
rect 1287 1105 1291 1161
rect 1227 1101 1291 1105
rect 1353 1161 1417 1165
rect 1353 1105 1357 1161
rect 1357 1105 1413 1161
rect 1413 1105 1417 1161
rect 1353 1101 1417 1105
rect 1479 1161 1543 1165
rect 1479 1105 1483 1161
rect 1483 1105 1539 1161
rect 1539 1105 1543 1161
rect 1479 1101 1543 1105
rect 1605 1161 1669 1165
rect 1605 1105 1609 1161
rect 1609 1105 1665 1161
rect 1665 1105 1669 1161
rect 1605 1101 1669 1105
rect 1731 1161 1795 1165
rect 1731 1105 1735 1161
rect 1735 1105 1791 1161
rect 1791 1105 1795 1161
rect 1731 1101 1795 1105
rect 1857 1161 1921 1165
rect 1857 1105 1861 1161
rect 1861 1105 1917 1161
rect 1917 1105 1921 1161
rect 1857 1101 1921 1105
rect 1983 1161 2047 1165
rect 1983 1105 1987 1161
rect 1987 1105 2043 1161
rect 2043 1105 2047 1161
rect 1983 1101 2047 1105
rect 1 1016 65 1020
rect 1 960 5 1016
rect 5 960 61 1016
rect 61 960 65 1016
rect 1 956 65 960
rect 1 890 65 894
rect 1 834 5 890
rect 5 834 61 890
rect 61 834 65 890
rect 1 830 65 834
rect 1 764 65 768
rect 1 708 5 764
rect 5 708 61 764
rect 61 708 65 764
rect 1 704 65 708
rect 1 638 65 642
rect 1 582 5 638
rect 5 582 61 638
rect 61 582 65 638
rect 1 578 65 582
rect 1 512 65 516
rect 1 456 5 512
rect 5 456 61 512
rect 61 456 65 512
rect 1 452 65 456
rect 1 386 65 390
rect 1 330 5 386
rect 5 330 61 386
rect 61 330 65 386
rect 1 326 65 330
rect 1 260 65 264
rect 1 204 5 260
rect 5 204 61 260
rect 61 204 65 260
rect 1 200 65 204
rect 1 134 65 138
rect 1 78 5 134
rect 5 78 61 134
rect 61 78 65 134
rect 1 74 65 78
rect 1101 1035 1165 1039
rect 1101 979 1105 1035
rect 1105 979 1161 1035
rect 1161 979 1165 1035
rect 1101 975 1165 979
rect 1101 909 1165 913
rect 1101 853 1105 909
rect 1105 853 1161 909
rect 1161 853 1165 909
rect 1101 849 1165 853
rect 1101 783 1165 787
rect 1101 727 1105 783
rect 1105 727 1161 783
rect 1161 727 1165 783
rect 1101 723 1165 727
rect 1101 657 1165 661
rect 1101 601 1105 657
rect 1105 601 1161 657
rect 1161 601 1165 657
rect 1101 597 1165 601
rect 1101 531 1165 535
rect 1101 475 1105 531
rect 1105 475 1161 531
rect 1161 475 1165 531
rect 1101 471 1165 475
rect 1101 405 1165 409
rect 1101 349 1105 405
rect 1105 349 1161 405
rect 1161 349 1165 405
rect 1101 345 1165 349
rect 1101 279 1165 283
rect 1101 223 1105 279
rect 1105 223 1161 279
rect 1161 223 1165 279
rect 1101 219 1165 223
rect 2201 1016 2265 1020
rect 2201 960 2205 1016
rect 2205 960 2261 1016
rect 2261 960 2265 1016
rect 2201 956 2265 960
rect 2201 890 2265 894
rect 2201 834 2205 890
rect 2205 834 2261 890
rect 2261 834 2265 890
rect 2201 830 2265 834
rect 2201 764 2265 768
rect 2201 708 2205 764
rect 2205 708 2261 764
rect 2261 708 2265 764
rect 2201 704 2265 708
rect 2201 638 2265 642
rect 2201 582 2205 638
rect 2205 582 2261 638
rect 2261 582 2265 638
rect 2201 578 2265 582
rect 2201 512 2265 516
rect 2201 456 2205 512
rect 2205 456 2261 512
rect 2261 456 2265 512
rect 2201 452 2265 456
rect 2201 386 2265 390
rect 2201 330 2205 386
rect 2205 330 2261 386
rect 2261 330 2265 386
rect 2201 326 2265 330
rect 2201 260 2265 264
rect 2201 204 2205 260
rect 2205 204 2261 260
rect 2261 204 2265 260
rect 2201 200 2265 204
rect 2201 134 2265 138
rect 2201 78 2205 134
rect 2205 78 2261 134
rect 2261 78 2265 134
rect 2201 74 2265 78
rect 74 61 138 65
rect 74 5 78 61
rect 78 5 134 61
rect 134 5 138 61
rect 74 1 138 5
rect 200 61 264 65
rect 200 5 204 61
rect 204 5 260 61
rect 260 5 264 61
rect 200 1 264 5
rect 326 61 390 65
rect 326 5 330 61
rect 330 5 386 61
rect 386 5 390 61
rect 326 1 390 5
rect 452 61 516 65
rect 452 5 456 61
rect 456 5 512 61
rect 512 5 516 61
rect 452 1 516 5
rect 578 61 642 65
rect 578 5 582 61
rect 582 5 638 61
rect 638 5 642 61
rect 578 1 642 5
rect 704 61 768 65
rect 704 5 708 61
rect 708 5 764 61
rect 764 5 768 61
rect 704 1 768 5
rect 830 61 894 65
rect 830 5 834 61
rect 834 5 890 61
rect 890 5 894 61
rect 830 1 894 5
rect 956 61 1020 65
rect 956 5 960 61
rect 960 5 1016 61
rect 1016 5 1020 61
rect 956 1 1020 5
rect 1246 61 1310 65
rect 1246 5 1250 61
rect 1250 5 1306 61
rect 1306 5 1310 61
rect 1246 1 1310 5
rect 1372 61 1436 65
rect 1372 5 1376 61
rect 1376 5 1432 61
rect 1432 5 1436 61
rect 1372 1 1436 5
rect 1498 61 1562 65
rect 1498 5 1502 61
rect 1502 5 1558 61
rect 1558 5 1562 61
rect 1498 1 1562 5
rect 1624 61 1688 65
rect 1624 5 1628 61
rect 1628 5 1684 61
rect 1684 5 1688 61
rect 1624 1 1688 5
rect 1750 61 1814 65
rect 1750 5 1754 61
rect 1754 5 1810 61
rect 1810 5 1814 61
rect 1750 1 1814 5
rect 1876 61 1940 65
rect 1876 5 1880 61
rect 1880 5 1936 61
rect 1936 5 1940 61
rect 1876 1 1940 5
rect 2002 61 2066 65
rect 2002 5 2006 61
rect 2006 5 2062 61
rect 2062 5 2066 61
rect 2002 1 2066 5
rect 2128 61 2192 65
rect 2128 5 2132 61
rect 2132 5 2188 61
rect 2188 5 2192 61
rect 2128 1 2192 5
<< metal4 >>
rect 0 2265 2266 2266
rect 0 2201 74 2265
rect 138 2201 200 2265
rect 264 2201 326 2265
rect 390 2201 452 2265
rect 516 2201 578 2265
rect 642 2201 704 2265
rect 768 2201 830 2265
rect 894 2201 956 2265
rect 1020 2201 1246 2265
rect 1310 2201 1372 2265
rect 1436 2201 1498 2265
rect 1562 2201 1624 2265
rect 1688 2201 1750 2265
rect 1814 2201 1876 2265
rect 1940 2201 2002 2265
rect 2066 2201 2128 2265
rect 2192 2201 2266 2265
rect 0 2200 2266 2201
rect 0 2192 66 2200
rect 0 2128 1 2192
rect 65 2128 66 2192
rect 2200 2192 2266 2200
rect 0 2066 66 2128
rect 126 2080 2140 2140
rect 2200 2128 2201 2192
rect 2265 2128 2266 2192
rect 0 2002 1 2066
rect 65 2020 66 2066
rect 1086 2047 1180 2080
rect 65 2002 1026 2020
rect 0 1960 1026 2002
rect 1086 1983 1101 2047
rect 1165 1983 1180 2047
rect 2200 2066 2266 2128
rect 2200 2020 2201 2066
rect 0 1940 66 1960
rect 0 1876 1 1940
rect 65 1876 66 1940
rect 1086 1921 1180 1983
rect 1240 2002 2201 2020
rect 2265 2002 2266 2066
rect 1240 1960 2266 2002
rect 1086 1900 1101 1921
rect 0 1814 66 1876
rect 126 1857 1101 1900
rect 1165 1900 1180 1921
rect 2200 1940 2266 1960
rect 1165 1857 2140 1900
rect 126 1840 2140 1857
rect 2200 1876 2201 1940
rect 2265 1876 2266 1940
rect 0 1750 1 1814
rect 65 1780 66 1814
rect 1086 1795 1180 1840
rect 65 1750 1026 1780
rect 0 1720 1026 1750
rect 1086 1731 1101 1795
rect 1165 1731 1180 1795
rect 2200 1814 2266 1876
rect 2200 1780 2201 1814
rect 0 1688 66 1720
rect 0 1624 1 1688
rect 65 1624 66 1688
rect 1086 1669 1180 1731
rect 1240 1750 2201 1780
rect 2265 1750 2266 1814
rect 1240 1720 2266 1750
rect 1086 1660 1101 1669
rect 0 1562 66 1624
rect 126 1605 1101 1660
rect 1165 1660 1180 1669
rect 2200 1688 2266 1720
rect 1165 1605 2140 1660
rect 126 1600 2140 1605
rect 2200 1624 2201 1688
rect 2265 1624 2266 1688
rect 0 1498 1 1562
rect 65 1540 66 1562
rect 1086 1543 1180 1600
rect 65 1498 1026 1540
rect 0 1480 1026 1498
rect 0 1436 66 1480
rect 0 1372 1 1436
rect 65 1372 66 1436
rect 1086 1479 1101 1543
rect 1165 1479 1180 1543
rect 2200 1562 2266 1624
rect 2200 1540 2201 1562
rect 1240 1498 2201 1540
rect 2265 1498 2266 1562
rect 1240 1480 2266 1498
rect 1086 1420 1180 1479
rect 2200 1436 2266 1480
rect 0 1310 66 1372
rect 126 1417 2140 1420
rect 126 1360 1101 1417
rect 0 1246 1 1310
rect 65 1300 66 1310
rect 1086 1353 1101 1360
rect 1165 1360 2140 1417
rect 2200 1372 2201 1436
rect 2265 1372 2266 1436
rect 1165 1353 1180 1360
rect 65 1246 1026 1300
rect 0 1240 1026 1246
rect 1086 1291 1180 1353
rect 2200 1310 2266 1372
rect 2200 1300 2201 1310
rect 0 1026 66 1240
rect 1086 1227 1101 1291
rect 1165 1227 1180 1291
rect 1240 1246 2201 1300
rect 2265 1246 2266 1310
rect 1240 1240 2266 1246
rect 1086 1180 1180 1227
rect 126 1165 2140 1180
rect 126 1101 219 1165
rect 283 1101 345 1165
rect 409 1101 471 1165
rect 535 1101 597 1165
rect 661 1101 723 1165
rect 787 1101 849 1165
rect 913 1101 975 1165
rect 1039 1101 1101 1165
rect 1165 1101 1227 1165
rect 1291 1101 1353 1165
rect 1417 1101 1479 1165
rect 1543 1101 1605 1165
rect 1669 1101 1731 1165
rect 1795 1101 1857 1165
rect 1921 1101 1983 1165
rect 2047 1101 2140 1165
rect 126 1086 2140 1101
rect 1086 1039 1180 1086
rect 0 1020 1026 1026
rect 0 956 1 1020
rect 65 966 1026 1020
rect 1086 975 1101 1039
rect 1165 975 1180 1039
rect 2200 1026 2266 1240
rect 65 956 66 966
rect 0 894 66 956
rect 1086 913 1180 975
rect 1240 1020 2266 1026
rect 1240 966 2201 1020
rect 1086 906 1101 913
rect 0 830 1 894
rect 65 830 66 894
rect 126 849 1101 906
rect 1165 906 1180 913
rect 2200 956 2201 966
rect 2265 956 2266 1020
rect 1165 849 2140 906
rect 126 846 2140 849
rect 2200 894 2266 956
rect 0 786 66 830
rect 1086 787 1180 846
rect 0 768 1026 786
rect 0 704 1 768
rect 65 726 1026 768
rect 65 704 66 726
rect 0 642 66 704
rect 1086 723 1101 787
rect 1165 723 1180 787
rect 2200 830 2201 894
rect 2265 830 2266 894
rect 2200 786 2266 830
rect 1240 768 2266 786
rect 1240 726 2201 768
rect 1086 666 1180 723
rect 2200 704 2201 726
rect 2265 704 2266 768
rect 0 578 1 642
rect 65 578 66 642
rect 126 661 2140 666
rect 126 606 1101 661
rect 0 546 66 578
rect 1086 597 1101 606
rect 1165 606 2140 661
rect 2200 642 2266 704
rect 1165 597 1180 606
rect 0 516 1026 546
rect 0 452 1 516
rect 65 486 1026 516
rect 1086 535 1180 597
rect 2200 578 2201 642
rect 2265 578 2266 642
rect 2200 546 2266 578
rect 65 452 66 486
rect 0 390 66 452
rect 1086 471 1101 535
rect 1165 471 1180 535
rect 1240 516 2266 546
rect 1240 486 2201 516
rect 1086 426 1180 471
rect 2200 452 2201 486
rect 2265 452 2266 516
rect 0 326 1 390
rect 65 326 66 390
rect 126 409 2140 426
rect 126 366 1101 409
rect 0 306 66 326
rect 1086 345 1101 366
rect 1165 366 2140 409
rect 2200 390 2266 452
rect 1165 345 1180 366
rect 0 264 1026 306
rect 0 200 1 264
rect 65 246 1026 264
rect 1086 283 1180 345
rect 2200 326 2201 390
rect 2265 326 2266 390
rect 2200 306 2266 326
rect 65 200 66 246
rect 0 138 66 200
rect 1086 219 1101 283
rect 1165 219 1180 283
rect 1240 264 2266 306
rect 1240 246 2201 264
rect 1086 186 1180 219
rect 2200 200 2201 246
rect 2265 200 2266 264
rect 0 74 1 138
rect 65 74 66 138
rect 126 126 2140 186
rect 2200 138 2266 200
rect 0 66 66 74
rect 2200 74 2201 138
rect 2265 74 2266 138
rect 2200 66 2266 74
rect 0 65 2266 66
rect 0 1 74 65
rect 138 1 200 65
rect 264 1 326 65
rect 390 1 452 65
rect 516 1 578 65
rect 642 1 704 65
rect 768 1 830 65
rect 894 1 956 65
rect 1020 1 1246 65
rect 1310 1 1372 65
rect 1436 1 1498 65
rect 1562 1 1624 65
rect 1688 1 1750 65
rect 1814 1 1876 65
rect 1940 1 2002 65
rect 2066 1 2128 65
rect 2192 1 2266 65
rect 0 0 2266 1
<< labels >>
flabel metal2 s 1450 1421 1469 1441 0 FreeSans 200 0 0 0 C0
port 1 nsew
flabel metal2 s 1485 1362 1521 1386 0 FreeSans 200 0 0 0 C1
port 2 nsew
flabel pwell s 1551 1747 1572 1796 0 FreeSans 400 0 0 0 SUB
port 3 nsew
<< properties >>
string GDS_END 418054
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 380518
string path 56.250 0.825 0.400 0.825 
string device primitive
<< end >>
