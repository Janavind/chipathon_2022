magic
tech sky130B
magscale 1 2
timestamp 1666199351
use sky130_fd_pr__dfl1__example_55959141808187  sky130_fd_pr__dfl1__example_55959141808187_0
timestamp 1666199351
transform 1 0 -42 0 1 21
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808187  sky130_fd_pr__dfl1__example_55959141808187_1
timestamp 1666199351
transform 1 0 7511 0 1 -327
box 0 0 1 1
<< properties >>
string GDS_END 32657196
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 32656036
<< end >>
