magic
tech sky130A
magscale 1 2
timestamp 1666199351
<< nwell >>
rect -38 261 1786 582
<< pwell >>
rect 1 21 1743 203
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 331 47 361 177
rect 415 47 445 177
rect 499 47 529 177
rect 583 47 613 177
rect 667 47 697 177
rect 855 47 885 177
rect 939 47 969 177
rect 1023 47 1053 177
rect 1107 47 1137 177
rect 1191 47 1221 177
rect 1275 47 1305 177
rect 1359 47 1389 177
rect 1443 47 1473 177
rect 1631 47 1661 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 331 297 361 497
rect 415 297 445 497
rect 499 297 529 497
rect 583 297 613 497
rect 667 297 697 497
rect 855 297 885 497
rect 939 297 969 497
rect 1023 297 1053 497
rect 1107 297 1137 497
rect 1191 297 1221 497
rect 1275 297 1305 497
rect 1359 297 1389 497
rect 1443 297 1473 497
rect 1631 297 1661 497
<< ndiff >>
rect 27 163 79 177
rect 27 129 35 163
rect 69 129 79 163
rect 27 95 79 129
rect 27 61 35 95
rect 69 61 79 95
rect 27 47 79 61
rect 109 163 163 177
rect 109 129 119 163
rect 153 129 163 163
rect 109 95 163 129
rect 109 61 119 95
rect 153 61 163 95
rect 109 47 163 61
rect 193 95 247 177
rect 193 61 203 95
rect 237 61 247 95
rect 193 47 247 61
rect 277 163 331 177
rect 277 129 287 163
rect 321 129 331 163
rect 277 95 331 129
rect 277 61 287 95
rect 321 61 331 95
rect 277 47 331 61
rect 361 95 415 177
rect 361 61 371 95
rect 405 61 415 95
rect 361 47 415 61
rect 445 163 499 177
rect 445 129 455 163
rect 489 129 499 163
rect 445 95 499 129
rect 445 61 455 95
rect 489 61 499 95
rect 445 47 499 61
rect 529 95 583 177
rect 529 61 539 95
rect 573 61 583 95
rect 529 47 583 61
rect 613 163 667 177
rect 613 129 623 163
rect 657 129 667 163
rect 613 95 667 129
rect 613 61 623 95
rect 657 61 667 95
rect 613 47 667 61
rect 697 95 855 177
rect 697 61 707 95
rect 741 61 811 95
rect 845 61 855 95
rect 697 47 855 61
rect 885 163 939 177
rect 885 129 895 163
rect 929 129 939 163
rect 885 95 939 129
rect 885 61 895 95
rect 929 61 939 95
rect 885 47 939 61
rect 969 95 1023 177
rect 969 61 979 95
rect 1013 61 1023 95
rect 969 47 1023 61
rect 1053 163 1107 177
rect 1053 129 1063 163
rect 1097 129 1107 163
rect 1053 95 1107 129
rect 1053 61 1063 95
rect 1097 61 1107 95
rect 1053 47 1107 61
rect 1137 95 1191 177
rect 1137 61 1147 95
rect 1181 61 1191 95
rect 1137 47 1191 61
rect 1221 163 1275 177
rect 1221 129 1231 163
rect 1265 129 1275 163
rect 1221 95 1275 129
rect 1221 61 1231 95
rect 1265 61 1275 95
rect 1221 47 1275 61
rect 1305 95 1359 177
rect 1305 61 1315 95
rect 1349 61 1359 95
rect 1305 47 1359 61
rect 1389 163 1443 177
rect 1389 129 1399 163
rect 1433 129 1443 163
rect 1389 95 1443 129
rect 1389 61 1399 95
rect 1433 61 1443 95
rect 1389 47 1443 61
rect 1473 95 1525 177
rect 1473 61 1483 95
rect 1517 61 1525 95
rect 1473 47 1525 61
rect 1579 163 1631 177
rect 1579 129 1587 163
rect 1621 129 1631 163
rect 1579 95 1631 129
rect 1579 61 1587 95
rect 1621 61 1631 95
rect 1579 47 1631 61
rect 1661 163 1717 177
rect 1661 129 1671 163
rect 1705 129 1717 163
rect 1661 95 1717 129
rect 1661 61 1671 95
rect 1705 61 1717 95
rect 1661 47 1717 61
<< pdiff >>
rect 27 479 79 497
rect 27 445 35 479
rect 69 445 79 479
rect 27 411 79 445
rect 27 377 35 411
rect 69 377 79 411
rect 27 343 79 377
rect 27 309 35 343
rect 69 309 79 343
rect 27 297 79 309
rect 109 477 163 497
rect 109 443 119 477
rect 153 443 163 477
rect 109 409 163 443
rect 109 375 119 409
rect 153 375 163 409
rect 109 297 163 375
rect 193 477 247 497
rect 193 443 203 477
rect 237 443 247 477
rect 193 409 247 443
rect 193 375 203 409
rect 237 375 247 409
rect 193 341 247 375
rect 193 307 203 341
rect 237 307 247 341
rect 193 297 247 307
rect 277 477 331 497
rect 277 443 287 477
rect 321 443 331 477
rect 277 409 331 443
rect 277 375 287 409
rect 321 375 331 409
rect 277 297 331 375
rect 361 477 415 497
rect 361 443 371 477
rect 405 443 415 477
rect 361 409 415 443
rect 361 375 371 409
rect 405 375 415 409
rect 361 341 415 375
rect 361 307 371 341
rect 405 307 415 341
rect 361 297 415 307
rect 445 409 499 497
rect 445 375 455 409
rect 489 375 499 409
rect 445 341 499 375
rect 445 307 455 341
rect 489 307 499 341
rect 445 297 499 307
rect 529 477 583 497
rect 529 443 539 477
rect 573 443 583 477
rect 529 409 583 443
rect 529 375 539 409
rect 573 375 583 409
rect 529 297 583 375
rect 613 409 667 497
rect 613 375 623 409
rect 657 375 667 409
rect 613 341 667 375
rect 613 307 623 341
rect 657 307 667 341
rect 613 297 667 307
rect 697 477 749 497
rect 697 443 707 477
rect 741 443 749 477
rect 697 409 749 443
rect 697 375 707 409
rect 741 375 749 409
rect 697 297 749 375
rect 803 477 855 497
rect 803 443 811 477
rect 845 443 855 477
rect 803 409 855 443
rect 803 375 811 409
rect 845 375 855 409
rect 803 297 855 375
rect 885 409 939 497
rect 885 375 895 409
rect 929 375 939 409
rect 885 341 939 375
rect 885 307 895 341
rect 929 307 939 341
rect 885 297 939 307
rect 969 477 1023 497
rect 969 443 979 477
rect 1013 443 1023 477
rect 969 409 1023 443
rect 969 375 979 409
rect 1013 375 1023 409
rect 969 297 1023 375
rect 1053 409 1107 497
rect 1053 375 1063 409
rect 1097 375 1107 409
rect 1053 341 1107 375
rect 1053 307 1063 341
rect 1097 307 1107 341
rect 1053 297 1107 307
rect 1137 477 1191 497
rect 1137 443 1147 477
rect 1181 443 1191 477
rect 1137 409 1191 443
rect 1137 375 1147 409
rect 1181 375 1191 409
rect 1137 341 1191 375
rect 1137 307 1147 341
rect 1181 307 1191 341
rect 1137 297 1191 307
rect 1221 409 1275 497
rect 1221 375 1231 409
rect 1265 375 1275 409
rect 1221 341 1275 375
rect 1221 307 1231 341
rect 1265 307 1275 341
rect 1221 297 1275 307
rect 1305 477 1359 497
rect 1305 443 1315 477
rect 1349 443 1359 477
rect 1305 409 1359 443
rect 1305 375 1315 409
rect 1349 375 1359 409
rect 1305 297 1359 375
rect 1389 409 1443 497
rect 1389 375 1399 409
rect 1433 375 1443 409
rect 1389 341 1443 375
rect 1389 307 1399 341
rect 1433 307 1443 341
rect 1389 297 1443 307
rect 1473 477 1525 497
rect 1473 443 1483 477
rect 1517 443 1525 477
rect 1473 409 1525 443
rect 1473 375 1483 409
rect 1517 375 1525 409
rect 1473 297 1525 375
rect 1579 479 1631 497
rect 1579 445 1587 479
rect 1621 445 1631 479
rect 1579 411 1631 445
rect 1579 377 1587 411
rect 1621 377 1631 411
rect 1579 343 1631 377
rect 1579 309 1587 343
rect 1621 309 1631 343
rect 1579 297 1631 309
rect 1661 479 1717 497
rect 1661 445 1671 479
rect 1705 445 1717 479
rect 1661 411 1717 445
rect 1661 377 1671 411
rect 1705 377 1717 411
rect 1661 343 1717 377
rect 1661 309 1671 343
rect 1705 309 1717 343
rect 1661 297 1717 309
<< ndiffc >>
rect 35 129 69 163
rect 35 61 69 95
rect 119 129 153 163
rect 119 61 153 95
rect 203 61 237 95
rect 287 129 321 163
rect 287 61 321 95
rect 371 61 405 95
rect 455 129 489 163
rect 455 61 489 95
rect 539 61 573 95
rect 623 129 657 163
rect 623 61 657 95
rect 707 61 741 95
rect 811 61 845 95
rect 895 129 929 163
rect 895 61 929 95
rect 979 61 1013 95
rect 1063 129 1097 163
rect 1063 61 1097 95
rect 1147 61 1181 95
rect 1231 129 1265 163
rect 1231 61 1265 95
rect 1315 61 1349 95
rect 1399 129 1433 163
rect 1399 61 1433 95
rect 1483 61 1517 95
rect 1587 129 1621 163
rect 1587 61 1621 95
rect 1671 129 1705 163
rect 1671 61 1705 95
<< pdiffc >>
rect 35 445 69 479
rect 35 377 69 411
rect 35 309 69 343
rect 119 443 153 477
rect 119 375 153 409
rect 203 443 237 477
rect 203 375 237 409
rect 203 307 237 341
rect 287 443 321 477
rect 287 375 321 409
rect 371 443 405 477
rect 371 375 405 409
rect 371 307 405 341
rect 455 375 489 409
rect 455 307 489 341
rect 539 443 573 477
rect 539 375 573 409
rect 623 375 657 409
rect 623 307 657 341
rect 707 443 741 477
rect 707 375 741 409
rect 811 443 845 477
rect 811 375 845 409
rect 895 375 929 409
rect 895 307 929 341
rect 979 443 1013 477
rect 979 375 1013 409
rect 1063 375 1097 409
rect 1063 307 1097 341
rect 1147 443 1181 477
rect 1147 375 1181 409
rect 1147 307 1181 341
rect 1231 375 1265 409
rect 1231 307 1265 341
rect 1315 443 1349 477
rect 1315 375 1349 409
rect 1399 375 1433 409
rect 1399 307 1433 341
rect 1483 443 1517 477
rect 1483 375 1517 409
rect 1587 445 1621 479
rect 1587 377 1621 411
rect 1587 309 1621 343
rect 1671 445 1705 479
rect 1671 377 1705 411
rect 1671 309 1705 343
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 331 497 361 523
rect 415 497 445 523
rect 499 497 529 523
rect 583 497 613 523
rect 667 497 697 523
rect 855 497 885 523
rect 939 497 969 523
rect 1023 497 1053 523
rect 1107 497 1137 523
rect 1191 497 1221 523
rect 1275 497 1305 523
rect 1359 497 1389 523
rect 1443 497 1473 523
rect 1631 497 1661 523
rect 79 265 109 297
rect 163 265 193 297
rect 247 265 277 297
rect 331 265 361 297
rect 79 249 361 265
rect 79 215 95 249
rect 129 215 163 249
rect 197 215 231 249
rect 265 215 299 249
rect 333 215 361 249
rect 79 199 361 215
rect 79 177 109 199
rect 163 177 193 199
rect 247 177 277 199
rect 331 177 361 199
rect 415 265 445 297
rect 499 265 529 297
rect 583 265 613 297
rect 667 265 697 297
rect 415 249 697 265
rect 415 215 431 249
rect 465 215 499 249
rect 533 215 567 249
rect 601 215 635 249
rect 669 215 697 249
rect 415 199 697 215
rect 415 177 445 199
rect 499 177 529 199
rect 583 177 613 199
rect 667 177 697 199
rect 855 265 885 297
rect 939 265 969 297
rect 1023 265 1053 297
rect 1107 265 1137 297
rect 855 249 1137 265
rect 855 215 871 249
rect 905 215 939 249
rect 973 215 1007 249
rect 1041 215 1075 249
rect 1109 215 1137 249
rect 855 199 1137 215
rect 855 177 885 199
rect 939 177 969 199
rect 1023 177 1053 199
rect 1107 177 1137 199
rect 1191 265 1221 297
rect 1275 265 1305 297
rect 1359 265 1389 297
rect 1443 265 1473 297
rect 1631 265 1661 297
rect 1191 249 1544 265
rect 1191 215 1343 249
rect 1377 215 1411 249
rect 1445 215 1494 249
rect 1528 215 1544 249
rect 1191 199 1544 215
rect 1631 249 1712 265
rect 1631 215 1662 249
rect 1696 215 1712 249
rect 1631 199 1712 215
rect 1191 177 1221 199
rect 1275 177 1305 199
rect 1359 177 1389 199
rect 1443 177 1473 199
rect 1631 177 1661 199
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 331 21 361 47
rect 415 21 445 47
rect 499 21 529 47
rect 583 21 613 47
rect 667 21 697 47
rect 855 21 885 47
rect 939 21 969 47
rect 1023 21 1053 47
rect 1107 21 1137 47
rect 1191 21 1221 47
rect 1275 21 1305 47
rect 1359 21 1389 47
rect 1443 21 1473 47
rect 1631 21 1661 47
<< polycont >>
rect 95 215 129 249
rect 163 215 197 249
rect 231 215 265 249
rect 299 215 333 249
rect 431 215 465 249
rect 499 215 533 249
rect 567 215 601 249
rect 635 215 669 249
rect 871 215 905 249
rect 939 215 973 249
rect 1007 215 1041 249
rect 1075 215 1109 249
rect 1343 215 1377 249
rect 1411 215 1445 249
rect 1494 215 1528 249
rect 1662 215 1696 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 19 479 85 493
rect 19 445 35 479
rect 69 445 85 479
rect 19 411 85 445
rect 19 377 35 411
rect 69 377 85 411
rect 19 343 85 377
rect 119 477 161 527
rect 153 443 161 477
rect 119 409 161 443
rect 153 375 161 409
rect 119 359 161 375
rect 195 477 245 493
rect 195 443 203 477
rect 237 443 245 477
rect 195 409 245 443
rect 195 375 203 409
rect 237 375 245 409
rect 19 309 35 343
rect 69 325 85 343
rect 195 341 245 375
rect 279 477 329 527
rect 279 443 287 477
rect 321 443 329 477
rect 279 409 329 443
rect 279 375 287 409
rect 321 375 329 409
rect 279 359 329 375
rect 363 477 749 493
rect 363 443 371 477
rect 405 459 539 477
rect 405 443 413 459
rect 363 409 413 443
rect 531 443 539 459
rect 573 459 707 477
rect 573 443 581 459
rect 363 375 371 409
rect 405 375 413 409
rect 195 325 203 341
rect 69 309 203 325
rect 19 307 203 309
rect 237 325 245 341
rect 363 341 413 375
rect 363 325 371 341
rect 237 307 371 325
rect 405 307 413 341
rect 19 291 413 307
rect 447 409 497 425
rect 447 375 455 409
rect 489 375 497 409
rect 447 341 497 375
rect 531 409 581 443
rect 699 443 707 459
rect 741 443 749 477
rect 531 375 539 409
rect 573 375 581 409
rect 531 359 581 375
rect 615 409 665 425
rect 615 375 623 409
rect 657 375 665 409
rect 447 307 455 341
rect 489 325 497 341
rect 615 341 665 375
rect 699 409 749 443
rect 699 375 707 409
rect 741 375 749 409
rect 699 359 749 375
rect 803 477 1525 493
rect 803 443 811 477
rect 845 459 979 477
rect 845 443 853 459
rect 803 409 853 443
rect 971 443 979 459
rect 1013 459 1147 477
rect 1013 443 1021 459
rect 803 375 811 409
rect 845 375 853 409
rect 803 359 853 375
rect 887 409 937 425
rect 887 375 895 409
rect 929 375 937 409
rect 615 325 623 341
rect 489 307 623 325
rect 657 325 665 341
rect 887 341 937 375
rect 971 409 1021 443
rect 1139 443 1147 459
rect 1181 459 1315 477
rect 1181 443 1189 459
rect 971 375 979 409
rect 1013 375 1021 409
rect 971 359 1021 375
rect 1055 409 1105 425
rect 1055 375 1063 409
rect 1097 375 1105 409
rect 887 325 895 341
rect 657 307 895 325
rect 929 325 937 341
rect 1055 341 1105 375
rect 1055 325 1063 341
rect 929 307 1063 325
rect 1097 307 1105 341
rect 447 291 1105 307
rect 1139 409 1189 443
rect 1307 443 1315 459
rect 1349 459 1483 477
rect 1349 443 1357 459
rect 1139 375 1147 409
rect 1181 375 1189 409
rect 1139 341 1189 375
rect 1139 307 1147 341
rect 1181 307 1189 341
rect 1139 291 1189 307
rect 1223 409 1273 425
rect 1223 375 1231 409
rect 1265 375 1273 409
rect 1223 341 1273 375
rect 1307 409 1357 443
rect 1475 443 1483 459
rect 1517 443 1525 477
rect 1307 375 1315 409
rect 1349 375 1357 409
rect 1307 359 1357 375
rect 1391 409 1441 425
rect 1391 375 1399 409
rect 1433 375 1441 409
rect 1223 307 1231 341
rect 1265 325 1273 341
rect 1391 341 1441 375
rect 1475 409 1525 443
rect 1475 375 1483 409
rect 1517 375 1525 409
rect 1475 359 1525 375
rect 1570 479 1637 493
rect 1570 445 1587 479
rect 1621 445 1637 479
rect 1570 411 1637 445
rect 1570 377 1587 411
rect 1621 377 1637 411
rect 1391 325 1399 341
rect 1265 307 1399 325
rect 1433 307 1441 341
rect 1570 343 1637 377
rect 1570 325 1587 343
rect 1223 291 1441 307
rect 1494 309 1587 325
rect 1621 309 1637 343
rect 1494 291 1637 309
rect 1671 479 1717 527
rect 1705 445 1717 479
rect 1671 411 1717 445
rect 1705 377 1717 411
rect 1671 343 1717 377
rect 1705 309 1717 343
rect 1671 291 1717 309
rect 79 249 361 257
rect 79 215 95 249
rect 129 215 163 249
rect 197 215 231 249
rect 265 215 299 249
rect 333 215 361 249
rect 415 249 750 257
rect 415 215 431 249
rect 465 215 499 249
rect 533 215 567 249
rect 601 215 635 249
rect 669 215 750 249
rect 797 249 1137 257
rect 797 215 871 249
rect 905 215 939 249
rect 973 215 1007 249
rect 1041 215 1075 249
rect 1109 215 1137 249
rect 1223 181 1293 291
rect 1494 257 1528 291
rect 1327 249 1528 257
rect 1327 215 1343 249
rect 1377 215 1411 249
rect 1445 215 1494 249
rect 1562 249 1731 257
rect 1562 215 1662 249
rect 1696 215 1731 249
rect 1494 181 1528 215
rect 35 163 69 179
rect 35 95 69 129
rect 35 17 69 61
rect 103 163 1449 181
rect 103 129 119 163
rect 153 145 287 163
rect 153 129 169 145
rect 103 95 169 129
rect 271 129 287 145
rect 321 145 455 163
rect 321 129 337 145
rect 103 61 119 95
rect 153 61 169 95
rect 103 51 169 61
rect 203 95 237 111
rect 203 17 237 61
rect 271 95 337 129
rect 439 129 455 145
rect 489 145 623 163
rect 489 129 505 145
rect 271 61 287 95
rect 321 61 337 95
rect 271 51 337 61
rect 371 95 405 111
rect 371 17 405 61
rect 439 95 505 129
rect 607 129 623 145
rect 657 145 895 163
rect 657 129 673 145
rect 439 61 455 95
rect 489 61 505 95
rect 439 51 505 61
rect 539 95 573 111
rect 539 17 573 61
rect 607 95 673 129
rect 879 129 895 145
rect 929 145 1063 163
rect 929 129 945 145
rect 607 61 623 95
rect 657 61 673 95
rect 607 51 673 61
rect 707 95 845 111
rect 741 61 811 95
rect 707 17 845 61
rect 879 95 945 129
rect 1047 129 1063 145
rect 1097 145 1231 163
rect 1097 129 1113 145
rect 879 61 895 95
rect 929 61 945 95
rect 879 51 945 61
rect 979 95 1013 111
rect 979 17 1013 61
rect 1047 95 1113 129
rect 1215 129 1231 145
rect 1265 145 1399 163
rect 1265 129 1281 145
rect 1047 61 1063 95
rect 1097 61 1113 95
rect 1047 51 1113 61
rect 1147 95 1181 111
rect 1147 17 1181 61
rect 1215 95 1281 129
rect 1383 129 1399 145
rect 1433 129 1449 163
rect 1494 163 1637 181
rect 1494 147 1587 163
rect 1215 61 1231 95
rect 1265 61 1281 95
rect 1215 51 1281 61
rect 1315 95 1349 111
rect 1315 17 1349 61
rect 1383 95 1449 129
rect 1562 129 1587 147
rect 1621 129 1637 163
rect 1383 61 1399 95
rect 1433 61 1449 95
rect 1383 51 1449 61
rect 1483 95 1517 111
rect 1483 17 1517 61
rect 1562 95 1637 129
rect 1562 61 1587 95
rect 1621 61 1637 95
rect 1562 51 1637 61
rect 1671 163 1717 181
rect 1705 129 1717 163
rect 1671 95 1717 129
rect 1705 61 1717 95
rect 1671 17 1717 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
<< metal1 >>
rect 0 561 1748 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 0 496 1748 527
rect 0 17 1748 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
rect 0 -48 1748 -17
<< labels >>
flabel locali s 578 221 612 255 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel locali s 210 221 244 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 1686 221 1720 255 0 FreeSans 400 0 0 0 D_N
port 4 nsew signal input
flabel locali s 950 221 984 255 0 FreeSans 400 0 0 0 C
port 3 nsew signal input
flabel locali s 1226 357 1260 391 0 FreeSans 400 0 0 0 Y
port 9 nsew signal output
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 nor4b_4
rlabel metal1 s 0 -48 1748 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1748 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1748 544
string GDS_END 1181110
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1167616
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 8.740 0.000 
<< end >>
