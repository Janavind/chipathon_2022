magic
tech sky130A
magscale 1 2
timestamp 1666199351
<< nwell >>
rect -38 261 2246 582
<< pwell >>
rect 347 21 1863 157
rect 29 -17 63 17
<< locali >>
rect 115 333 166 493
rect 287 333 338 490
rect 465 333 510 493
rect 631 333 682 490
rect 803 333 851 490
rect 981 333 1056 490
rect 1185 333 1235 490
rect 1357 333 1407 490
rect 1529 333 1579 490
rect 1701 333 1751 490
rect 1873 333 1921 490
rect 2045 333 2096 490
rect 115 291 2096 333
rect 465 283 1751 291
rect 465 56 510 283
rect 631 56 682 283
rect 803 56 851 283
rect 981 56 1051 283
rect 1185 56 1235 283
rect 1357 56 1407 283
rect 1529 56 1579 283
rect 1701 56 1751 283
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2208 561
rect 28 299 81 527
rect 200 367 252 527
rect 373 367 424 527
rect 544 367 596 527
rect 717 367 768 527
rect 893 367 944 527
rect 1098 424 1150 527
rect 1098 367 1149 424
rect 1271 367 1322 527
rect 1443 367 1494 527
rect 1615 367 1666 527
rect 1787 367 1838 527
rect 1959 367 2010 527
rect 2130 367 2182 527
rect 69 221 305 255
rect 339 221 397 255
rect 69 179 431 221
rect 371 17 425 122
rect 544 17 597 122
rect 716 17 769 122
rect 893 17 946 122
rect 1098 17 1151 122
rect 1270 17 1315 122
rect 1442 17 1495 122
rect 1614 17 1667 122
rect 1786 221 1869 255
rect 1903 221 1961 255
rect 1995 221 2142 255
rect 1786 179 2142 221
rect 1786 17 1839 122
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2208 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 305 221 339 255
rect 397 221 431 255
rect 1869 221 1903 255
rect 1961 221 1995 255
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
<< metal1 >>
rect 0 561 2208 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2208 561
rect 0 496 2208 527
rect 293 255 443 261
rect 293 221 305 255
rect 339 221 397 255
rect 431 252 443 255
rect 1857 255 2007 261
rect 1857 252 1869 255
rect 431 224 1869 252
rect 431 221 443 224
rect 293 215 443 221
rect 1857 221 1869 224
rect 1903 221 1961 255
rect 1995 221 2007 255
rect 1857 215 2007 221
rect 0 17 2208 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2208 17
rect 0 -48 2208 -17
<< labels >>
rlabel metal1 s 1857 215 2007 224 6 A
port 1 nsew signal input
rlabel metal1 s 293 215 443 224 6 A
port 1 nsew signal input
rlabel metal1 s 293 224 2007 252 6 A
port 1 nsew signal input
rlabel metal1 s 1857 252 2007 261 6 A
port 1 nsew signal input
rlabel metal1 s 293 252 443 261 6 A
port 1 nsew signal input
rlabel metal1 s 0 -48 2208 48 8 VGND
port 2 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 17 8 VNB
port 3 nsew ground bidirectional
rlabel nwell s -38 261 2246 582 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 496 2208 592 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 1701 56 1751 283 6 Y
port 6 nsew signal output
rlabel locali s 1529 56 1579 283 6 Y
port 6 nsew signal output
rlabel locali s 1357 56 1407 283 6 Y
port 6 nsew signal output
rlabel locali s 1185 56 1235 283 6 Y
port 6 nsew signal output
rlabel locali s 981 56 1051 283 6 Y
port 6 nsew signal output
rlabel locali s 803 56 851 283 6 Y
port 6 nsew signal output
rlabel locali s 631 56 682 283 6 Y
port 6 nsew signal output
rlabel locali s 465 56 510 283 6 Y
port 6 nsew signal output
rlabel locali s 465 283 1751 291 6 Y
port 6 nsew signal output
rlabel locali s 115 291 2096 333 6 Y
port 6 nsew signal output
rlabel locali s 2045 333 2096 490 6 Y
port 6 nsew signal output
rlabel locali s 1873 333 1921 490 6 Y
port 6 nsew signal output
rlabel locali s 1701 333 1751 490 6 Y
port 6 nsew signal output
rlabel locali s 1529 333 1579 490 6 Y
port 6 nsew signal output
rlabel locali s 1357 333 1407 490 6 Y
port 6 nsew signal output
rlabel locali s 1185 333 1235 490 6 Y
port 6 nsew signal output
rlabel locali s 981 333 1056 490 6 Y
port 6 nsew signal output
rlabel locali s 803 333 851 490 6 Y
port 6 nsew signal output
rlabel locali s 631 333 682 490 6 Y
port 6 nsew signal output
rlabel locali s 465 333 510 493 6 Y
port 6 nsew signal output
rlabel locali s 287 333 338 490 6 Y
port 6 nsew signal output
rlabel locali s 115 333 166 493 6 Y
port 6 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2208 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3349990
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3337002
<< end >>
