magic
tech sky130B
magscale 1 2
timestamp 1666464484
use sky130_fd_pr__hvdfl1sd2__example_55959141808178  sky130_fd_pr__hvdfl1sd2__example_55959141808178_0
timestamp 1666464484
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808178  sky130_fd_pr__hvdfl1sd2__example_55959141808178_1
timestamp 1666464484
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808178  sky130_fd_pr__hvdfl1sd2__example_55959141808178_2
timestamp 1666464484
transform 1 0 256 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808178  sky130_fd_pr__hvdfl1sd2__example_55959141808178_3
timestamp 1666464484
transform 1 0 412 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808178  sky130_fd_pr__hvdfl1sd2__example_55959141808178_4
timestamp 1666464484
transform 1 0 568 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808178  sky130_fd_pr__hvdfl1sd2__example_55959141808178_5
timestamp 1666464484
transform 1 0 724 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808178  sky130_fd_pr__hvdfl1sd2__example_55959141808178_6
timestamp 1666464484
transform 1 0 880 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808178  sky130_fd_pr__hvdfl1sd2__example_55959141808178_7
timestamp 1666464484
transform 1 0 1036 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 43513828
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 43509662
<< end >>
