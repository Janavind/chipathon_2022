magic
tech sky130A
timestamp 1666464484
<< properties >>
string GDS_END 3298718
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 3297950
<< end >>
