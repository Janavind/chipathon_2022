magic
tech sky130A
magscale 1 2
timestamp 1666464484
use sky130_fd_pr__hvdftpl1s__example_55959141808646  sky130_fd_pr__hvdftpl1s__example_55959141808646_0
timestamp 1666464484
transform -1 0 -77 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 1500774
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 1499916
<< end >>
