magic
tech sky130A
magscale 1 2
timestamp 1666464484
<< locali >>
rect 0 1397 846 1431
rect 430 686 464 1167
rect 430 652 559 686
rect 657 652 691 686
rect 345 485 379 551
rect 212 361 246 427
rect 79 237 113 303
rect 0 -17 846 17
use sky130_sram_1kbyte_1rw1r_8x1024_8_pdriver_0  sky130_sram_1kbyte_1rw1r_8x1024_8_pdriver_0_0
timestamp 1666464484
transform 1 0 478 0 1 0
box -36 -17 404 1471
use sky130_sram_1kbyte_1rw1r_8x1024_8_pnand3  sky130_sram_1kbyte_1rw1r_8x1024_8_pnand3_0
timestamp 1666464484
transform 1 0 0 0 1 0
box -36 -17 514 1471
<< labels >>
rlabel locali s 674 669 674 669 4 Z
port 1 nsew
rlabel locali s 96 270 96 270 4 A
port 2 nsew
rlabel locali s 229 394 229 394 4 B
port 3 nsew
rlabel locali s 362 518 362 518 4 C
port 4 nsew
rlabel locali s 423 0 423 0 4 gnd
port 5 nsew
rlabel locali s 423 1414 423 1414 4 vdd
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 846 1414
string GDS_END 348542
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_8x1024_8.gds
string GDS_START 347294
<< end >>
