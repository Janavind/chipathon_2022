magic
tech sky130B
magscale 1 2
timestamp 1666199351
<< nwell >>
rect -38 261 1510 582
<< pwell >>
rect 1 21 1471 203
rect 30 -17 64 21
<< locali >>
rect 1034 373 1455 417
rect 20 289 715 325
rect 20 207 277 289
rect 332 249 601 255
rect 331 215 601 249
rect 332 207 601 215
rect 649 207 715 289
rect 1226 255 1270 339
rect 1000 207 1270 255
rect 1386 299 1455 373
rect 355 165 1271 173
rect 1421 165 1455 299
rect 355 139 1455 165
rect 355 135 666 139
rect 775 125 1455 139
rect 775 123 1009 125
rect 775 51 839 123
rect 975 51 1009 123
rect 1143 123 1455 125
rect 1143 51 1177 123
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 19 417 69 493
rect 103 451 169 527
rect 203 421 237 493
rect 271 455 337 527
rect 371 421 405 493
rect 439 455 505 527
rect 539 421 573 493
rect 607 455 673 527
rect 707 451 1454 493
rect 707 421 741 451
rect 203 417 741 421
rect 19 359 741 417
rect 775 357 982 417
rect 926 339 982 357
rect 749 289 766 323
rect 800 289 892 323
rect 926 289 1192 339
rect 749 255 892 289
rect 749 207 951 255
rect 1318 265 1352 289
rect 1318 199 1387 265
rect 113 139 321 173
rect 19 17 79 117
rect 113 106 155 139
rect 190 17 237 105
rect 271 101 321 139
rect 271 51 673 101
rect 707 17 741 105
rect 873 17 939 89
rect 1043 17 1109 89
rect 1211 17 1277 89
rect 1383 17 1454 89
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 766 289 800 323
rect 1318 289 1352 323
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
<< metal1 >>
rect 0 561 1472 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 0 496 1472 527
rect 754 323 812 329
rect 754 289 766 323
rect 800 320 812 323
rect 1306 323 1364 329
rect 1306 320 1318 323
rect 800 292 1318 320
rect 800 289 812 292
rect 754 283 812 289
rect 1306 289 1318 292
rect 1352 289 1364 323
rect 1306 283 1364 289
rect 0 17 1472 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
rect 0 -48 1472 -17
<< labels >>
rlabel locali s 332 207 601 215 6 A1
port 1 nsew signal input
rlabel locali s 331 215 601 249 6 A1
port 1 nsew signal input
rlabel locali s 332 249 601 255 6 A1
port 1 nsew signal input
rlabel locali s 649 207 715 289 6 A2
port 2 nsew signal input
rlabel locali s 20 207 277 289 6 A2
port 2 nsew signal input
rlabel locali s 20 289 715 325 6 A2
port 2 nsew signal input
rlabel metal1 s 1306 283 1364 292 6 B1
port 3 nsew signal input
rlabel metal1 s 754 283 812 292 6 B1
port 3 nsew signal input
rlabel metal1 s 754 292 1364 320 6 B1
port 3 nsew signal input
rlabel metal1 s 1306 320 1364 329 6 B1
port 3 nsew signal input
rlabel metal1 s 754 320 812 329 6 B1
port 3 nsew signal input
rlabel locali s 1000 207 1270 255 6 C1
port 4 nsew signal input
rlabel locali s 1226 255 1270 339 6 C1
port 4 nsew signal input
rlabel metal1 s 0 -48 1472 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 21 1471 203 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 1510 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 1472 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1143 51 1177 123 6 Y
port 9 nsew signal output
rlabel locali s 1143 123 1455 125 6 Y
port 9 nsew signal output
rlabel locali s 975 51 1009 123 6 Y
port 9 nsew signal output
rlabel locali s 775 51 839 123 6 Y
port 9 nsew signal output
rlabel locali s 775 123 1009 125 6 Y
port 9 nsew signal output
rlabel locali s 775 125 1455 139 6 Y
port 9 nsew signal output
rlabel locali s 355 135 666 139 6 Y
port 9 nsew signal output
rlabel locali s 355 139 1455 165 6 Y
port 9 nsew signal output
rlabel locali s 1421 165 1455 299 6 Y
port 9 nsew signal output
rlabel locali s 355 165 1271 173 6 Y
port 9 nsew signal output
rlabel locali s 1386 299 1455 373 6 Y
port 9 nsew signal output
rlabel locali s 1034 373 1455 417 6 Y
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1472 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3604130
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3593550
<< end >>
