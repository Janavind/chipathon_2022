magic
tech sky130B
magscale 1 2
timestamp 1666199351
use sky130_fd_pr__dfl1sd__example_55959141808336  sky130_fd_pr__dfl1sd__example_55959141808336_0
timestamp 1666199351
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808337  sky130_fd_pr__hvdfl1sd2__example_55959141808337_0
timestamp 1666199351
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808337  sky130_fd_pr__hvdfl1sd2__example_55959141808337_1
timestamp 1666199351
transform 1 0 256 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808338  sky130_fd_pr__hvdfl1sd__example_55959141808338_0
timestamp 1666199351
transform 1 0 412 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 32244072
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 32241984
<< end >>
