magic
tech sky130A
magscale 1 2
timestamp 1666464484
<< nwell >>
rect 0 236 1215 668
<< pwell >>
rect 827 150 1193 176
rect 40 14 1193 150
rect 827 -76 1193 14
<< mvnmos >>
rect 119 40 219 124
rect 275 40 375 124
rect 431 40 531 124
rect 619 40 719 124
rect 906 -50 1006 150
<< mvpmos >>
rect 119 302 219 602
rect 275 302 375 602
rect 431 302 531 602
rect 619 302 719 602
rect 888 402 988 602
<< mvndiff >>
rect 853 132 906 150
rect 66 86 119 124
rect 66 52 74 86
rect 108 52 119 86
rect 66 40 119 52
rect 219 86 275 124
rect 219 52 230 86
rect 264 52 275 86
rect 219 40 275 52
rect 375 86 431 124
rect 375 52 386 86
rect 420 52 431 86
rect 375 40 431 52
rect 531 86 619 124
rect 531 52 558 86
rect 592 52 619 86
rect 531 40 619 52
rect 719 86 772 124
rect 719 52 730 86
rect 764 52 772 86
rect 719 40 772 52
rect 853 98 861 132
rect 895 98 906 132
rect 853 64 906 98
rect 853 30 861 64
rect 895 30 906 64
rect 853 -4 906 30
rect 853 -38 861 -4
rect 895 -38 906 -4
rect 853 -50 906 -38
rect 1006 132 1059 150
rect 1006 98 1017 132
rect 1051 98 1059 132
rect 1006 64 1059 98
rect 1006 30 1017 64
rect 1051 30 1059 64
rect 1006 -4 1059 30
rect 1006 -38 1017 -4
rect 1051 -38 1059 -4
rect 1006 -50 1059 -38
<< mvpdiff >>
rect 66 590 119 602
rect 66 556 74 590
rect 108 556 119 590
rect 66 522 119 556
rect 66 488 74 522
rect 108 488 119 522
rect 66 454 119 488
rect 66 420 74 454
rect 108 420 119 454
rect 66 386 119 420
rect 66 352 74 386
rect 108 352 119 386
rect 66 302 119 352
rect 219 590 275 602
rect 219 556 230 590
rect 264 556 275 590
rect 219 522 275 556
rect 219 488 230 522
rect 264 488 275 522
rect 219 454 275 488
rect 219 420 230 454
rect 264 420 275 454
rect 219 386 275 420
rect 219 352 230 386
rect 264 352 275 386
rect 219 302 275 352
rect 375 590 431 602
rect 375 556 386 590
rect 420 556 431 590
rect 375 522 431 556
rect 375 488 386 522
rect 420 488 431 522
rect 375 454 431 488
rect 375 420 386 454
rect 420 420 431 454
rect 375 386 431 420
rect 375 352 386 386
rect 420 352 431 386
rect 375 302 431 352
rect 531 590 619 602
rect 531 556 542 590
rect 576 556 619 590
rect 531 522 619 556
rect 531 488 542 522
rect 576 488 619 522
rect 531 454 619 488
rect 531 420 542 454
rect 576 420 619 454
rect 531 386 619 420
rect 531 352 542 386
rect 576 352 619 386
rect 531 302 619 352
rect 719 590 775 602
rect 719 556 730 590
rect 764 556 775 590
rect 719 522 775 556
rect 719 488 730 522
rect 764 488 775 522
rect 719 454 775 488
rect 719 420 730 454
rect 764 420 775 454
rect 719 386 775 420
rect 835 590 888 602
rect 835 556 843 590
rect 877 556 888 590
rect 835 522 888 556
rect 835 488 843 522
rect 877 488 888 522
rect 835 454 888 488
rect 835 420 843 454
rect 877 420 888 454
rect 835 402 888 420
rect 988 590 1041 602
rect 988 556 999 590
rect 1033 556 1041 590
rect 988 522 1041 556
rect 988 488 999 522
rect 1033 488 1041 522
rect 988 454 1041 488
rect 988 420 999 454
rect 1033 420 1041 454
rect 988 402 1041 420
rect 719 352 730 386
rect 764 352 775 386
rect 719 302 775 352
<< mvndiffc >>
rect 74 52 108 86
rect 230 52 264 86
rect 386 52 420 86
rect 558 52 592 86
rect 730 52 764 86
rect 861 98 895 132
rect 861 30 895 64
rect 861 -38 895 -4
rect 1017 98 1051 132
rect 1017 30 1051 64
rect 1017 -38 1051 -4
<< mvpdiffc >>
rect 74 556 108 590
rect 74 488 108 522
rect 74 420 108 454
rect 74 352 108 386
rect 230 556 264 590
rect 230 488 264 522
rect 230 420 264 454
rect 230 352 264 386
rect 386 556 420 590
rect 386 488 420 522
rect 386 420 420 454
rect 386 352 420 386
rect 542 556 576 590
rect 542 488 576 522
rect 542 420 576 454
rect 542 352 576 386
rect 730 556 764 590
rect 730 488 764 522
rect 730 420 764 454
rect 843 556 877 590
rect 843 488 877 522
rect 843 420 877 454
rect 999 556 1033 590
rect 999 488 1033 522
rect 999 420 1033 454
rect 730 352 764 386
<< mvpsubdiff >>
rect 1133 126 1167 150
rect 1133 8 1167 92
rect 1133 -50 1167 -26
<< mvnsubdiff >>
rect 1115 578 1149 602
rect 1115 505 1149 544
rect 1115 432 1149 471
rect 1115 360 1149 398
rect 1115 302 1149 326
<< mvpsubdiffcont >>
rect 1133 92 1167 126
rect 1133 -26 1167 8
<< mvnsubdiffcont >>
rect 1115 544 1149 578
rect 1115 471 1149 505
rect 1115 398 1149 432
rect 1115 326 1149 360
<< poly >>
rect 119 602 219 628
rect 275 602 375 628
rect 431 602 531 628
rect 619 602 719 628
rect 888 602 988 628
rect 888 356 988 402
rect 888 340 1093 356
rect 888 306 975 340
rect 1009 306 1043 340
rect 1077 306 1093 340
rect 119 276 219 302
rect 275 276 375 302
rect 431 276 531 302
rect 119 252 531 276
rect 619 270 719 302
rect 888 290 1093 306
rect 119 218 135 252
rect 169 218 219 252
rect 253 218 302 252
rect 336 218 531 252
rect 119 150 531 218
rect 573 254 719 270
rect 573 220 589 254
rect 623 220 657 254
rect 691 220 719 254
rect 573 204 719 220
rect 119 124 219 150
rect 275 124 375 150
rect 431 124 531 150
rect 619 124 719 204
rect 873 232 1007 248
rect 873 198 889 232
rect 923 198 957 232
rect 991 198 1007 232
rect 873 182 1007 198
rect 906 150 1006 182
rect 119 14 219 40
rect 275 14 375 40
rect 431 14 531 40
rect 619 14 719 40
rect 906 -76 1006 -50
<< polycont >>
rect 975 306 1009 340
rect 1043 306 1077 340
rect 135 218 169 252
rect 219 218 253 252
rect 302 218 336 252
rect 589 220 623 254
rect 657 220 691 254
rect 889 198 923 232
rect 957 198 991 232
<< locali >>
rect 230 640 576 674
rect 74 590 108 606
rect 74 522 108 556
rect 74 454 108 488
rect 74 386 108 420
rect 74 336 108 352
rect 230 590 264 640
rect 230 522 264 556
rect 230 454 264 488
rect 230 386 264 420
rect 230 336 264 352
rect 386 590 420 606
rect 386 522 420 556
rect 386 454 420 488
rect 386 386 420 420
rect 386 270 420 352
rect 542 590 576 640
rect 542 522 576 556
rect 542 454 576 488
rect 542 386 576 420
rect 542 336 576 352
rect 725 590 773 606
rect 725 556 730 590
rect 764 556 773 590
rect 725 522 773 556
rect 725 488 730 522
rect 764 488 773 522
rect 725 454 773 488
rect 725 420 730 454
rect 764 420 773 454
rect 725 386 773 420
rect 725 352 730 386
rect 764 352 773 386
rect 725 271 773 352
rect 807 590 877 606
rect 807 556 843 590
rect 807 522 877 556
rect 807 488 843 522
rect 807 454 877 488
rect 999 590 1149 606
rect 1033 578 1149 590
rect 1033 556 1115 578
rect 999 544 1115 556
rect 999 522 1149 544
rect 1033 505 1149 522
rect 1033 488 1115 505
rect 999 483 1115 488
rect 807 420 843 454
rect 807 404 877 420
rect 911 471 1115 483
rect 911 454 1149 471
rect 911 420 999 454
rect 1033 432 1149 454
rect 1033 420 1115 432
rect 386 254 691 270
rect 119 218 135 252
rect 169 218 219 252
rect 253 218 302 252
rect 336 218 352 252
rect 386 220 589 254
rect 623 220 657 254
rect 386 204 691 220
rect 74 86 108 130
rect 74 36 108 52
rect 230 86 264 102
rect 230 2 264 52
rect 386 86 420 204
rect 725 170 759 271
rect 807 237 855 404
rect 911 398 1115 420
rect 911 390 1149 398
rect 911 388 950 390
rect 907 384 950 388
rect 905 380 950 384
rect 902 378 949 380
rect 902 374 946 378
rect 902 370 944 374
rect 902 248 941 370
rect 1115 360 1149 390
rect 975 340 1077 356
rect 1009 306 1043 340
rect 975 290 1077 306
rect 1115 302 1149 326
rect 659 136 759 170
rect 793 182 855 237
rect 889 232 991 248
rect 923 198 957 232
rect 889 182 991 198
rect 386 36 420 52
rect 558 86 592 102
rect 558 2 592 52
rect 230 -32 592 2
rect 659 2 696 136
rect 793 102 827 182
rect 1025 148 1077 290
rect 730 86 827 102
rect 764 52 827 86
rect 730 36 827 52
rect 861 132 895 148
rect 861 64 895 98
rect 861 2 895 30
rect 659 -4 895 2
rect 659 -32 861 -4
rect 861 -54 895 -38
rect 1017 132 1077 148
rect 1051 98 1077 132
rect 1017 64 1077 98
rect 1051 30 1077 64
rect 1017 -4 1077 30
rect 1051 -38 1077 -4
rect 1017 -54 1077 -38
rect 1133 126 1167 150
rect 1133 8 1167 92
rect 1133 -50 1167 -26
use sky130_fd_pr__nfet_01v8__example_55959141808109  sky130_fd_pr__nfet_01v8__example_55959141808109_0
timestamp 1666464484
transform -1 0 1006 0 1 -50
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808110  sky130_fd_pr__nfet_01v8__example_55959141808110_0
timestamp 1666464484
transform 1 0 619 0 1 40
box -17 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808111  sky130_fd_pr__nfet_01v8__example_55959141808111_0
timestamp 1666464484
transform 1 0 431 0 1 40
box -1 0 117 1
use sky130_fd_pr__nfet_01v8__example_55959141808112  sky130_fd_pr__nfet_01v8__example_55959141808112_0
timestamp 1666464484
transform 1 0 275 0 1 40
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808113  sky130_fd_pr__nfet_01v8__example_55959141808113_0
timestamp 1666464484
transform 1 0 119 0 1 40
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808103  sky130_fd_pr__pfet_01v8__example_55959141808103_0
timestamp 1666464484
transform 1 0 619 0 -1 602
box -33 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808105  sky130_fd_pr__pfet_01v8__example_55959141808105_0
timestamp 1666464484
transform 1 0 275 0 -1 602
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_55959141808107  sky130_fd_pr__pfet_01v8__example_55959141808107_0
timestamp 1666464484
transform -1 0 988 0 -1 602
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808108  sky130_fd_pr__pfet_01v8__example_55959141808108_0
timestamp 1666464484
transform 1 0 119 0 -1 602
box -1 0 101 1
<< labels >>
flabel locali s 1017 27 1051 93 3 FreeSans 200 180 0 0 VGND
port 1 nsew
flabel locali s 74 405 108 471 3 FreeSans 200 0 0 0 VCC_IO
port 2 nsew
flabel locali s 74 62 108 128 3 FreeSans 200 0 0 0 VGND
port 1 nsew
flabel locali s 119 218 135 252 3 FreeSans 200 0 0 0 IN
port 3 nsew
flabel locali s 1063 405 1097 471 0 FreeSans 200 0 0 0 VCC_IO
port 2 nsew
flabel locali s 543 218 559 252 3 FreeSans 200 0 0 0 OUT
port 4 nsew
flabel locali s 1133 66 1167 150 0 FreeSans 200 0 0 0 VGND
port 1 nsew
flabel locali s 433 -12 433 -12 7 FreeSans 200 0 0 0 INT_N
port 5 nsew
flabel locali s 434 658 434 658 7 FreeSans 200 0 0 0 INT_P
port 6 nsew
<< properties >>
string GDS_END 33982688
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 33977068
<< end >>
