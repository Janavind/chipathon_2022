magic
tech sky130B
timestamp 1666464484
<< properties >>
string GDS_END 1499836
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 1497656
<< end >>
