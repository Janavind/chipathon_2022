magic
tech sky130A
magscale 1 2
timestamp 1666199351
<< metal1 >>
rect 12486 -407 12538 -351
<< metal2 >>
rect 7956 15977 8019 15991
rect 7956 15927 7969 15977
tri 7969 15927 8019 15977 nw
rect 675 -407 721 -361
rect 1084 -407 1130 -328
rect 1226 -407 1278 -355
rect 2551 -407 2603 -363
rect 3262 -407 3314 -306
rect 4471 -407 4523 -340
rect 5320 -407 5372 -379
rect 5698 -407 5750 -355
rect 6150 -407 6202 -351
rect 6363 -407 6415 -363
rect 7092 -407 7144 -351
rect 7678 -407 7730 -318
rect 9049 -407 9101 -355
rect 9971 -407 10023 -355
rect 13367 -407 13419 -355
rect 13655 -407 13785 -363
rect 15256 -407 15384 -363
rect 15522 -407 15574 -363
rect 15741 -407 15781 -363
rect 15943 -407 15983 -215
<< metal3 >>
rect 80 -407 204 -244
rect 9173 -407 9239 -355
rect 12564 -407 12778 -260
rect 15716 -407 15782 -254
rect 15848 -407 15914 -244
<< metal4 >>
rect 0 34750 254 39593
rect 15746 34750 16000 39593
rect 0 13600 254 18593
rect 15746 13600 16000 18593
rect 0 12410 254 13300
rect 15746 12410 16000 13300
rect 0 11240 254 12130
rect 15746 11240 16000 12130
rect 0 10874 254 10940
rect 15746 10874 16000 10940
rect 0 10218 254 10814
rect 15746 10218 16000 10814
rect 0 9922 254 10158
rect 15746 9922 16000 10158
rect 0 9266 254 9862
rect 15746 9266 16000 9862
rect 0 9140 254 9206
rect 15746 9140 16000 9206
rect 0 7910 254 8840
rect 15746 7910 16000 8840
rect 0 6940 254 7630
rect 15746 6940 16000 7630
rect 0 5970 254 6660
rect 15746 5970 16000 6660
rect 0 4760 254 5690
rect 15746 4760 16000 5690
rect 0 3550 254 4480
rect 15746 3550 16000 4480
rect 0 2580 254 3270
rect 15746 2580 16000 3270
rect 0 1370 254 2300
rect 15746 1370 16000 2300
rect 0 0 254 1090
rect 15746 0 16000 1090
<< metal5 >>
rect 0 34750 254 39593
rect 15746 34750 16000 39593
rect 6423 24687 10731 28996
rect 0 13600 254 18590
rect 15746 13600 16000 18590
rect 0 12430 254 13280
rect 15746 12430 16000 13280
rect 0 11260 254 12110
rect 15746 11260 16000 12110
rect 0 9140 254 10940
rect 15746 9140 16000 10940
rect 0 7930 254 8820
rect 15746 7930 16000 8820
rect 0 6960 254 7610
rect 15746 6960 16000 7610
rect 0 5990 254 6640
rect 15746 5990 16000 6640
rect 0 4780 254 5670
rect 15746 4780 16000 5670
rect 0 3570 254 4460
rect 15746 3570 16000 4460
rect 0 2600 254 3250
rect 15746 2600 16000 3250
rect 0 1390 254 2280
rect 15746 1390 16000 2280
rect 0 20 254 1070
rect 15746 20 16000 1070
use sky130_fd_io__overlay_gpiov2  sky130_fd_io__overlay_gpiov2_0
timestamp 1666199351
transform 1 0 0 0 1 -407
box 0 407 16000 40000
use sky130_fd_io__top_gpiov2  sky130_fd_io__top_gpiov2_0
timestamp 1666199351
transform 1 0 0 0 1 -407
box -143 -136 16134 40000
<< labels >>
flabel metal4 s 0 10218 254 10814 3 FreeSans 650 0 0 0 AMUXBUS_A
port 28 nsew
flabel metal4 s 15746 10218 16000 10814 3 FreeSans 650 180 0 0 AMUXBUS_A
port 28 nsew
flabel metal4 s 0 9266 254 9862 3 FreeSans 650 0 0 0 AMUXBUS_B
port 29 nsew
flabel metal4 s 15746 9266 16000 9862 3 FreeSans 650 180 0 0 AMUXBUS_B
port 29 nsew
flabel metal1 s 12486 -407 12538 -351 0 FreeSans 500 270 0 0 ANALOG_EN
port 22 nsew
flabel metal3 s 9173 -407 9239 -355 0 FreeSans 500 270 0 0 ANALOG_POL
port 26 nsew
flabel metal2 s 6150 -407 6202 -351 0 FreeSans 500 270 0 0 ANALOG_SEL
port 23 nsew
flabel metal2 s 5698 -407 5750 -355 0 FreeSans 500 270 0 0 DM[2]
port 6 nsew
flabel metal2 s 13367 -407 13419 -355 0 FreeSans 500 270 0 0 DM[1]
port 7 nsew
flabel metal2 s 9971 -407 10023 -355 0 FreeSans 500 270 0 0 DM[0]
port 8 nsew
flabel metal2 s 7092 -407 7144 -351 0 FreeSans 500 270 0 0 ENABLE_H
port 13 nsew
flabel metal2 s 7678 -407 7730 -318 0 FreeSans 500 270 0 0 ENABLE_INP_H
port 15 nsew
flabel metal2 s 2551 -407 2603 -363 0 FreeSans 500 270 0 0 ENABLE_VDDA_H
port 14 nsew
flabel metal3 s 15716 -407 15782 -254 0 FreeSans 500 270 0 0 ENABLE_VDDIO
port 24 nsew
flabel metal2 s 3262 -407 3314 -306 0 FreeSans 500 270 0 0 ENABLE_VSWITCH_H
port 25 nsew
flabel metal2 s 6363 -407 6415 -363 0 FreeSans 500 270 0 0 HLD_H_N
port 9 nsew
flabel metal2 s 5320 -407 5372 -379 0 FreeSans 500 270 0 0 HLD_OVR
port 21 nsew
flabel metal2 s 1084 -407 1130 -328 0 FreeSans 500 270 0 0 IB_MODE_SEL
port 12 nsew
flabel metal3 s 15848 -407 15914 -244 0 FreeSans 500 270 0 0 IN
port 10 nsew
flabel metal3 s 80 -407 204 -244 0 FreeSans 800 0 0 0 IN_H
port 1 nsew
flabel metal2 s 9049 -407 9101 -355 0 FreeSans 500 270 0 0 INP_DIS
port 11 nsew
flabel metal2 s 675 -407 721 -361 0 FreeSans 500 270 0 0 OE_N
port 16 nsew
flabel metal2 s 4471 -407 4523 -340 0 FreeSans 500 0 0 0 OUT
port 27 nsew
flabel metal5 s 6423 24687 10731 28996 0 FreeSans 2000 0 0 0 PAD
port 5 nsew
flabel metal2 s 15256 -407 15384 -363 0 FreeSans 500 270 0 0 PAD_A_ESD_0_H
port 3 nsew
flabel metal2 s 13655 -407 13785 -363 0 FreeSans 500 270 0 0 PAD_A_ESD_1_H
port 4 nsew
flabel metal3 s 12564 -407 12778 -260 0 FreeSans 500 270 0 0 PAD_A_NOESD_H
port 2 nsew
flabel metal2 s 15522 -407 15574 -363 0 FreeSans 500 270 0 0 SLOW
port 19 nsew
flabel metal2 s 15741 -407 15781 -363 0 FreeSans 500 270 0 0 TIE_HI_ESD
port 17 nsew
flabel metal2 s 15943 -407 15983 -215 0 FreeSans 500 270 0 0 TIE_LO_ESD
port 18 nsew
flabel metal5 s 0 1390 254 2280 3 FreeSans 650 0 0 0 VCCD
port 36 nsew
flabel metal4 s 0 1370 254 2300 3 FreeSans 650 0 0 0 VCCD
port 36 nsew
flabel metal5 s 15746 1390 16000 2280 3 FreeSans 650 180 0 0 VCCD
port 36 nsew
flabel metal4 s 15746 1370 16000 2300 3 FreeSans 650 180 0 0 VCCD
port 36 nsew
flabel metal5 s 0 20 254 1070 3 FreeSans 650 0 0 0 VCCHIB
port 34 nsew
flabel metal4 s 0 0 254 1090 3 FreeSans 650 0 0 0 VCCHIB
port 34 nsew
flabel metal5 s 15746 20 16000 1070 3 FreeSans 650 180 0 0 VCCHIB
port 34 nsew
flabel metal4 s 15746 0 16000 1090 3 FreeSans 650 180 0 0 VCCHIB
port 34 nsew
flabel metal5 s 0 2600 193 3250 3 FreeSans 650 0 0 0 VDDA
port 31 nsew
flabel metal4 s 0 2580 193 3270 3 FreeSans 650 0 0 0 VDDA
port 31 nsew
flabel metal5 s 15807 2600 16000 3250 3 FreeSans 650 180 0 0 VDDA
port 31 nsew
flabel metal4 s 15807 2580 16000 3270 3 FreeSans 650 180 0 0 VDDA
port 31 nsew
flabel metal5 s 0 13600 254 18590 3 FreeSans 650 0 0 0 VDDIO
port 35 nsew
flabel metal5 s 0 3570 254 4460 3 FreeSans 650 0 0 0 VDDIO
port 35 nsew
flabel metal4 s 0 3550 254 4480 3 FreeSans 650 0 0 0 VDDIO
port 35 nsew
flabel metal4 s 0 13600 254 18593 3 FreeSans 650 0 0 0 VDDIO
port 35 nsew
flabel metal5 s 15746 13600 16000 18590 3 FreeSans 650 180 0 0 VDDIO
port 35 nsew
flabel metal5 s 15746 3570 16000 4460 3 FreeSans 650 180 0 0 VDDIO
port 35 nsew
flabel metal4 s 15746 3550 16000 4480 3 FreeSans 650 180 0 0 VDDIO
port 35 nsew
flabel metal4 s 15746 13600 16000 18593 3 FreeSans 650 180 0 0 VDDIO
port 35 nsew
flabel metal5 s 0 12430 254 13280 3 FreeSans 650 0 0 0 VDDIO_Q
port 33 nsew
flabel metal4 s 0 12410 254 13300 3 FreeSans 650 0 0 0 VDDIO_Q
port 33 nsew
flabel metal5 s 15746 12430 16000 13280 3 FreeSans 650 180 0 0 VDDIO_Q
port 33 nsew
flabel metal4 s 15746 12410 16000 13300 3 FreeSans 650 180 0 0 VDDIO_Q
port 33 nsew
flabel metal5 s 0 9140 254 10940 3 FreeSans 650 0 0 0 VSSA
port 30 nsew
flabel metal5 s 0 6961 254 7610 3 FreeSans 650 0 0 0 VSSA
port 30 nsew
flabel metal4 s 0 9140 254 9206 3 FreeSans 650 0 0 0 VSSA
port 30 nsew
flabel metal4 s 0 9922 254 10158 3 FreeSans 650 0 0 0 VSSA
port 30 nsew
flabel metal4 s 0 10874 254 10940 3 FreeSans 650 0 0 0 VSSA
port 30 nsew
flabel metal4 s 0 6940 254 7630 3 FreeSans 650 0 0 0 VSSA
port 30 nsew
flabel metal5 s 15746 9140 16000 10940 3 FreeSans 650 180 0 0 VSSA
port 30 nsew
flabel metal5 s 15746 6961 16000 7610 3 FreeSans 650 180 0 0 VSSA
port 30 nsew
flabel metal4 s 15746 9922 16000 10158 3 FreeSans 650 180 0 0 VSSA
port 30 nsew
flabel metal4 s 15746 10874 16000 10940 3 FreeSans 650 180 0 0 VSSA
port 30 nsew
flabel metal4 s 15746 9140 16000 9206 3 FreeSans 650 180 0 0 VSSA
port 30 nsew
flabel metal4 s 15746 6940 16000 7630 3 FreeSans 650 180 0 0 VSSA
port 30 nsew
flabel metal5 s 0 7930 254 8820 3 FreeSans 650 0 0 0 VSSD
port 38 nsew
flabel metal4 s 0 7910 254 8840 3 FreeSans 650 0 0 0 VSSD
port 38 nsew
flabel metal5 s 15746 7930 16000 8820 3 FreeSans 650 180 0 0 VSSD
port 38 nsew
flabel metal4 s 15746 7910 16000 8840 3 FreeSans 650 180 0 0 VSSD
port 38 nsew
flabel metal4 s 0 34750 254 39593 3 FreeSans 650 0 0 0 VSSIO
port 37 nsew
flabel metal5 s 0 4780 254 5670 3 FreeSans 650 0 0 0 VSSIO
port 37 nsew
flabel metal4 s 127 37171 127 37171 3 FreeSans 650 0 0 0 VSSIO
port 37 nsew
flabel metal4 s 0 4760 254 5690 3 FreeSans 650 0 0 0 VSSIO
port 37 nsew
flabel metal4 s 15746 34750 16000 39593 3 FreeSans 650 180 0 0 VSSIO
port 37 nsew
flabel metal5 s 15746 4780 16000 5670 3 FreeSans 650 180 0 0 VSSIO
port 37 nsew
flabel metal4 s 15746 4760 16000 5690 3 FreeSans 650 180 0 0 VSSIO
port 37 nsew
flabel metal4 s 15873 37171 15873 37171 3 FreeSans 650 180 0 0 VSSIO
port 37 nsew
flabel metal5 s 0 11260 254 12110 3 FreeSans 650 0 0 0 VSSIO_Q
port 39 nsew
flabel metal4 s 0 11240 254 12130 3 FreeSans 650 0 0 0 VSSIO_Q
port 39 nsew
flabel metal5 s 15746 11260 16000 12110 3 FreeSans 650 180 0 0 VSSIO_Q
port 39 nsew
flabel metal4 s 15746 11240 16000 12130 3 FreeSans 650 180 0 0 VSSIO_Q
port 39 nsew
flabel metal5 s 0 5990 254 6640 3 FreeSans 650 0 0 0 VSWITCH
port 32 nsew
flabel metal4 s 0 5970 254 6660 3 FreeSans 650 0 0 0 VSWITCH
port 32 nsew
flabel metal5 s 15746 5990 16000 6640 3 FreeSans 650 180 0 0 VSWITCH
port 32 nsew
flabel metal4 s 15746 5970 16000 6660 3 FreeSans 650 180 0 0 VSWITCH
port 32 nsew
flabel metal2 s 1226 -407 1278 -355 0 FreeSans 500 270 0 0 VTRIP_SEL
port 20 nsew
<< properties >>
string FIXED_BBOX 0 0 16000 39593
string GDS_END 2545096
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io.gds
string GDS_START 2527264
<< end >>
