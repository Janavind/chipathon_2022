magic
tech sky130A
timestamp 1666464484
<< obsm1 >>
rect 62 62 45468 44584
<< obsm2 >>
rect 62 62 45468 44584
<< metal3 >>
rect 136 44336 45394 44510
rect 476 43996 45054 44170
rect 45424 39848 45530 39886
rect 45424 39576 45530 39614
rect 0 18496 106 18534
rect 0 17952 106 17990
rect 0 17136 106 17174
rect 0 16592 106 16630
rect 0 15776 106 15814
rect 0 15096 106 15134
rect 0 14280 106 14318
rect 45424 9860 45530 9898
rect 45424 8976 45530 9014
rect 45424 8432 45530 8470
rect 45424 7548 45530 7586
rect 45424 7004 45530 7042
rect 45424 6188 45530 6226
rect 45424 5508 45530 5546
rect 0 5100 106 5138
rect 0 4284 106 4322
rect 0 4148 106 4186
rect 476 476 45054 650
rect 136 136 45394 310
<< obsm3 >>
rect 62 44570 45468 44584
rect 62 44276 76 44570
rect 45454 44276 45468 44570
rect 62 44230 45468 44276
rect 62 43936 416 44230
rect 45114 43936 45468 44230
rect 62 39946 45468 43936
rect 62 39788 45364 39946
rect 62 39674 45468 39788
rect 62 39516 45364 39674
rect 62 18594 45468 39516
rect 166 18436 45468 18594
rect 62 18050 45468 18436
rect 166 17892 45468 18050
rect 62 17234 45468 17892
rect 166 17076 45468 17234
rect 62 16690 45468 17076
rect 166 16532 45468 16690
rect 62 15874 45468 16532
rect 166 15716 45468 15874
rect 62 15194 45468 15716
rect 166 15036 45468 15194
rect 62 14378 45468 15036
rect 166 14220 45468 14378
rect 62 9958 45468 14220
rect 62 9800 45364 9958
rect 62 9074 45468 9800
rect 62 8916 45364 9074
rect 62 8530 45468 8916
rect 62 8372 45364 8530
rect 62 7646 45468 8372
rect 62 7488 45364 7646
rect 62 7102 45468 7488
rect 62 6944 45364 7102
rect 62 6286 45468 6944
rect 62 6128 45364 6286
rect 62 5606 45468 6128
rect 62 5448 45364 5606
rect 62 5198 45468 5448
rect 166 5040 45468 5198
rect 62 4382 45468 5040
rect 166 4088 45468 4382
rect 62 710 45468 4088
rect 62 416 416 710
rect 45114 416 45468 710
rect 62 370 45468 416
rect 62 76 76 370
rect 45454 76 45468 370
rect 62 62 45468 76
<< metal4 >>
rect 136 136 310 44510
rect 12784 44540 12822 44646
rect 15300 44540 15338 44646
rect 17816 44540 17854 44646
rect 20332 44540 20370 44646
rect 22780 44540 22818 44646
rect 25228 44540 25266 44646
rect 27812 44540 27850 44646
rect 30328 44540 30366 44646
rect 37264 44540 37302 44646
rect 37808 44540 37846 44646
rect 38352 44540 38390 44646
rect 476 476 650 44170
rect 44880 476 45054 44170
rect 6460 0 6498 106
rect 7140 0 7178 106
rect 7684 0 7722 106
rect 8228 0 8266 106
rect 8840 0 8878 106
rect 9452 0 9490 106
rect 9996 0 10034 106
rect 10540 0 10578 106
rect 11152 0 11190 106
rect 11696 0 11734 106
rect 12376 0 12414 106
rect 12648 0 12686 106
rect 12852 0 12890 106
rect 15232 0 15270 106
rect 17748 0 17786 106
rect 20264 0 20302 106
rect 22780 0 22818 106
rect 25228 0 25266 106
rect 27744 0 27782 106
rect 30260 0 30298 106
rect 45220 136 45394 44510
<< obsm4 >>
rect 62 44570 12724 44584
rect 62 76 76 44570
rect 370 44480 12724 44570
rect 12882 44480 15240 44584
rect 15398 44480 17756 44584
rect 17914 44480 20272 44584
rect 20430 44480 22720 44584
rect 22878 44480 25168 44584
rect 25326 44480 27752 44584
rect 27910 44480 30268 44584
rect 30426 44480 37204 44584
rect 37362 44480 37748 44584
rect 37906 44480 38292 44584
rect 38450 44570 45468 44584
rect 38450 44480 45160 44570
rect 370 44230 45160 44480
rect 370 416 416 44230
rect 710 416 44820 44230
rect 45114 416 45160 44230
rect 370 166 45160 416
rect 370 76 6400 166
rect 62 62 6400 76
rect 6558 62 7080 166
rect 7238 62 7624 166
rect 7782 62 8168 166
rect 8326 62 8780 166
rect 8938 62 9392 166
rect 9550 62 9936 166
rect 10094 62 10480 166
rect 10638 62 11092 166
rect 11250 62 11636 166
rect 11794 62 12316 166
rect 12474 62 12588 166
rect 12746 62 12792 166
rect 12950 62 15172 166
rect 15330 62 17688 166
rect 17846 62 20204 166
rect 20362 62 22720 166
rect 22878 62 25168 166
rect 25326 62 27684 166
rect 27842 62 30200 166
rect 30358 76 45160 166
rect 45454 76 45468 44570
rect 30358 62 45468 76
<< labels >>
rlabel metal4 s 8840 0 8878 106 6 din0[0]
port 8 nsew default input
rlabel metal4 s 9452 0 9490 106 6 din0[1]
port 7 nsew default input
rlabel metal4 s 9996 0 10034 106 6 din0[2]
port 6 nsew default input
rlabel metal4 s 10540 0 10578 106 6 din0[3]
port 5 nsew default input
rlabel metal4 s 11152 0 11190 106 6 din0[4]
port 4 nsew default input
rlabel metal4 s 11696 0 11734 106 6 din0[5]
port 3 nsew default input
rlabel metal4 s 12376 0 12414 106 6 din0[6]
port 2 nsew default input
rlabel metal4 s 12852 0 12890 106 6 din0[7]
port 1 nsew default input
rlabel metal4 s 6460 0 6498 106 6 addr0[0]
port 18 nsew default input
rlabel metal4 s 7140 0 7178 106 6 addr0[1]
port 17 nsew default input
rlabel metal4 s 7684 0 7722 106 6 addr0[2]
port 16 nsew default input
rlabel metal3 s 0 14280 106 14318 6 addr0[3]
port 15 nsew default input
rlabel metal3 s 0 15096 106 15134 6 addr0[4]
port 14 nsew default input
rlabel metal3 s 0 15776 106 15814 6 addr0[5]
port 13 nsew default input
rlabel metal3 s 0 16592 106 16630 6 addr0[6]
port 12 nsew default input
rlabel metal3 s 0 17136 106 17174 6 addr0[7]
port 11 nsew default input
rlabel metal3 s 0 17952 106 17990 6 addr0[8]
port 10 nsew default input
rlabel metal3 s 0 18496 106 18534 6 addr0[9]
port 9 nsew default input
rlabel metal4 s 38352 44540 38390 44646 6 addr1[0]
port 28 nsew default input
rlabel metal4 s 37808 44540 37846 44646 6 addr1[1]
port 27 nsew default input
rlabel metal4 s 37264 44540 37302 44646 6 addr1[2]
port 26 nsew default input
rlabel metal3 s 45424 9860 45530 9898 6 addr1[3]
port 25 nsew default input
rlabel metal3 s 45424 8976 45530 9014 6 addr1[4]
port 24 nsew default input
rlabel metal3 s 45424 8432 45530 8470 6 addr1[5]
port 23 nsew default input
rlabel metal3 s 45424 7548 45530 7586 6 addr1[6]
port 22 nsew default input
rlabel metal3 s 45424 7004 45530 7042 6 addr1[7]
port 21 nsew default input
rlabel metal3 s 45424 6188 45530 6226 6 addr1[8]
port 20 nsew default input
rlabel metal3 s 45424 5508 45530 5546 6 addr1[9]
port 19 nsew default input
rlabel metal3 s 0 4284 106 4322 6 csb0
port 29 nsew default input
rlabel metal3 s 45424 39848 45530 39886 6 csb1
port 30 nsew default input
rlabel metal3 s 0 5100 106 5138 6 web0
port 31 nsew default input
rlabel metal3 s 0 4148 106 4186 6 clk0
port 32 nsew default input
rlabel metal3 s 45424 39576 45530 39614 6 clk1
port 33 nsew default input
rlabel metal4 s 8228 0 8266 106 6 wmask0[0]
port 34 nsew default input
rlabel metal4 s 12648 0 12686 106 6 dout0[0]
port 42 nsew default output
rlabel metal4 s 15232 0 15270 106 6 dout0[1]
port 41 nsew default output
rlabel metal4 s 17748 0 17786 106 6 dout0[2]
port 40 nsew default output
rlabel metal4 s 20264 0 20302 106 6 dout0[3]
port 39 nsew default output
rlabel metal4 s 22780 0 22818 106 6 dout0[4]
port 38 nsew default output
rlabel metal4 s 25228 0 25266 106 6 dout0[5]
port 37 nsew default output
rlabel metal4 s 27744 0 27782 106 6 dout0[6]
port 36 nsew default output
rlabel metal4 s 30260 0 30298 106 6 dout0[7]
port 35 nsew default output
rlabel metal4 s 12784 44540 12822 44646 6 dout1[0]
port 50 nsew default output
rlabel metal4 s 15300 44540 15338 44646 6 dout1[1]
port 49 nsew default output
rlabel metal4 s 17816 44540 17854 44646 6 dout1[2]
port 48 nsew default output
rlabel metal4 s 20332 44540 20370 44646 6 dout1[3]
port 47 nsew default output
rlabel metal4 s 22780 44540 22818 44646 6 dout1[4]
port 46 nsew default output
rlabel metal4 s 25228 44540 25266 44646 6 dout1[5]
port 45 nsew default output
rlabel metal4 s 27812 44540 27850 44646 6 dout1[6]
port 44 nsew default output
rlabel metal4 s 30328 44540 30366 44646 6 dout1[7]
port 43 nsew default output
rlabel metal4 s 476 476 650 44170 6 vccd1
port 51 nsew power bidirectional abutment
rlabel metal3 s 476 476 45054 650 6 vccd1
port 51 nsew power bidirectional abutment
rlabel metal3 s 476 43996 45054 44170 6 vccd1
port 51 nsew power bidirectional abutment
rlabel metal4 s 44880 476 45054 44170 6 vccd1
port 51 nsew power bidirectional abutment
rlabel metal3 s 136 44336 45394 44510 6 vssd1
port 52 nsew ground bidirectional abutment
rlabel metal3 s 136 136 45394 310 6 vssd1
port 52 nsew ground bidirectional abutment
rlabel metal4 s 45220 136 45394 44510 6 vssd1
port 52 nsew ground bidirectional abutment
rlabel metal4 s 136 136 310 44510 6 vssd1
port 52 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 45530 44646
string LEFclass BLOCK
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 9277678
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_8x1024_8.gds
string GDS_START 7724596
<< end >>
