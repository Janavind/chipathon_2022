magic
tech sky130A
magscale 1 2
timestamp 1666464484
<< nwell >>
rect -38 261 590 582
<< pwell >>
rect 362 163 551 203
rect 1 27 551 163
rect 30 -17 64 27
rect 362 21 551 27
<< locali >>
rect 18 425 349 483
rect 18 151 88 265
rect 122 199 264 323
rect 481 299 535 493
rect 298 199 379 265
rect 501 152 535 299
rect 481 83 535 152
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 18 357 336 391
rect 383 367 439 527
rect 18 299 82 357
rect 302 333 336 357
rect 302 299 447 333
rect 413 265 447 299
rect 413 199 467 265
rect 413 165 447 199
rect 125 131 447 165
rect 19 17 85 117
rect 125 61 159 131
rect 199 17 265 97
rect 299 61 333 131
rect 367 17 443 97
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
<< metal1 >>
rect 0 561 552 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 0 496 552 527
rect 0 17 552 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
rect 0 -48 552 -17
<< labels >>
rlabel locali s 298 199 379 265 6 A
port 1 nsew signal input
rlabel locali s 18 425 349 483 6 B
port 2 nsew signal input
rlabel locali s 122 199 264 323 6 C
port 3 nsew signal input
rlabel locali s 18 151 88 265 6 D
port 4 nsew signal input
rlabel metal1 s 0 -48 552 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 362 21 551 27 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 30 -17 64 27 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 27 551 163 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 362 163 551 203 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 590 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 552 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 481 83 535 152 6 X
port 9 nsew signal output
rlabel locali s 501 152 535 299 6 X
port 9 nsew signal output
rlabel locali s 481 299 535 493 6 X
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 552 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1054298
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1048276
<< end >>
