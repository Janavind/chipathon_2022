magic
tech sky130A
timestamp 1666199351
<< properties >>
string GDS_END 4360
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_2kbyte_1rw1r_32x512_8.gds
string GDS_START 3908
<< end >>
