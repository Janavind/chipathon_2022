magic
tech sky130A
magscale 1 2
timestamp 1666464484
<< nwell >>
rect -38 261 1694 582
<< pwell >>
rect 1 201 1341 203
rect 1 23 1652 201
rect 1 21 197 23
rect 655 21 845 23
rect 1256 21 1652 23
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 177
rect 186 93 216 177
rect 409 49 439 177
rect 497 49 527 177
rect 739 47 769 177
rect 925 49 955 177
rect 1076 49 1106 133
rect 1235 49 1265 177
rect 1355 47 1385 167
rect 1455 47 1485 175
rect 1539 47 1569 175
<< scpmoshvt >>
rect 83 297 113 497
rect 186 297 216 425
rect 396 325 426 493
rect 493 297 523 465
rect 705 297 735 497
rect 925 297 955 465
rect 1076 297 1106 425
rect 1251 329 1281 457
rect 1354 329 1384 497
rect 1455 297 1485 497
rect 1539 297 1569 497
<< ndiff >>
rect 27 129 79 177
rect 27 95 35 129
rect 69 95 79 129
rect 27 47 79 95
rect 109 93 186 177
rect 216 169 301 177
rect 216 135 255 169
rect 289 135 301 169
rect 216 93 301 135
rect 355 165 409 177
rect 355 131 365 165
rect 399 131 409 165
rect 109 89 171 93
rect 109 55 119 89
rect 153 55 171 89
rect 109 47 171 55
rect 355 49 409 131
rect 439 91 497 177
rect 439 57 451 91
rect 485 57 497 91
rect 439 49 497 57
rect 527 91 597 177
rect 527 57 551 91
rect 585 57 597 91
rect 527 49 597 57
rect 681 157 739 177
rect 681 123 695 157
rect 729 123 739 157
rect 681 89 739 123
rect 681 55 695 89
rect 729 55 739 89
rect 681 47 739 55
rect 769 165 821 177
rect 769 131 779 165
rect 813 131 821 165
rect 769 124 821 131
rect 769 47 819 124
rect 875 104 925 177
rect 873 97 925 104
rect 873 63 881 97
rect 915 63 925 97
rect 873 49 925 63
rect 955 133 1055 177
rect 1131 169 1235 177
rect 1131 135 1177 169
rect 1211 135 1235 169
rect 1131 133 1235 135
rect 955 126 1076 133
rect 955 92 965 126
rect 999 92 1076 126
rect 955 49 1076 92
rect 1106 49 1235 133
rect 1265 167 1315 177
rect 1405 167 1455 175
rect 1265 93 1355 167
rect 1265 59 1277 93
rect 1311 59 1355 93
rect 1265 49 1355 59
rect 1282 47 1355 49
rect 1385 142 1455 167
rect 1385 108 1411 142
rect 1445 108 1455 142
rect 1385 47 1455 108
rect 1485 97 1539 175
rect 1485 63 1495 97
rect 1529 63 1539 97
rect 1485 47 1539 63
rect 1569 101 1626 175
rect 1569 67 1579 101
rect 1613 67 1626 101
rect 1569 47 1626 67
<< pdiff >>
rect 27 477 83 497
rect 27 443 39 477
rect 73 443 83 477
rect 27 409 83 443
rect 27 375 39 409
rect 73 375 83 409
rect 27 341 83 375
rect 27 307 39 341
rect 73 307 83 341
rect 27 297 83 307
rect 113 477 171 497
rect 113 443 124 477
rect 158 443 171 477
rect 113 425 171 443
rect 113 297 186 425
rect 216 341 272 425
rect 216 307 226 341
rect 260 307 272 341
rect 331 413 396 493
rect 331 379 352 413
rect 386 379 396 413
rect 331 325 396 379
rect 426 481 478 493
rect 426 447 436 481
rect 470 465 478 481
rect 653 481 705 497
rect 470 447 493 465
rect 426 325 493 447
rect 216 297 272 307
rect 443 297 493 325
rect 523 423 599 465
rect 653 447 661 481
rect 695 447 705 481
rect 653 435 705 447
rect 523 339 600 423
rect 523 305 554 339
rect 588 305 600 339
rect 523 297 600 305
rect 654 297 705 435
rect 735 343 787 497
rect 735 309 745 343
rect 779 309 787 343
rect 735 297 787 309
rect 841 405 925 465
rect 841 371 849 405
rect 883 371 925 405
rect 841 297 925 371
rect 955 425 1054 465
rect 1296 489 1354 497
rect 1296 457 1308 489
rect 1166 425 1251 457
rect 955 409 1076 425
rect 955 375 1005 409
rect 1039 375 1076 409
rect 955 341 1076 375
rect 955 307 1005 341
rect 1039 307 1076 341
rect 955 297 1076 307
rect 1106 421 1251 425
rect 1106 387 1207 421
rect 1241 387 1251 421
rect 1106 329 1251 387
rect 1281 455 1308 457
rect 1342 455 1354 489
rect 1281 329 1354 455
rect 1384 341 1455 497
rect 1384 329 1411 341
rect 1106 297 1201 329
rect 1399 307 1411 329
rect 1445 307 1455 341
rect 1399 297 1455 307
rect 1485 489 1539 497
rect 1485 455 1495 489
rect 1529 455 1539 489
rect 1485 297 1539 455
rect 1569 477 1626 497
rect 1569 443 1580 477
rect 1614 443 1626 477
rect 1569 409 1626 443
rect 1569 375 1580 409
rect 1614 375 1626 409
rect 1569 297 1626 375
<< ndiffc >>
rect 35 95 69 129
rect 255 135 289 169
rect 365 131 399 165
rect 119 55 153 89
rect 451 57 485 91
rect 551 57 585 91
rect 695 123 729 157
rect 695 55 729 89
rect 779 131 813 165
rect 881 63 915 97
rect 1177 135 1211 169
rect 965 92 999 126
rect 1277 59 1311 93
rect 1411 108 1445 142
rect 1495 63 1529 97
rect 1579 67 1613 101
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 39 307 73 341
rect 124 443 158 477
rect 226 307 260 341
rect 352 379 386 413
rect 436 447 470 481
rect 661 447 695 481
rect 554 305 588 339
rect 745 309 779 343
rect 849 371 883 405
rect 1005 375 1039 409
rect 1005 307 1039 341
rect 1207 387 1241 421
rect 1308 455 1342 489
rect 1411 307 1445 341
rect 1495 455 1529 489
rect 1580 443 1614 477
rect 1580 375 1614 409
<< poly >>
rect 83 497 113 523
rect 396 493 426 519
rect 186 425 216 483
rect 493 465 523 504
rect 705 497 735 523
rect 83 265 113 297
rect 186 265 216 297
rect 396 271 426 325
rect 925 493 1281 523
rect 1354 497 1384 523
rect 1455 497 1485 523
rect 1539 497 1569 523
rect 925 465 955 493
rect 1251 457 1281 493
rect 1076 425 1106 451
rect 396 265 439 271
rect 493 265 523 297
rect 78 249 144 265
rect 78 215 100 249
rect 134 215 144 249
rect 78 199 144 215
rect 186 249 439 265
rect 186 215 366 249
rect 400 215 439 249
rect 186 199 439 215
rect 481 249 535 265
rect 481 215 491 249
rect 525 215 535 249
rect 705 247 735 297
rect 925 247 955 297
rect 1076 265 1106 297
rect 1251 265 1281 329
rect 705 217 955 247
rect 481 199 535 215
rect 79 177 109 199
rect 186 177 216 199
rect 409 177 439 199
rect 497 177 527 199
rect 739 177 769 217
rect 925 177 955 217
rect 997 249 1106 265
rect 997 215 1007 249
rect 1041 215 1106 249
rect 997 199 1106 215
rect 186 67 216 93
rect 79 21 109 47
rect 409 21 439 49
rect 497 21 527 49
rect 1076 133 1106 199
rect 1235 249 1289 265
rect 1354 256 1384 329
rect 1455 265 1485 297
rect 1539 265 1569 297
rect 1354 255 1385 256
rect 1235 215 1245 249
rect 1279 215 1289 249
rect 1235 199 1289 215
rect 1331 239 1385 255
rect 1331 205 1341 239
rect 1375 205 1385 239
rect 1235 177 1265 199
rect 1331 189 1385 205
rect 1427 249 1485 265
rect 1427 215 1437 249
rect 1471 215 1485 249
rect 1427 199 1485 215
rect 1527 249 1581 265
rect 1527 215 1537 249
rect 1571 215 1581 249
rect 1527 199 1581 215
rect 1355 167 1385 189
rect 1455 175 1485 199
rect 1539 175 1569 199
rect 739 21 769 47
rect 925 21 955 49
rect 1076 23 1106 49
rect 1235 21 1265 49
rect 1355 21 1385 47
rect 1455 21 1485 47
rect 1539 21 1569 47
<< polycont >>
rect 100 215 134 249
rect 366 215 400 249
rect 491 215 525 249
rect 1007 215 1041 249
rect 1245 215 1279 249
rect 1341 205 1375 239
rect 1437 215 1471 249
rect 1537 215 1571 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 17 477 73 493
rect 17 443 39 477
rect 107 477 174 527
rect 645 481 711 527
rect 1479 489 1546 527
rect 107 443 124 477
rect 158 443 174 477
rect 210 447 436 481
rect 470 447 504 481
rect 645 447 661 481
rect 695 447 711 481
rect 778 455 1308 489
rect 1342 455 1397 489
rect 1479 455 1495 489
rect 1529 455 1546 489
rect 1580 477 1639 493
rect 17 409 73 443
rect 210 409 244 447
rect 778 413 812 455
rect 17 375 39 409
rect 17 341 73 375
rect 17 307 39 341
rect 17 288 73 307
rect 107 375 244 409
rect 312 379 352 413
rect 386 379 812 413
rect 849 405 883 421
rect 17 185 66 288
rect 107 265 141 375
rect 187 307 226 341
rect 260 307 504 341
rect 100 249 141 265
rect 134 215 141 249
rect 100 199 141 215
rect 17 129 69 185
rect 106 173 141 199
rect 106 139 221 173
rect 17 95 35 129
rect 17 70 69 95
rect 103 89 153 105
rect 103 55 119 89
rect 103 17 153 55
rect 187 85 221 139
rect 255 169 289 307
rect 470 265 504 307
rect 538 305 554 339
rect 588 323 615 339
rect 559 289 581 305
rect 559 275 615 289
rect 323 249 436 265
rect 323 215 366 249
rect 400 215 436 249
rect 470 249 525 265
rect 470 215 491 249
rect 470 199 525 215
rect 255 119 289 135
rect 349 165 425 181
rect 349 131 365 165
rect 399 159 425 165
rect 559 159 593 275
rect 649 241 683 379
rect 729 309 745 343
rect 779 309 813 343
rect 729 289 813 309
rect 399 131 593 159
rect 349 125 593 131
rect 627 207 683 241
rect 627 91 661 207
rect 765 187 813 289
rect 414 85 451 91
rect 187 57 451 85
rect 485 57 501 91
rect 535 57 551 91
rect 585 57 661 91
rect 695 157 729 173
rect 695 89 729 123
rect 187 51 501 57
rect 799 165 813 187
rect 765 131 779 153
rect 765 83 813 131
rect 849 119 883 371
rect 917 178 951 455
rect 1614 443 1639 477
rect 1580 421 1639 443
rect 987 375 1005 409
rect 1039 375 1070 409
rect 987 341 1070 375
rect 987 307 1005 341
rect 1039 323 1070 341
rect 1177 387 1207 421
rect 1241 409 1639 421
rect 1241 387 1580 409
rect 1039 307 1041 323
rect 987 289 1041 307
rect 1075 289 1143 323
rect 990 249 1075 254
rect 990 215 1007 249
rect 1041 215 1075 249
rect 990 199 1075 215
rect 1033 187 1075 199
rect 917 165 959 178
rect 917 144 999 165
rect 925 131 999 144
rect 965 126 999 131
rect 1033 153 1041 187
rect 1033 126 1075 153
rect 849 85 857 119
rect 695 17 729 55
rect 849 63 881 85
rect 915 63 931 97
rect 965 64 999 92
rect 1109 85 1143 289
rect 1177 169 1211 387
rect 1542 375 1580 387
rect 1614 375 1639 409
rect 1245 289 1361 323
rect 1395 307 1411 341
rect 1445 307 1559 341
rect 1395 299 1559 307
rect 1245 249 1279 289
rect 1525 265 1559 299
rect 1245 199 1279 215
rect 1313 239 1375 255
rect 1313 205 1341 239
rect 1409 249 1491 265
rect 1409 215 1437 249
rect 1471 215 1491 249
rect 1525 249 1571 265
rect 1525 215 1537 249
rect 1313 189 1375 205
rect 1525 199 1571 215
rect 1313 187 1354 189
rect 1313 153 1317 187
rect 1351 153 1354 187
rect 1525 181 1559 199
rect 1313 146 1354 153
rect 1411 150 1559 181
rect 1403 147 1559 150
rect 1177 119 1211 135
rect 1403 142 1461 147
rect 1403 119 1411 142
rect 1245 85 1277 93
rect 849 53 931 63
rect 1109 59 1277 85
rect 1311 59 1338 93
rect 1403 85 1409 119
rect 1445 108 1461 142
rect 1605 117 1639 375
rect 1443 85 1461 108
rect 1403 59 1461 85
rect 1495 97 1529 113
rect 1109 51 1338 59
rect 1495 17 1529 63
rect 1579 101 1639 117
rect 1613 67 1639 101
rect 1579 51 1639 67
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 581 305 588 323
rect 588 305 615 323
rect 581 289 615 305
rect 765 165 799 187
rect 765 153 779 165
rect 779 153 799 165
rect 1041 289 1075 323
rect 1041 153 1075 187
rect 857 97 891 119
rect 857 85 881 97
rect 881 85 891 97
rect 1317 153 1351 187
rect 1409 108 1411 119
rect 1411 108 1443 119
rect 1409 85 1443 108
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
<< metal1 >>
rect 0 561 1656 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 0 496 1656 527
rect 569 323 627 329
rect 569 289 581 323
rect 615 320 627 323
rect 1029 323 1087 329
rect 1029 320 1041 323
rect 615 292 1041 320
rect 615 289 627 292
rect 569 283 627 289
rect 1029 289 1041 292
rect 1075 289 1087 323
rect 1029 283 1087 289
rect 753 187 811 193
rect 753 153 765 187
rect 799 184 811 187
rect 1029 187 1087 193
rect 1029 184 1041 187
rect 799 156 1041 184
rect 799 153 811 156
rect 753 147 811 153
rect 1029 153 1041 156
rect 1075 184 1087 187
rect 1305 187 1363 193
rect 1305 184 1317 187
rect 1075 156 1317 184
rect 1075 153 1087 156
rect 1029 147 1087 153
rect 1305 153 1317 156
rect 1351 153 1363 187
rect 1305 147 1363 153
rect 845 119 903 125
rect 845 85 857 119
rect 891 116 903 119
rect 1397 119 1455 125
rect 1397 116 1409 119
rect 891 88 1409 116
rect 891 85 903 88
rect 845 79 903 85
rect 1397 85 1409 88
rect 1443 85 1455 119
rect 1397 79 1455 85
rect 0 17 1656 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
rect 0 -48 1656 -17
<< labels >>
flabel locali s 29 357 63 391 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 1317 289 1351 323 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 397 221 431 255 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 1409 221 1443 255 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 xnor3_1
rlabel metal1 s 0 -48 1656 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1656 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1656 544
string GDS_END 596416
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 584810
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 8.280 0.000 
<< end >>
