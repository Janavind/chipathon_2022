magic
tech sky130A
magscale 1 2
timestamp 1666464484
use sky130_fd_pr__dfl1sd2__example_55959141808518  sky130_fd_pr__dfl1sd2__example_55959141808518_0
timestamp 1666464484
transform 1 0 160 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808518  sky130_fd_pr__dfl1sd2__example_55959141808518_1
timestamp 1666464484
transform 1 0 376 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808518  sky130_fd_pr__dfl1sd2__example_55959141808518_2
timestamp 1666464484
transform 1 0 592 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808518  sky130_fd_pr__dfl1sd2__example_55959141808518_3
timestamp 1666464484
transform 1 0 808 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808518  sky130_fd_pr__dfl1sd2__example_55959141808518_4
timestamp 1666464484
transform 1 0 1024 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_55959141808517  sky130_fd_pr__dfl1sd__example_55959141808517_0
timestamp 1666464484
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_55959141808517  sky130_fd_pr__dfl1sd__example_55959141808517_1
timestamp 1666464484
transform 1 0 1240 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 42402304
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 42398802
<< end >>
