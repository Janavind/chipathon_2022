magic
tech sky130B
magscale 1 2
timestamp 1666199351
<< locali >>
rect 383 1369 667 1388
rect 383 1263 400 1369
rect 650 1263 667 1369
rect 383 1251 667 1263
rect 383 125 667 137
rect 383 19 400 125
rect 650 19 667 125
rect 383 0 667 19
<< viali >>
rect 400 1263 650 1369
rect 400 19 650 125
<< obsli1 >>
rect 190 1225 256 1291
rect 794 1225 860 1291
rect 190 1203 230 1225
rect 820 1203 860 1225
rect 41 1179 230 1203
rect 41 1145 60 1179
rect 94 1145 230 1179
rect 41 1107 230 1145
rect 41 1073 60 1107
rect 94 1073 230 1107
rect 41 1035 230 1073
rect 41 1001 60 1035
rect 94 1001 230 1035
rect 41 963 230 1001
rect 41 929 60 963
rect 94 929 230 963
rect 41 891 230 929
rect 41 857 60 891
rect 94 857 230 891
rect 41 819 230 857
rect 41 785 60 819
rect 94 785 230 819
rect 41 747 230 785
rect 41 713 60 747
rect 94 713 230 747
rect 41 675 230 713
rect 41 641 60 675
rect 94 641 230 675
rect 41 603 230 641
rect 41 569 60 603
rect 94 569 230 603
rect 41 531 230 569
rect 41 497 60 531
rect 94 497 230 531
rect 41 459 230 497
rect 41 425 60 459
rect 94 425 230 459
rect 41 387 230 425
rect 41 353 60 387
rect 94 353 230 387
rect 41 315 230 353
rect 41 281 60 315
rect 94 281 230 315
rect 41 243 230 281
rect 41 209 60 243
rect 94 209 230 243
rect 41 185 230 209
rect 352 185 386 1203
rect 508 185 542 1203
rect 664 185 698 1203
rect 820 1179 1009 1203
rect 820 1145 956 1179
rect 990 1145 1009 1179
rect 820 1107 1009 1145
rect 820 1073 956 1107
rect 990 1073 1009 1107
rect 820 1035 1009 1073
rect 820 1001 956 1035
rect 990 1001 1009 1035
rect 820 963 1009 1001
rect 820 929 956 963
rect 990 929 1009 963
rect 820 891 1009 929
rect 820 857 956 891
rect 990 857 1009 891
rect 820 819 1009 857
rect 820 785 956 819
rect 990 785 1009 819
rect 820 747 1009 785
rect 820 713 956 747
rect 990 713 1009 747
rect 820 675 1009 713
rect 820 641 956 675
rect 990 641 1009 675
rect 820 603 1009 641
rect 820 569 956 603
rect 990 569 1009 603
rect 820 531 1009 569
rect 820 497 956 531
rect 990 497 1009 531
rect 820 459 1009 497
rect 820 425 956 459
rect 990 425 1009 459
rect 820 387 1009 425
rect 820 353 956 387
rect 990 353 1009 387
rect 820 315 1009 353
rect 820 281 956 315
rect 990 281 1009 315
rect 820 243 1009 281
rect 820 209 956 243
rect 990 209 1009 243
rect 820 185 1009 209
rect 190 163 230 185
rect 820 163 860 185
rect 190 97 256 163
rect 794 97 860 163
<< obsli1c >>
rect 60 1145 94 1179
rect 60 1073 94 1107
rect 60 1001 94 1035
rect 60 929 94 963
rect 60 857 94 891
rect 60 785 94 819
rect 60 713 94 747
rect 60 641 94 675
rect 60 569 94 603
rect 60 497 94 531
rect 60 425 94 459
rect 60 353 94 387
rect 60 281 94 315
rect 60 209 94 243
rect 956 1145 990 1179
rect 956 1073 990 1107
rect 956 1001 990 1035
rect 956 929 990 963
rect 956 857 990 891
rect 956 785 990 819
rect 956 713 990 747
rect 956 641 990 675
rect 956 569 990 603
rect 956 497 990 531
rect 956 425 990 459
rect 956 353 990 387
rect 956 281 990 315
rect 956 209 990 243
<< metal1 >>
rect 380 1369 670 1388
rect 380 1263 400 1369
rect 650 1263 670 1369
rect 380 1251 670 1263
rect 41 1179 100 1191
rect 41 1145 60 1179
rect 94 1145 100 1179
rect 41 1107 100 1145
rect 41 1073 60 1107
rect 94 1073 100 1107
rect 41 1035 100 1073
rect 41 1001 60 1035
rect 94 1001 100 1035
rect 41 963 100 1001
rect 41 929 60 963
rect 94 929 100 963
rect 41 891 100 929
rect 41 857 60 891
rect 94 857 100 891
rect 41 819 100 857
rect 41 785 60 819
rect 94 785 100 819
rect 41 747 100 785
rect 41 713 60 747
rect 94 713 100 747
rect 41 675 100 713
rect 41 641 60 675
rect 94 641 100 675
rect 41 603 100 641
rect 41 569 60 603
rect 94 569 100 603
rect 41 531 100 569
rect 41 497 60 531
rect 94 497 100 531
rect 41 459 100 497
rect 41 425 60 459
rect 94 425 100 459
rect 41 387 100 425
rect 41 353 60 387
rect 94 353 100 387
rect 41 315 100 353
rect 41 281 60 315
rect 94 281 100 315
rect 41 243 100 281
rect 41 209 60 243
rect 94 209 100 243
rect 41 197 100 209
rect 950 1179 1009 1191
rect 950 1145 956 1179
rect 990 1145 1009 1179
rect 950 1107 1009 1145
rect 950 1073 956 1107
rect 990 1073 1009 1107
rect 950 1035 1009 1073
rect 950 1001 956 1035
rect 990 1001 1009 1035
rect 950 963 1009 1001
rect 950 929 956 963
rect 990 929 1009 963
rect 950 891 1009 929
rect 950 857 956 891
rect 990 857 1009 891
rect 950 819 1009 857
rect 950 785 956 819
rect 990 785 1009 819
rect 950 747 1009 785
rect 950 713 956 747
rect 990 713 1009 747
rect 950 675 1009 713
rect 950 641 956 675
rect 990 641 1009 675
rect 950 603 1009 641
rect 950 569 956 603
rect 990 569 1009 603
rect 950 531 1009 569
rect 950 497 956 531
rect 990 497 1009 531
rect 950 459 1009 497
rect 950 425 956 459
rect 990 425 1009 459
rect 950 387 1009 425
rect 950 353 956 387
rect 990 353 1009 387
rect 950 315 1009 353
rect 950 281 956 315
rect 990 281 1009 315
rect 950 243 1009 281
rect 950 209 956 243
rect 990 209 1009 243
rect 950 197 1009 209
rect 380 125 670 137
rect 380 19 400 125
rect 650 19 670 125
rect 380 0 670 19
<< obsm1 >>
rect 343 197 395 1191
rect 499 197 551 1191
rect 655 197 707 1191
<< metal2 >>
rect 14 719 1036 1191
rect 14 197 1036 669
<< labels >>
rlabel metal2 s 14 719 1036 1191 6 DRAIN
port 1 nsew
rlabel viali s 400 1263 650 1369 6 GATE
port 2 nsew
rlabel viali s 400 19 650 125 6 GATE
port 2 nsew
rlabel locali s 383 1251 667 1388 6 GATE
port 2 nsew
rlabel locali s 383 0 667 137 6 GATE
port 2 nsew
rlabel metal1 s 380 1251 670 1388 6 GATE
port 2 nsew
rlabel metal1 s 380 0 670 137 6 GATE
port 2 nsew
rlabel metal2 s 14 197 1036 669 6 SOURCE
port 3 nsew
rlabel metal1 s 41 197 100 1191 6 SUBSTRATE
port 4 nsew
rlabel metal1 s 950 197 1009 1191 6 SUBSTRATE
port 4 nsew
<< properties >>
string FIXED_BBOX 14 0 1036 1388
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 8463040
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 8440388
string device primitive
<< end >>
