magic
tech sky130A
magscale 1 2
timestamp 1666199351
<< nwell >>
rect -36 679 1808 1471
<< pwell >>
rect 1636 25 1738 159
<< psubdiff >>
rect 1662 109 1712 133
rect 1662 75 1670 109
rect 1704 75 1712 109
rect 1662 51 1712 75
<< nsubdiff >>
rect 1662 1339 1712 1363
rect 1662 1305 1670 1339
rect 1704 1305 1712 1339
rect 1662 1281 1712 1305
<< psubdiffcont >>
rect 1670 75 1704 109
<< nsubdiffcont >>
rect 1670 1305 1704 1339
<< poly >>
rect 114 740 144 907
rect 48 724 144 740
rect 48 690 64 724
rect 98 690 144 724
rect 48 674 144 690
rect 114 507 144 674
<< polycont >>
rect 64 690 98 724
<< locali >>
rect 0 1397 1772 1431
rect 62 1130 96 1397
rect 274 1130 308 1397
rect 490 1130 524 1397
rect 706 1130 740 1397
rect 922 1130 956 1397
rect 1138 1130 1172 1397
rect 1354 1130 1388 1397
rect 1566 1130 1600 1397
rect 1670 1339 1704 1397
rect 1670 1289 1704 1305
rect 64 724 98 740
rect 64 674 98 690
rect 814 724 848 1096
rect 814 690 865 724
rect 814 318 848 690
rect 62 17 96 218
rect 274 17 308 218
rect 490 17 524 218
rect 706 17 740 218
rect 922 17 956 218
rect 1138 17 1172 218
rect 1354 17 1388 218
rect 1566 17 1600 218
rect 1670 109 1704 125
rect 1670 17 1704 75
rect 0 -17 1772 17
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_16  sky130_sram_2kbyte_1rw1r_32x512_8_contact_16_0
timestamp 1666199351
transform 1 0 48 0 1 674
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_28  sky130_sram_2kbyte_1rw1r_32x512_8_contact_28_0
timestamp 1666199351
transform 1 0 1662 0 1 1281
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_29  sky130_sram_2kbyte_1rw1r_32x512_8_contact_29_0
timestamp 1666199351
transform 1 0 1662 0 1 51
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_nmos_m14_w2_000_sli_dli_da_p  sky130_sram_2kbyte_1rw1r_32x512_8_nmos_m14_w2_000_sli_dli_da_p_0
timestamp 1666199351
transform 1 0 54 0 1 51
box -26 -26 1580 456
use sky130_sram_2kbyte_1rw1r_32x512_8_pmos_m14_w2_000_sli_dli_da_p  sky130_sram_2kbyte_1rw1r_32x512_8_pmos_m14_w2_000_sli_dli_da_p_0
timestamp 1666199351
transform 1 0 54 0 1 963
box -59 -56 1613 454
<< labels >>
rlabel locali s 81 707 81 707 4 A
port 1 nsew
rlabel locali s 848 707 848 707 4 Z
port 2 nsew
rlabel locali s 886 0 886 0 4 gnd
port 3 nsew
rlabel locali s 886 1414 886 1414 4 vdd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 1772 1414
string GDS_END 360640
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_2kbyte_1rw1r_32x512_8.gds
string GDS_START 357874
<< end >>
