magic
tech sky130B
magscale 1 2
timestamp 1666199351
<< locali >>
rect 1935 8820 1969 8836
rect 1935 8770 1969 8786
rect 11919 8820 11953 8836
rect 11919 8770 11953 8786
rect 21903 8820 21937 8836
rect 21903 8770 21937 8786
rect 31887 8820 31921 8836
rect 31887 8770 31921 8786
<< viali >>
rect 1935 8786 1969 8820
rect 11919 8786 11953 8820
rect 21903 8786 21937 8820
rect 31887 8786 31921 8820
<< metal1 >>
rect 1923 8820 1981 8826
rect 1923 8786 1935 8820
rect 1969 8817 1981 8820
rect 10717 8817 10723 8829
rect 1969 8789 10723 8817
rect 1969 8786 1981 8789
rect 1923 8780 1981 8786
rect 10717 8777 10723 8789
rect 10775 8777 10781 8829
rect 11907 8820 11965 8826
rect 11907 8786 11919 8820
rect 11953 8817 11965 8820
rect 20701 8817 20707 8829
rect 11953 8789 20707 8817
rect 11953 8786 11965 8789
rect 11907 8780 11965 8786
rect 20701 8777 20707 8789
rect 20759 8777 20765 8829
rect 21891 8820 21949 8826
rect 21891 8786 21903 8820
rect 21937 8817 21949 8820
rect 30685 8817 30691 8829
rect 21937 8789 30691 8817
rect 21937 8786 21949 8789
rect 21891 8780 21949 8786
rect 30685 8777 30691 8789
rect 30743 8777 30749 8829
rect 31875 8820 31933 8826
rect 31875 8786 31887 8820
rect 31921 8817 31933 8820
rect 40669 8817 40675 8829
rect 31921 8789 40675 8817
rect 31921 8786 31933 8789
rect 31875 8780 31933 8786
rect 40669 8777 40675 8789
rect 40727 8777 40733 8829
rect 1629 7905 1689 7961
rect 2877 7905 2937 7961
rect 4125 7905 4185 7961
rect 5373 7905 5433 7961
rect 6621 7905 6681 7961
rect 7869 7905 7929 7961
rect 9117 7905 9177 7961
rect 10365 7905 10425 7961
rect 11613 7905 11673 7961
rect 12861 7905 12921 7961
rect 14109 7905 14169 7961
rect 15357 7905 15417 7961
rect 16605 7905 16665 7961
rect 17853 7905 17913 7961
rect 19101 7905 19161 7961
rect 20349 7905 20409 7961
rect 21597 7905 21657 7961
rect 22845 7905 22905 7961
rect 24093 7905 24153 7961
rect 25341 7905 25401 7961
rect 26589 7905 26649 7961
rect 27837 7905 27897 7961
rect 29085 7905 29145 7961
rect 30333 7905 30393 7961
rect 31581 7905 31641 7961
rect 32829 7905 32889 7961
rect 34077 7905 34137 7961
rect 35325 7905 35385 7961
rect 36573 7905 36633 7961
rect 37821 7905 37881 7961
rect 39069 7905 39129 7961
rect 40317 7905 40377 7961
rect 10717 7871 10723 7880
rect 1473 7837 10723 7871
rect 10717 7828 10723 7837
rect 10775 7871 10781 7880
rect 20701 7871 20707 7880
rect 10775 7837 10833 7871
rect 11457 7837 20707 7871
rect 10775 7828 10781 7837
rect 20701 7828 20707 7837
rect 20759 7871 20765 7880
rect 30685 7871 30691 7880
rect 20759 7837 20817 7871
rect 21441 7837 30691 7871
rect 20759 7828 20765 7837
rect 30685 7828 30691 7837
rect 30743 7871 30749 7880
rect 40669 7871 40675 7880
rect 30743 7837 30801 7871
rect 31425 7837 40675 7871
rect 30743 7828 30749 7837
rect 40669 7828 40675 7837
rect 40727 7871 40733 7880
rect 40727 7837 40785 7871
rect 40727 7828 40733 7837
rect 1501 5888 1529 5954
rect 1501 5860 1601 5888
rect 1478 5448 1524 5702
rect 1573 4572 1601 5860
rect 1703 5808 1731 5954
rect 2749 5888 2777 5954
rect 2749 5860 2849 5888
rect 1646 5780 1731 5808
rect 1646 4560 1674 5780
rect 2726 5448 2772 5702
rect 2821 4572 2849 5860
rect 2951 5808 2979 5954
rect 3997 5888 4025 5954
rect 3997 5860 4097 5888
rect 2894 5780 2979 5808
rect 2894 4560 2922 5780
rect 3974 5448 4020 5702
rect 4069 4572 4097 5860
rect 4199 5808 4227 5954
rect 5245 5888 5273 5954
rect 5245 5860 5345 5888
rect 4142 5780 4227 5808
rect 4142 4560 4170 5780
rect 5222 5448 5268 5702
rect 5317 4572 5345 5860
rect 5447 5808 5475 5954
rect 6493 5888 6521 5954
rect 6493 5860 6593 5888
rect 5390 5780 5475 5808
rect 5390 4560 5418 5780
rect 6470 5448 6516 5702
rect 6565 4572 6593 5860
rect 6695 5808 6723 5954
rect 7741 5888 7769 5954
rect 7741 5860 7841 5888
rect 6638 5780 6723 5808
rect 6638 4560 6666 5780
rect 7718 5448 7764 5702
rect 7813 4572 7841 5860
rect 7943 5808 7971 5954
rect 8989 5888 9017 5954
rect 8989 5860 9089 5888
rect 7886 5780 7971 5808
rect 7886 4560 7914 5780
rect 8966 5448 9012 5702
rect 9061 4572 9089 5860
rect 9191 5808 9219 5954
rect 10237 5888 10265 5954
rect 10237 5860 10337 5888
rect 9134 5780 9219 5808
rect 9134 4560 9162 5780
rect 10214 5448 10260 5702
rect 10309 4572 10337 5860
rect 10439 5808 10467 5954
rect 11485 5888 11513 5954
rect 11485 5860 11585 5888
rect 10382 5780 10467 5808
rect 10382 4560 10410 5780
rect 11462 5448 11508 5702
rect 11557 4572 11585 5860
rect 11687 5808 11715 5954
rect 12733 5888 12761 5954
rect 12733 5860 12833 5888
rect 11630 5780 11715 5808
rect 11630 4560 11658 5780
rect 12710 5448 12756 5702
rect 12805 4572 12833 5860
rect 12935 5808 12963 5954
rect 13981 5888 14009 5954
rect 13981 5860 14081 5888
rect 12878 5780 12963 5808
rect 12878 4560 12906 5780
rect 13958 5448 14004 5702
rect 14053 4572 14081 5860
rect 14183 5808 14211 5954
rect 15229 5888 15257 5954
rect 15229 5860 15329 5888
rect 14126 5780 14211 5808
rect 14126 4560 14154 5780
rect 15206 5448 15252 5702
rect 15301 4572 15329 5860
rect 15431 5808 15459 5954
rect 16477 5888 16505 5954
rect 16477 5860 16577 5888
rect 15374 5780 15459 5808
rect 15374 4560 15402 5780
rect 16454 5448 16500 5702
rect 16549 4572 16577 5860
rect 16679 5808 16707 5954
rect 17725 5888 17753 5954
rect 17725 5860 17825 5888
rect 16622 5780 16707 5808
rect 16622 4560 16650 5780
rect 17702 5448 17748 5702
rect 17797 4572 17825 5860
rect 17927 5808 17955 5954
rect 18973 5888 19001 5954
rect 18973 5860 19073 5888
rect 17870 5780 17955 5808
rect 17870 4560 17898 5780
rect 18950 5448 18996 5702
rect 19045 4572 19073 5860
rect 19175 5808 19203 5954
rect 20221 5888 20249 5954
rect 20221 5860 20321 5888
rect 19118 5780 19203 5808
rect 19118 4560 19146 5780
rect 20198 5448 20244 5702
rect 20293 4572 20321 5860
rect 20423 5808 20451 5954
rect 21469 5888 21497 5954
rect 21469 5860 21569 5888
rect 20366 5780 20451 5808
rect 20366 4560 20394 5780
rect 21446 5448 21492 5702
rect 21541 4572 21569 5860
rect 21671 5808 21699 5954
rect 22717 5888 22745 5954
rect 22717 5860 22817 5888
rect 21614 5780 21699 5808
rect 21614 4560 21642 5780
rect 22694 5448 22740 5702
rect 22789 4572 22817 5860
rect 22919 5808 22947 5954
rect 23965 5888 23993 5954
rect 23965 5860 24065 5888
rect 22862 5780 22947 5808
rect 22862 4560 22890 5780
rect 23942 5448 23988 5702
rect 24037 4572 24065 5860
rect 24167 5808 24195 5954
rect 25213 5888 25241 5954
rect 25213 5860 25313 5888
rect 24110 5780 24195 5808
rect 24110 4560 24138 5780
rect 25190 5448 25236 5702
rect 25285 4572 25313 5860
rect 25415 5808 25443 5954
rect 26461 5888 26489 5954
rect 26461 5860 26561 5888
rect 25358 5780 25443 5808
rect 25358 4560 25386 5780
rect 26438 5448 26484 5702
rect 26533 4572 26561 5860
rect 26663 5808 26691 5954
rect 27709 5888 27737 5954
rect 27709 5860 27809 5888
rect 26606 5780 26691 5808
rect 26606 4560 26634 5780
rect 27686 5448 27732 5702
rect 27781 4572 27809 5860
rect 27911 5808 27939 5954
rect 28957 5888 28985 5954
rect 28957 5860 29057 5888
rect 27854 5780 27939 5808
rect 27854 4560 27882 5780
rect 28934 5448 28980 5702
rect 29029 4572 29057 5860
rect 29159 5808 29187 5954
rect 30205 5888 30233 5954
rect 30205 5860 30305 5888
rect 29102 5780 29187 5808
rect 29102 4560 29130 5780
rect 30182 5448 30228 5702
rect 30277 4572 30305 5860
rect 30407 5808 30435 5954
rect 31453 5888 31481 5954
rect 31453 5860 31553 5888
rect 30350 5780 30435 5808
rect 30350 4560 30378 5780
rect 31430 5448 31476 5702
rect 31525 4572 31553 5860
rect 31655 5808 31683 5954
rect 32701 5888 32729 5954
rect 32701 5860 32801 5888
rect 31598 5780 31683 5808
rect 31598 4560 31626 5780
rect 32678 5448 32724 5702
rect 32773 4572 32801 5860
rect 32903 5808 32931 5954
rect 33949 5888 33977 5954
rect 33949 5860 34049 5888
rect 32846 5780 32931 5808
rect 32846 4560 32874 5780
rect 33926 5448 33972 5702
rect 34021 4572 34049 5860
rect 34151 5808 34179 5954
rect 35197 5888 35225 5954
rect 35197 5860 35297 5888
rect 34094 5780 34179 5808
rect 34094 4560 34122 5780
rect 35174 5448 35220 5702
rect 35269 4572 35297 5860
rect 35399 5808 35427 5954
rect 36445 5888 36473 5954
rect 36445 5860 36545 5888
rect 35342 5780 35427 5808
rect 35342 4560 35370 5780
rect 36422 5448 36468 5702
rect 36517 4572 36545 5860
rect 36647 5808 36675 5954
rect 37693 5888 37721 5954
rect 37693 5860 37793 5888
rect 36590 5780 36675 5808
rect 36590 4560 36618 5780
rect 37670 5448 37716 5702
rect 37765 4572 37793 5860
rect 37895 5808 37923 5954
rect 38941 5888 38969 5954
rect 38941 5860 39041 5888
rect 37838 5780 37923 5808
rect 37838 4560 37866 5780
rect 38918 5448 38964 5702
rect 39013 4572 39041 5860
rect 39143 5808 39171 5954
rect 40189 5888 40217 5954
rect 40189 5860 40289 5888
rect 39086 5780 39171 5808
rect 39086 4560 39114 5780
rect 40166 5448 40212 5702
rect 40261 4572 40289 5860
rect 40391 5808 40419 5954
rect 40334 5780 40419 5808
rect 40334 4560 40362 5780
rect 1573 3380 1601 3446
rect 1454 3352 1601 3380
rect 1454 2946 1482 3352
rect 1646 3300 1674 3446
rect 2821 3380 2849 3446
rect 2702 3352 2849 3380
rect 1646 3272 1946 3300
rect 1918 3070 1946 3272
rect 2702 2946 2730 3352
rect 2894 3300 2922 3446
rect 4069 3380 4097 3446
rect 3950 3352 4097 3380
rect 2894 3272 3194 3300
rect 3166 3070 3194 3272
rect 3950 2946 3978 3352
rect 4142 3300 4170 3446
rect 5317 3380 5345 3446
rect 5198 3352 5345 3380
rect 4142 3272 4442 3300
rect 4414 3070 4442 3272
rect 5198 2946 5226 3352
rect 5390 3300 5418 3446
rect 6565 3380 6593 3446
rect 6446 3352 6593 3380
rect 5390 3272 5690 3300
rect 5662 3070 5690 3272
rect 6446 2946 6474 3352
rect 6638 3300 6666 3446
rect 7813 3380 7841 3446
rect 7694 3352 7841 3380
rect 6638 3272 6938 3300
rect 6910 3070 6938 3272
rect 7694 2946 7722 3352
rect 7886 3300 7914 3446
rect 9061 3380 9089 3446
rect 8942 3352 9089 3380
rect 7886 3272 8186 3300
rect 8158 3070 8186 3272
rect 8942 2946 8970 3352
rect 9134 3300 9162 3446
rect 10309 3380 10337 3446
rect 10190 3352 10337 3380
rect 9134 3272 9434 3300
rect 9406 3070 9434 3272
rect 10190 2946 10218 3352
rect 10382 3300 10410 3446
rect 11557 3380 11585 3446
rect 11438 3352 11585 3380
rect 10382 3272 10682 3300
rect 10654 3070 10682 3272
rect 11438 2946 11466 3352
rect 11630 3300 11658 3446
rect 12805 3380 12833 3446
rect 12686 3352 12833 3380
rect 11630 3272 11930 3300
rect 11902 3070 11930 3272
rect 12686 2946 12714 3352
rect 12878 3300 12906 3446
rect 14053 3380 14081 3446
rect 13934 3352 14081 3380
rect 12878 3272 13178 3300
rect 13150 3070 13178 3272
rect 13934 2946 13962 3352
rect 14126 3300 14154 3446
rect 15301 3380 15329 3446
rect 15182 3352 15329 3380
rect 14126 3272 14426 3300
rect 14398 3070 14426 3272
rect 15182 2946 15210 3352
rect 15374 3300 15402 3446
rect 16549 3380 16577 3446
rect 16430 3352 16577 3380
rect 15374 3272 15674 3300
rect 15646 3070 15674 3272
rect 16430 2946 16458 3352
rect 16622 3300 16650 3446
rect 17797 3380 17825 3446
rect 17678 3352 17825 3380
rect 16622 3272 16922 3300
rect 16894 3070 16922 3272
rect 17678 2946 17706 3352
rect 17870 3300 17898 3446
rect 19045 3380 19073 3446
rect 18926 3352 19073 3380
rect 17870 3272 18170 3300
rect 18142 3070 18170 3272
rect 18926 2946 18954 3352
rect 19118 3300 19146 3446
rect 20293 3380 20321 3446
rect 20174 3352 20321 3380
rect 19118 3272 19418 3300
rect 19390 3070 19418 3272
rect 20174 2946 20202 3352
rect 20366 3300 20394 3446
rect 21541 3380 21569 3446
rect 21422 3352 21569 3380
rect 20366 3272 20666 3300
rect 20638 3070 20666 3272
rect 21422 2946 21450 3352
rect 21614 3300 21642 3446
rect 22789 3380 22817 3446
rect 22670 3352 22817 3380
rect 21614 3272 21914 3300
rect 21886 3070 21914 3272
rect 22670 2946 22698 3352
rect 22862 3300 22890 3446
rect 24037 3380 24065 3446
rect 23918 3352 24065 3380
rect 22862 3272 23162 3300
rect 23134 3070 23162 3272
rect 23918 2946 23946 3352
rect 24110 3300 24138 3446
rect 25285 3380 25313 3446
rect 25166 3352 25313 3380
rect 24110 3272 24410 3300
rect 24382 3070 24410 3272
rect 25166 2946 25194 3352
rect 25358 3300 25386 3446
rect 26533 3380 26561 3446
rect 26414 3352 26561 3380
rect 25358 3272 25658 3300
rect 25630 3070 25658 3272
rect 26414 2946 26442 3352
rect 26606 3300 26634 3446
rect 27781 3380 27809 3446
rect 27662 3352 27809 3380
rect 26606 3272 26906 3300
rect 26878 3070 26906 3272
rect 27662 2946 27690 3352
rect 27854 3300 27882 3446
rect 29029 3380 29057 3446
rect 28910 3352 29057 3380
rect 27854 3272 28154 3300
rect 28126 3070 28154 3272
rect 28910 2946 28938 3352
rect 29102 3300 29130 3446
rect 30277 3380 30305 3446
rect 30158 3352 30305 3380
rect 29102 3272 29402 3300
rect 29374 3070 29402 3272
rect 30158 2946 30186 3352
rect 30350 3300 30378 3446
rect 31525 3380 31553 3446
rect 31406 3352 31553 3380
rect 30350 3272 30650 3300
rect 30622 3070 30650 3272
rect 31406 2946 31434 3352
rect 31598 3300 31626 3446
rect 32773 3380 32801 3446
rect 32654 3352 32801 3380
rect 31598 3272 31898 3300
rect 31870 3070 31898 3272
rect 32654 2946 32682 3352
rect 32846 3300 32874 3446
rect 34021 3380 34049 3446
rect 33902 3352 34049 3380
rect 32846 3272 33146 3300
rect 33118 3070 33146 3272
rect 33902 2946 33930 3352
rect 34094 3300 34122 3446
rect 35269 3380 35297 3446
rect 35150 3352 35297 3380
rect 34094 3272 34394 3300
rect 34366 3070 34394 3272
rect 35150 2946 35178 3352
rect 35342 3300 35370 3446
rect 36517 3380 36545 3446
rect 36398 3352 36545 3380
rect 35342 3272 35642 3300
rect 35614 3070 35642 3272
rect 36398 2946 36426 3352
rect 36590 3300 36618 3446
rect 37765 3380 37793 3446
rect 37646 3352 37793 3380
rect 36590 3272 36890 3300
rect 36862 3070 36890 3272
rect 37646 2946 37674 3352
rect 37838 3300 37866 3446
rect 39013 3380 39041 3446
rect 38894 3352 39041 3380
rect 37838 3272 38138 3300
rect 38110 3070 38138 3272
rect 38894 2946 38922 3352
rect 39086 3300 39114 3446
rect 40261 3380 40289 3446
rect 40142 3352 40289 3380
rect 39086 3272 39386 3300
rect 39358 3070 39386 3272
rect 40142 2946 40170 3352
rect 40334 3300 40362 3446
rect 40334 3272 40634 3300
rect 40606 3070 40634 3272
rect 1454 1192 1482 1258
rect 1440 1164 1482 1192
rect 816 252 844 1006
rect 1280 252 1308 1006
rect 1440 252 1468 1164
rect 1918 1112 1946 1258
rect 1904 1084 1946 1112
rect 2050 1112 2078 1258
rect 2514 1192 2542 1258
rect 2702 1192 2730 1258
rect 2514 1164 2556 1192
rect 2050 1084 2092 1112
rect 1904 252 1932 1084
rect 2064 252 2092 1084
rect 2528 252 2556 1164
rect 2688 1164 2730 1192
rect 2688 252 2716 1164
rect 3166 1112 3194 1258
rect 3152 1084 3194 1112
rect 3298 1112 3326 1258
rect 3762 1192 3790 1258
rect 3950 1192 3978 1258
rect 3762 1164 3804 1192
rect 3298 1084 3340 1112
rect 3152 252 3180 1084
rect 3312 252 3340 1084
rect 3776 252 3804 1164
rect 3936 1164 3978 1192
rect 3936 252 3964 1164
rect 4414 1112 4442 1258
rect 4400 1084 4442 1112
rect 4546 1112 4574 1258
rect 5010 1192 5038 1258
rect 5198 1192 5226 1258
rect 5010 1164 5052 1192
rect 4546 1084 4588 1112
rect 4400 252 4428 1084
rect 4560 252 4588 1084
rect 5024 252 5052 1164
rect 5184 1164 5226 1192
rect 5184 252 5212 1164
rect 5662 1112 5690 1258
rect 5648 1084 5690 1112
rect 5794 1112 5822 1258
rect 6258 1192 6286 1258
rect 6446 1192 6474 1258
rect 6258 1164 6300 1192
rect 5794 1084 5836 1112
rect 5648 252 5676 1084
rect 5808 252 5836 1084
rect 6272 252 6300 1164
rect 6432 1164 6474 1192
rect 6432 252 6460 1164
rect 6910 1112 6938 1258
rect 6896 1084 6938 1112
rect 7042 1112 7070 1258
rect 7506 1192 7534 1258
rect 7694 1192 7722 1258
rect 7506 1164 7548 1192
rect 7042 1084 7084 1112
rect 6896 252 6924 1084
rect 7056 252 7084 1084
rect 7520 252 7548 1164
rect 7680 1164 7722 1192
rect 7680 252 7708 1164
rect 8158 1112 8186 1258
rect 8144 1084 8186 1112
rect 8290 1112 8318 1258
rect 8754 1192 8782 1258
rect 8942 1192 8970 1258
rect 8754 1164 8796 1192
rect 8290 1084 8332 1112
rect 8144 252 8172 1084
rect 8304 252 8332 1084
rect 8768 252 8796 1164
rect 8928 1164 8970 1192
rect 8928 252 8956 1164
rect 9406 1112 9434 1258
rect 9392 1084 9434 1112
rect 9538 1112 9566 1258
rect 10002 1192 10030 1258
rect 10190 1192 10218 1258
rect 10002 1164 10044 1192
rect 9538 1084 9580 1112
rect 9392 252 9420 1084
rect 9552 252 9580 1084
rect 10016 252 10044 1164
rect 10176 1164 10218 1192
rect 10176 252 10204 1164
rect 10654 1112 10682 1258
rect 10640 1084 10682 1112
rect 10786 1112 10814 1258
rect 11250 1192 11278 1258
rect 11438 1192 11466 1258
rect 11250 1164 11292 1192
rect 10786 1084 10828 1112
rect 10640 252 10668 1084
rect 10800 252 10828 1084
rect 11264 252 11292 1164
rect 11424 1164 11466 1192
rect 11424 252 11452 1164
rect 11902 1112 11930 1258
rect 11888 1084 11930 1112
rect 12034 1112 12062 1258
rect 12498 1192 12526 1258
rect 12686 1192 12714 1258
rect 12498 1164 12540 1192
rect 12034 1084 12076 1112
rect 11888 252 11916 1084
rect 12048 252 12076 1084
rect 12512 252 12540 1164
rect 12672 1164 12714 1192
rect 12672 252 12700 1164
rect 13150 1112 13178 1258
rect 13136 1084 13178 1112
rect 13282 1112 13310 1258
rect 13746 1192 13774 1258
rect 13934 1192 13962 1258
rect 13746 1164 13788 1192
rect 13282 1084 13324 1112
rect 13136 252 13164 1084
rect 13296 252 13324 1084
rect 13760 252 13788 1164
rect 13920 1164 13962 1192
rect 13920 252 13948 1164
rect 14398 1112 14426 1258
rect 14384 1084 14426 1112
rect 14530 1112 14558 1258
rect 14994 1192 15022 1258
rect 15182 1192 15210 1258
rect 14994 1164 15036 1192
rect 14530 1084 14572 1112
rect 14384 252 14412 1084
rect 14544 252 14572 1084
rect 15008 252 15036 1164
rect 15168 1164 15210 1192
rect 15168 252 15196 1164
rect 15646 1112 15674 1258
rect 15632 1084 15674 1112
rect 15778 1112 15806 1258
rect 16242 1192 16270 1258
rect 16430 1192 16458 1258
rect 16242 1164 16284 1192
rect 15778 1084 15820 1112
rect 15632 252 15660 1084
rect 15792 252 15820 1084
rect 16256 252 16284 1164
rect 16416 1164 16458 1192
rect 16416 252 16444 1164
rect 16894 1112 16922 1258
rect 16880 1084 16922 1112
rect 17026 1112 17054 1258
rect 17490 1192 17518 1258
rect 17678 1192 17706 1258
rect 17490 1164 17532 1192
rect 17026 1084 17068 1112
rect 16880 252 16908 1084
rect 17040 252 17068 1084
rect 17504 252 17532 1164
rect 17664 1164 17706 1192
rect 17664 252 17692 1164
rect 18142 1112 18170 1258
rect 18128 1084 18170 1112
rect 18274 1112 18302 1258
rect 18738 1192 18766 1258
rect 18926 1192 18954 1258
rect 18738 1164 18780 1192
rect 18274 1084 18316 1112
rect 18128 252 18156 1084
rect 18288 252 18316 1084
rect 18752 252 18780 1164
rect 18912 1164 18954 1192
rect 18912 252 18940 1164
rect 19390 1112 19418 1258
rect 19376 1084 19418 1112
rect 19522 1112 19550 1258
rect 19986 1192 20014 1258
rect 20174 1192 20202 1258
rect 19986 1164 20028 1192
rect 19522 1084 19564 1112
rect 19376 252 19404 1084
rect 19536 252 19564 1084
rect 20000 252 20028 1164
rect 20160 1164 20202 1192
rect 20160 252 20188 1164
rect 20638 1112 20666 1258
rect 20624 1084 20666 1112
rect 20770 1112 20798 1258
rect 21234 1192 21262 1258
rect 21422 1192 21450 1258
rect 21234 1164 21276 1192
rect 20770 1084 20812 1112
rect 20624 252 20652 1084
rect 20784 252 20812 1084
rect 21248 252 21276 1164
rect 21408 1164 21450 1192
rect 21408 252 21436 1164
rect 21886 1112 21914 1258
rect 21872 1084 21914 1112
rect 22018 1112 22046 1258
rect 22482 1192 22510 1258
rect 22670 1192 22698 1258
rect 22482 1164 22524 1192
rect 22018 1084 22060 1112
rect 21872 252 21900 1084
rect 22032 252 22060 1084
rect 22496 252 22524 1164
rect 22656 1164 22698 1192
rect 22656 252 22684 1164
rect 23134 1112 23162 1258
rect 23120 1084 23162 1112
rect 23266 1112 23294 1258
rect 23730 1192 23758 1258
rect 23918 1192 23946 1258
rect 23730 1164 23772 1192
rect 23266 1084 23308 1112
rect 23120 252 23148 1084
rect 23280 252 23308 1084
rect 23744 252 23772 1164
rect 23904 1164 23946 1192
rect 23904 252 23932 1164
rect 24382 1112 24410 1258
rect 24368 1084 24410 1112
rect 24514 1112 24542 1258
rect 24978 1192 25006 1258
rect 25166 1192 25194 1258
rect 24978 1164 25020 1192
rect 24514 1084 24556 1112
rect 24368 252 24396 1084
rect 24528 252 24556 1084
rect 24992 252 25020 1164
rect 25152 1164 25194 1192
rect 25152 252 25180 1164
rect 25630 1112 25658 1258
rect 25616 1084 25658 1112
rect 25762 1112 25790 1258
rect 26226 1192 26254 1258
rect 26414 1192 26442 1258
rect 26226 1164 26268 1192
rect 25762 1084 25804 1112
rect 25616 252 25644 1084
rect 25776 252 25804 1084
rect 26240 252 26268 1164
rect 26400 1164 26442 1192
rect 26400 252 26428 1164
rect 26878 1112 26906 1258
rect 26864 1084 26906 1112
rect 27010 1112 27038 1258
rect 27474 1192 27502 1258
rect 27662 1192 27690 1258
rect 27474 1164 27516 1192
rect 27010 1084 27052 1112
rect 26864 252 26892 1084
rect 27024 252 27052 1084
rect 27488 252 27516 1164
rect 27648 1164 27690 1192
rect 27648 252 27676 1164
rect 28126 1112 28154 1258
rect 28112 1084 28154 1112
rect 28258 1112 28286 1258
rect 28722 1192 28750 1258
rect 28910 1192 28938 1258
rect 28722 1164 28764 1192
rect 28258 1084 28300 1112
rect 28112 252 28140 1084
rect 28272 252 28300 1084
rect 28736 252 28764 1164
rect 28896 1164 28938 1192
rect 28896 252 28924 1164
rect 29374 1112 29402 1258
rect 29360 1084 29402 1112
rect 29506 1112 29534 1258
rect 29970 1192 29998 1258
rect 30158 1192 30186 1258
rect 29970 1164 30012 1192
rect 29506 1084 29548 1112
rect 29360 252 29388 1084
rect 29520 252 29548 1084
rect 29984 252 30012 1164
rect 30144 1164 30186 1192
rect 30144 252 30172 1164
rect 30622 1112 30650 1258
rect 30608 1084 30650 1112
rect 30754 1112 30782 1258
rect 31218 1192 31246 1258
rect 31406 1192 31434 1258
rect 31218 1164 31260 1192
rect 30754 1084 30796 1112
rect 30608 252 30636 1084
rect 30768 252 30796 1084
rect 31232 252 31260 1164
rect 31392 1164 31434 1192
rect 31392 252 31420 1164
rect 31870 1112 31898 1258
rect 31856 1084 31898 1112
rect 32002 1112 32030 1258
rect 32466 1192 32494 1258
rect 32654 1192 32682 1258
rect 32466 1164 32508 1192
rect 32002 1084 32044 1112
rect 31856 252 31884 1084
rect 32016 252 32044 1084
rect 32480 252 32508 1164
rect 32640 1164 32682 1192
rect 32640 252 32668 1164
rect 33118 1112 33146 1258
rect 33104 1084 33146 1112
rect 33250 1112 33278 1258
rect 33714 1192 33742 1258
rect 33902 1192 33930 1258
rect 33714 1164 33756 1192
rect 33250 1084 33292 1112
rect 33104 252 33132 1084
rect 33264 252 33292 1084
rect 33728 252 33756 1164
rect 33888 1164 33930 1192
rect 33888 252 33916 1164
rect 34366 1112 34394 1258
rect 34352 1084 34394 1112
rect 34498 1112 34526 1258
rect 34962 1192 34990 1258
rect 35150 1192 35178 1258
rect 34962 1164 35004 1192
rect 34498 1084 34540 1112
rect 34352 252 34380 1084
rect 34512 252 34540 1084
rect 34976 252 35004 1164
rect 35136 1164 35178 1192
rect 35136 252 35164 1164
rect 35614 1112 35642 1258
rect 35600 1084 35642 1112
rect 35746 1112 35774 1258
rect 36210 1192 36238 1258
rect 36398 1192 36426 1258
rect 36210 1164 36252 1192
rect 35746 1084 35788 1112
rect 35600 252 35628 1084
rect 35760 252 35788 1084
rect 36224 252 36252 1164
rect 36384 1164 36426 1192
rect 36384 252 36412 1164
rect 36862 1112 36890 1258
rect 36848 1084 36890 1112
rect 36994 1112 37022 1258
rect 37458 1192 37486 1258
rect 37646 1192 37674 1258
rect 37458 1164 37500 1192
rect 36994 1084 37036 1112
rect 36848 252 36876 1084
rect 37008 252 37036 1084
rect 37472 252 37500 1164
rect 37632 1164 37674 1192
rect 37632 252 37660 1164
rect 38110 1112 38138 1258
rect 38096 1084 38138 1112
rect 38242 1112 38270 1258
rect 38706 1192 38734 1258
rect 38894 1192 38922 1258
rect 38706 1164 38748 1192
rect 38242 1084 38284 1112
rect 38096 252 38124 1084
rect 38256 252 38284 1084
rect 38720 252 38748 1164
rect 38880 1164 38922 1192
rect 38880 252 38908 1164
rect 39358 1112 39386 1258
rect 39344 1084 39386 1112
rect 39490 1112 39518 1258
rect 39954 1192 39982 1258
rect 40142 1192 40170 1258
rect 39954 1164 39996 1192
rect 39490 1084 39532 1112
rect 39344 252 39372 1084
rect 39504 252 39532 1084
rect 39968 252 39996 1164
rect 40128 1164 40170 1192
rect 40128 252 40156 1164
rect 40606 1112 40634 1258
rect 40592 1084 40634 1112
rect 40738 1112 40766 1258
rect 41202 1192 41230 1258
rect 41202 1164 41244 1192
rect 40738 1084 40780 1112
rect 40592 252 40620 1084
rect 40752 252 40780 1084
rect 41216 252 41244 1164
<< via1 >>
rect 10723 8777 10775 8829
rect 20707 8777 20759 8829
rect 30691 8777 30743 8829
rect 40675 8777 40727 8829
rect 10723 7828 10775 7880
rect 20707 7828 20759 7880
rect 30691 7828 30743 7880
rect 40675 7828 40727 7880
<< metal2 >>
rect 1360 9053 1388 9081
rect 11344 9053 11372 9081
rect 21328 9053 21356 9081
rect 31312 9053 31340 9081
rect 10723 8829 10775 8835
rect 10723 8771 10775 8777
rect 20707 8829 20759 8835
rect 20707 8771 20759 8777
rect 30691 8829 30743 8835
rect 30691 8771 30743 8777
rect 40675 8829 40727 8835
rect 40675 8771 40727 8777
rect 10735 7886 10763 8771
rect 20719 7886 20747 8771
rect 30703 7886 30731 8771
rect 40687 7886 40715 8771
rect 10723 7880 10775 7886
rect 10723 7822 10775 7828
rect 20707 7880 20759 7886
rect 20707 7822 20759 7828
rect 30691 7880 30743 7886
rect 30691 7822 30743 7828
rect 40675 7880 40727 7886
rect 40675 7822 40727 7828
<< metal3 >>
rect -49 9288 49 9386
rect 41261 9288 41359 9386
rect 0 8789 41310 8849
rect -49 8168 49 8266
rect 41261 8168 41359 8266
rect 1601 7725 1699 7823
rect 2849 7725 2947 7823
rect 4097 7725 4195 7823
rect 5345 7725 5443 7823
rect 6593 7725 6691 7823
rect 7841 7725 7939 7823
rect 9089 7725 9187 7823
rect 10337 7725 10435 7823
rect 11585 7725 11683 7823
rect 12833 7725 12931 7823
rect 14081 7725 14179 7823
rect 15329 7725 15427 7823
rect 16577 7725 16675 7823
rect 17825 7725 17923 7823
rect 19073 7725 19171 7823
rect 20321 7725 20419 7823
rect 21569 7725 21667 7823
rect 22817 7725 22915 7823
rect 24065 7725 24163 7823
rect 25313 7725 25411 7823
rect 26561 7725 26659 7823
rect 27809 7725 27907 7823
rect 29057 7725 29155 7823
rect 30305 7725 30403 7823
rect 31553 7725 31651 7823
rect 32801 7725 32899 7823
rect 34049 7725 34147 7823
rect 35297 7725 35395 7823
rect 36545 7725 36643 7823
rect 37793 7725 37891 7823
rect 39041 7725 39139 7823
rect 40289 7725 40387 7823
rect 1587 7309 1685 7407
rect 2835 7309 2933 7407
rect 4083 7309 4181 7407
rect 5331 7309 5429 7407
rect 6579 7309 6677 7407
rect 7827 7309 7925 7407
rect 9075 7309 9173 7407
rect 10323 7309 10421 7407
rect 11571 7309 11669 7407
rect 12819 7309 12917 7407
rect 14067 7309 14165 7407
rect 15315 7309 15413 7407
rect 16563 7309 16661 7407
rect 17811 7309 17909 7407
rect 19059 7309 19157 7407
rect 20307 7309 20405 7407
rect 21555 7309 21653 7407
rect 22803 7309 22901 7407
rect 24051 7309 24149 7407
rect 25299 7309 25397 7407
rect 26547 7309 26645 7407
rect 27795 7309 27893 7407
rect 29043 7309 29141 7407
rect 30291 7309 30389 7407
rect 31539 7309 31637 7407
rect 32787 7309 32885 7407
rect 34035 7309 34133 7407
rect 35283 7309 35381 7407
rect 36531 7309 36629 7407
rect 37779 7309 37877 7407
rect 39027 7309 39125 7407
rect 40275 7309 40373 7407
rect 1702 7107 1800 7205
rect 2950 7107 3048 7205
rect 4198 7107 4296 7205
rect 5446 7107 5544 7205
rect 6694 7107 6792 7205
rect 7942 7107 8040 7205
rect 9190 7107 9288 7205
rect 10438 7107 10536 7205
rect 11686 7107 11784 7205
rect 12934 7107 13032 7205
rect 14182 7107 14280 7205
rect 15430 7107 15528 7205
rect 16678 7107 16776 7205
rect 17926 7107 18024 7205
rect 19174 7107 19272 7205
rect 20422 7107 20520 7205
rect 21670 7107 21768 7205
rect 22918 7107 23016 7205
rect 24166 7107 24264 7205
rect 25414 7107 25512 7205
rect 26662 7107 26760 7205
rect 27910 7107 28008 7205
rect 29158 7107 29256 7205
rect 30406 7107 30504 7205
rect 31654 7107 31752 7205
rect 32902 7107 33000 7205
rect 34150 7107 34248 7205
rect 35398 7107 35496 7205
rect 36646 7107 36744 7205
rect 37894 7107 37992 7205
rect 39142 7107 39240 7205
rect 40390 7107 40488 7205
rect 1581 6775 1679 6873
rect 2829 6775 2927 6873
rect 4077 6775 4175 6873
rect 5325 6775 5423 6873
rect 6573 6775 6671 6873
rect 7821 6775 7919 6873
rect 9069 6775 9167 6873
rect 10317 6775 10415 6873
rect 11565 6775 11663 6873
rect 12813 6775 12911 6873
rect 14061 6775 14159 6873
rect 15309 6775 15407 6873
rect 16557 6775 16655 6873
rect 17805 6775 17903 6873
rect 19053 6775 19151 6873
rect 20301 6775 20399 6873
rect 21549 6775 21647 6873
rect 22797 6775 22895 6873
rect 24045 6775 24143 6873
rect 25293 6775 25391 6873
rect 26541 6775 26639 6873
rect 27789 6775 27887 6873
rect 29037 6775 29135 6873
rect 30285 6775 30383 6873
rect 31533 6775 31631 6873
rect 32781 6775 32879 6873
rect 34029 6775 34127 6873
rect 35277 6775 35375 6873
rect 36525 6775 36623 6873
rect 37773 6775 37871 6873
rect 39021 6775 39119 6873
rect 40269 6775 40367 6873
rect 1592 6338 1690 6436
rect 2840 6338 2938 6436
rect 4088 6338 4186 6436
rect 5336 6338 5434 6436
rect 6584 6338 6682 6436
rect 7832 6338 7930 6436
rect 9080 6338 9178 6436
rect 10328 6338 10426 6436
rect 11576 6338 11674 6436
rect 12824 6338 12922 6436
rect 14072 6338 14170 6436
rect 15320 6338 15418 6436
rect 16568 6338 16666 6436
rect 17816 6338 17914 6436
rect 19064 6338 19162 6436
rect 20312 6338 20410 6436
rect 21560 6338 21658 6436
rect 22808 6338 22906 6436
rect 24056 6338 24154 6436
rect 25304 6338 25402 6436
rect 26552 6338 26650 6436
rect 27800 6338 27898 6436
rect 29048 6338 29146 6436
rect 30296 6338 30394 6436
rect 31544 6338 31642 6436
rect 32792 6338 32890 6436
rect 34040 6338 34138 6436
rect 35288 6338 35386 6436
rect 36536 6338 36634 6436
rect 37784 6338 37882 6436
rect 39032 6338 39130 6436
rect 40280 6338 40378 6436
rect 1706 5545 1804 5643
rect 2954 5545 3052 5643
rect 4202 5545 4300 5643
rect 5450 5545 5548 5643
rect 6698 5545 6796 5643
rect 7946 5545 8044 5643
rect 9194 5545 9292 5643
rect 10442 5545 10540 5643
rect 11690 5545 11788 5643
rect 12938 5545 13036 5643
rect 14186 5545 14284 5643
rect 15434 5545 15532 5643
rect 16682 5545 16780 5643
rect 17930 5545 18028 5643
rect 19178 5545 19276 5643
rect 20426 5545 20524 5643
rect 21674 5545 21772 5643
rect 22922 5545 23020 5643
rect 24170 5545 24268 5643
rect 25418 5545 25516 5643
rect 26666 5545 26764 5643
rect 27914 5545 28012 5643
rect 29162 5545 29260 5643
rect 30410 5545 30508 5643
rect 31658 5545 31756 5643
rect 32906 5545 33004 5643
rect 34154 5545 34252 5643
rect 35402 5545 35500 5643
rect 36650 5545 36748 5643
rect 37898 5545 37996 5643
rect 39146 5545 39244 5643
rect 40394 5545 40492 5643
rect 1706 5223 1804 5321
rect 2954 5223 3052 5321
rect 4202 5223 4300 5321
rect 5450 5223 5548 5321
rect 6698 5223 6796 5321
rect 7946 5223 8044 5321
rect 9194 5223 9292 5321
rect 10442 5223 10540 5321
rect 11690 5223 11788 5321
rect 12938 5223 13036 5321
rect 14186 5223 14284 5321
rect 15434 5223 15532 5321
rect 16682 5223 16780 5321
rect 17930 5223 18028 5321
rect 19178 5223 19276 5321
rect 20426 5223 20524 5321
rect 21674 5223 21772 5321
rect 22922 5223 23020 5321
rect 24170 5223 24268 5321
rect 25418 5223 25516 5321
rect 26666 5223 26764 5321
rect 27914 5223 28012 5321
rect 29162 5223 29260 5321
rect 30410 5223 30508 5321
rect 31658 5223 31756 5321
rect 32906 5223 33004 5321
rect 34154 5223 34252 5321
rect 35402 5223 35500 5321
rect 36650 5223 36748 5321
rect 37898 5223 37996 5321
rect 39146 5223 39244 5321
rect 40394 5223 40492 5321
rect 1694 4385 1792 4483
rect 2942 4385 3040 4483
rect 4190 4385 4288 4483
rect 5438 4385 5536 4483
rect 6686 4385 6784 4483
rect 7934 4385 8032 4483
rect 9182 4385 9280 4483
rect 10430 4385 10528 4483
rect 11678 4385 11776 4483
rect 12926 4385 13024 4483
rect 14174 4385 14272 4483
rect 15422 4385 15520 4483
rect 16670 4385 16768 4483
rect 17918 4385 18016 4483
rect 19166 4385 19264 4483
rect 20414 4385 20512 4483
rect 21662 4385 21760 4483
rect 22910 4385 23008 4483
rect 24158 4385 24256 4483
rect 25406 4385 25504 4483
rect 26654 4385 26752 4483
rect 27902 4385 28000 4483
rect 29150 4385 29248 4483
rect 30398 4385 30496 4483
rect 31646 4385 31744 4483
rect 32894 4385 32992 4483
rect 34142 4385 34240 4483
rect 35390 4385 35488 4483
rect 36638 4385 36736 4483
rect 37886 4385 37984 4483
rect 39134 4385 39232 4483
rect 40382 4385 40480 4483
rect 1776 3611 1874 3709
rect 3024 3611 3122 3709
rect 4272 3611 4370 3709
rect 5520 3611 5618 3709
rect 6768 3611 6866 3709
rect 8016 3611 8114 3709
rect 9264 3611 9362 3709
rect 10512 3611 10610 3709
rect 11760 3611 11858 3709
rect 13008 3611 13106 3709
rect 14256 3611 14354 3709
rect 15504 3611 15602 3709
rect 16752 3611 16850 3709
rect 18000 3611 18098 3709
rect 19248 3611 19346 3709
rect 20496 3611 20594 3709
rect 21744 3611 21842 3709
rect 22992 3611 23090 3709
rect 24240 3611 24338 3709
rect 25488 3611 25586 3709
rect 26736 3611 26834 3709
rect 27984 3611 28082 3709
rect 29232 3611 29330 3709
rect 30480 3611 30578 3709
rect 31728 3611 31826 3709
rect 32976 3611 33074 3709
rect 34224 3611 34322 3709
rect 35472 3611 35570 3709
rect 36720 3611 36818 3709
rect 37968 3611 38066 3709
rect 39216 3611 39314 3709
rect 40464 3611 40562 3709
rect 0 3478 40562 3538
rect 0 2762 41310 2822
rect 0 2638 41310 2698
rect 1949 1862 2047 1960
rect 3197 1862 3295 1960
rect 4445 1862 4543 1960
rect 5693 1862 5791 1960
rect 6941 1862 7039 1960
rect 8189 1862 8287 1960
rect 9437 1862 9535 1960
rect 10685 1862 10783 1960
rect 11933 1862 12031 1960
rect 13181 1862 13279 1960
rect 14429 1862 14527 1960
rect 15677 1862 15775 1960
rect 16925 1862 17023 1960
rect 18173 1862 18271 1960
rect 19421 1862 19519 1960
rect 20669 1862 20767 1960
rect 21917 1862 22015 1960
rect 23165 1862 23263 1960
rect 24413 1862 24511 1960
rect 25661 1862 25759 1960
rect 26909 1862 27007 1960
rect 28157 1862 28255 1960
rect 29405 1862 29503 1960
rect 30653 1862 30751 1960
rect 31901 1862 31999 1960
rect 33149 1862 33247 1960
rect 34397 1862 34495 1960
rect 35645 1862 35743 1960
rect 36893 1862 36991 1960
rect 38141 1862 38239 1960
rect 39389 1862 39487 1960
rect 40637 1862 40735 1960
rect 0 951 41310 1011
rect 1132 313 1230 411
rect 1518 313 1616 411
rect 2380 313 2478 411
rect 2766 313 2864 411
rect 3628 313 3726 411
rect 4014 313 4112 411
rect 4876 313 4974 411
rect 5262 313 5360 411
rect 6124 313 6222 411
rect 6510 313 6608 411
rect 7372 313 7470 411
rect 7758 313 7856 411
rect 8620 313 8718 411
rect 9006 313 9104 411
rect 9868 313 9966 411
rect 10254 313 10352 411
rect 11116 313 11214 411
rect 11502 313 11600 411
rect 12364 313 12462 411
rect 12750 313 12848 411
rect 13612 313 13710 411
rect 13998 313 14096 411
rect 14860 313 14958 411
rect 15246 313 15344 411
rect 16108 313 16206 411
rect 16494 313 16592 411
rect 17356 313 17454 411
rect 17742 313 17840 411
rect 18604 313 18702 411
rect 18990 313 19088 411
rect 19852 313 19950 411
rect 20238 313 20336 411
rect 21100 313 21198 411
rect 21486 313 21584 411
rect 22348 313 22446 411
rect 22734 313 22832 411
rect 23596 313 23694 411
rect 23982 313 24080 411
rect 24844 313 24942 411
rect 25230 313 25328 411
rect 26092 313 26190 411
rect 26478 313 26576 411
rect 27340 313 27438 411
rect 27726 313 27824 411
rect 28588 313 28686 411
rect 28974 313 29072 411
rect 29836 313 29934 411
rect 30222 313 30320 411
rect 31084 313 31182 411
rect 31470 313 31568 411
rect 32332 313 32430 411
rect 32718 313 32816 411
rect 33580 313 33678 411
rect 33966 313 34064 411
rect 34828 313 34926 411
rect 35214 313 35312 411
rect 36076 313 36174 411
rect 36462 313 36560 411
rect 37324 313 37422 411
rect 37710 313 37808 411
rect 38572 313 38670 411
rect 38958 313 39056 411
rect 39820 313 39918 411
rect 40206 313 40304 411
rect 41068 313 41166 411
use sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_array  sky130_sram_1kbyte_1rw1r_32x256_8_column_mux_array_0
timestamp 1666199351
transform 1 0 0 0 -1 3194
box 0 87 41310 1936
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_0
timestamp 1666199351
transform 1 0 31875 0 1 8770
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_1
timestamp 1666199351
transform 1 0 21891 0 1 8770
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_2
timestamp 1666199351
transform 1 0 11907 0 1 8770
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_3
timestamp 1666199351
transform 1 0 1923 0 1 8770
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_0
timestamp 1666199351
transform 1 0 40669 0 1 8771
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_1
timestamp 1666199351
transform 1 0 40669 0 1 7822
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_2
timestamp 1666199351
transform 1 0 30685 0 1 8771
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_3
timestamp 1666199351
transform 1 0 30685 0 1 7822
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_4
timestamp 1666199351
transform 1 0 20701 0 1 8771
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_5
timestamp 1666199351
transform 1 0 20701 0 1 7822
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_6
timestamp 1666199351
transform 1 0 10717 0 1 8771
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_7
timestamp 1666199351
transform 1 0 10717 0 1 7822
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_precharge_array  sky130_sram_1kbyte_1rw1r_32x256_8_precharge_array_0
timestamp 1666199351
transform 1 0 0 0 -1 1006
box 0 -12 41310 768
use sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array  sky130_sram_1kbyte_1rw1r_32x256_8_sense_amp_array_0
timestamp 1666199351
transform 1 0 0 0 -1 5702
box 0 0 40999 2256
use sky130_sram_1kbyte_1rw1r_32x256_8_write_driver_array  sky130_sram_1kbyte_1rw1r_32x256_8_write_driver_array_0
timestamp 1666199351
transform 1 0 0 0 -1 7965
box 998 4 40942 2011
use sky130_sram_1kbyte_1rw1r_32x256_8_write_mask_and_array  sky130_sram_1kbyte_1rw1r_32x256_8_write_mask_and_array_0
timestamp 1666199351
transform 1 0 0 0 -1 9337
box -49 -49 41359 1177
<< labels >>
rlabel metal3 s 40394 5223 40492 5321 4 vdd
port 1 nsew
rlabel metal3 s 37773 6775 37871 6873 4 vdd
port 1 nsew
rlabel metal3 s 32781 6775 32879 6873 4 vdd
port 1 nsew
rlabel metal3 s 37793 7725 37891 7823 4 vdd
port 1 nsew
rlabel metal3 s 37898 5223 37996 5321 4 vdd
port 1 nsew
rlabel metal3 s 40289 7725 40387 7823 4 vdd
port 1 nsew
rlabel metal3 s 32801 7725 32899 7823 4 vdd
port 1 nsew
rlabel metal3 s 32906 5223 33004 5321 4 vdd
port 1 nsew
rlabel metal3 s 31553 7725 31651 7823 4 vdd
port 1 nsew
rlabel metal3 s 36525 6775 36623 6873 4 vdd
port 1 nsew
rlabel metal3 s 39146 5223 39244 5321 4 vdd
port 1 nsew
rlabel metal3 s 36545 7725 36643 7823 4 vdd
port 1 nsew
rlabel metal3 s 35277 6775 35375 6873 4 vdd
port 1 nsew
rlabel metal3 s 36650 5223 36748 5321 4 vdd
port 1 nsew
rlabel metal3 s 31533 6775 31631 6873 4 vdd
port 1 nsew
rlabel metal3 s 39021 6775 39119 6873 4 vdd
port 1 nsew
rlabel metal3 s 31658 5223 31756 5321 4 vdd
port 1 nsew
rlabel metal3 s 39041 7725 39139 7823 4 vdd
port 1 nsew
rlabel metal3 s 41261 8168 41359 8266 4 vdd
port 1 nsew
rlabel metal3 s 34049 7725 34147 7823 4 vdd
port 1 nsew
rlabel metal3 s 40269 6775 40367 6873 4 vdd
port 1 nsew
rlabel metal3 s 35297 7725 35395 7823 4 vdd
port 1 nsew
rlabel metal3 s 34029 6775 34127 6873 4 vdd
port 1 nsew
rlabel metal3 s 34154 5223 34252 5321 4 vdd
port 1 nsew
rlabel metal3 s 35402 5223 35500 5321 4 vdd
port 1 nsew
rlabel metal3 s 39146 5545 39244 5643 4 gnd
port 2 nsew
rlabel metal3 s 36646 7107 36744 7205 4 gnd
port 2 nsew
rlabel metal3 s 37894 7107 37992 7205 4 gnd
port 2 nsew
rlabel metal3 s 31539 7309 31637 7407 4 gnd
port 2 nsew
rlabel metal3 s 40390 7107 40488 7205 4 gnd
port 2 nsew
rlabel metal3 s 39027 7309 39125 7407 4 gnd
port 2 nsew
rlabel metal3 s 35402 5545 35500 5643 4 gnd
port 2 nsew
rlabel metal3 s 40280 6338 40378 6436 4 gnd
port 2 nsew
rlabel metal3 s 31544 6338 31642 6436 4 gnd
port 2 nsew
rlabel metal3 s 37779 7309 37877 7407 4 gnd
port 2 nsew
rlabel metal3 s 32792 6338 32890 6436 4 gnd
port 2 nsew
rlabel metal3 s 34040 6338 34138 6436 4 gnd
port 2 nsew
rlabel metal3 s 34150 7107 34248 7205 4 gnd
port 2 nsew
rlabel metal3 s 36650 5545 36748 5643 4 gnd
port 2 nsew
rlabel metal3 s 41261 9288 41359 9386 4 gnd
port 2 nsew
rlabel metal3 s 35283 7309 35381 7407 4 gnd
port 2 nsew
rlabel metal3 s 32902 7107 33000 7205 4 gnd
port 2 nsew
rlabel metal3 s 34154 5545 34252 5643 4 gnd
port 2 nsew
rlabel metal3 s 34035 7309 34133 7407 4 gnd
port 2 nsew
rlabel metal3 s 36536 6338 36634 6436 4 gnd
port 2 nsew
rlabel metal3 s 32787 7309 32885 7407 4 gnd
port 2 nsew
rlabel metal3 s 31654 7107 31752 7205 4 gnd
port 2 nsew
rlabel metal3 s 39032 6338 39130 6436 4 gnd
port 2 nsew
rlabel metal3 s 37898 5545 37996 5643 4 gnd
port 2 nsew
rlabel metal3 s 36531 7309 36629 7407 4 gnd
port 2 nsew
rlabel metal3 s 31658 5545 31756 5643 4 gnd
port 2 nsew
rlabel metal3 s 32906 5545 33004 5643 4 gnd
port 2 nsew
rlabel metal3 s 37784 6338 37882 6436 4 gnd
port 2 nsew
rlabel metal3 s 39142 7107 39240 7205 4 gnd
port 2 nsew
rlabel metal3 s 35398 7107 35496 7205 4 gnd
port 2 nsew
rlabel metal3 s 40275 7309 40373 7407 4 gnd
port 2 nsew
rlabel metal3 s 35288 6338 35386 6436 4 gnd
port 2 nsew
rlabel metal3 s 40394 5545 40492 5643 4 gnd
port 2 nsew
rlabel metal3 s 25313 7725 25411 7823 4 vdd
port 1 nsew
rlabel metal3 s 29158 7107 29256 7205 4 gnd
port 2 nsew
rlabel metal3 s 26561 7725 26659 7823 4 vdd
port 1 nsew
rlabel metal3 s 27789 6775 27887 6873 4 vdd
port 1 nsew
rlabel metal3 s 22817 7725 22915 7823 4 vdd
port 1 nsew
rlabel metal3 s 25293 6775 25391 6873 4 vdd
port 1 nsew
rlabel metal3 s 22922 5545 23020 5643 4 gnd
port 2 nsew
rlabel metal3 s 25299 7309 25397 7407 4 gnd
port 2 nsew
rlabel metal3 s 29162 5545 29260 5643 4 gnd
port 2 nsew
rlabel metal3 s 26666 5223 26764 5321 4 vdd
port 1 nsew
rlabel metal3 s 21549 6775 21647 6873 4 vdd
port 1 nsew
rlabel metal3 s 29037 6775 29135 6873 4 vdd
port 1 nsew
rlabel metal3 s 29162 5223 29260 5321 4 vdd
port 1 nsew
rlabel metal3 s 22918 7107 23016 7205 4 gnd
port 2 nsew
rlabel metal3 s 27800 6338 27898 6436 4 gnd
port 2 nsew
rlabel metal3 s 30305 7725 30403 7823 4 vdd
port 1 nsew
rlabel metal3 s 30291 7309 30389 7407 4 gnd
port 2 nsew
rlabel metal3 s 24170 5545 24268 5643 4 gnd
port 2 nsew
rlabel metal3 s 30296 6338 30394 6436 4 gnd
port 2 nsew
rlabel metal3 s 27809 7725 27907 7823 4 vdd
port 1 nsew
rlabel metal3 s 21555 7309 21653 7407 4 gnd
port 2 nsew
rlabel metal3 s 27914 5545 28012 5643 4 gnd
port 2 nsew
rlabel metal3 s 24065 7725 24163 7823 4 vdd
port 1 nsew
rlabel metal3 s 24170 5223 24268 5321 4 vdd
port 1 nsew
rlabel metal3 s 21674 5545 21772 5643 4 gnd
port 2 nsew
rlabel metal3 s 25418 5545 25516 5643 4 gnd
port 2 nsew
rlabel metal3 s 29057 7725 29155 7823 4 vdd
port 1 nsew
rlabel metal3 s 30410 5223 30508 5321 4 vdd
port 1 nsew
rlabel metal3 s 22922 5223 23020 5321 4 vdd
port 1 nsew
rlabel metal3 s 21560 6338 21658 6436 4 gnd
port 2 nsew
rlabel metal3 s 27914 5223 28012 5321 4 vdd
port 1 nsew
rlabel metal3 s 26666 5545 26764 5643 4 gnd
port 2 nsew
rlabel metal3 s 27910 7107 28008 7205 4 gnd
port 2 nsew
rlabel metal3 s 22797 6775 22895 6873 4 vdd
port 1 nsew
rlabel metal3 s 26541 6775 26639 6873 4 vdd
port 1 nsew
rlabel metal3 s 22803 7309 22901 7407 4 gnd
port 2 nsew
rlabel metal3 s 24045 6775 24143 6873 4 vdd
port 1 nsew
rlabel metal3 s 24056 6338 24154 6436 4 gnd
port 2 nsew
rlabel metal3 s 24051 7309 24149 7407 4 gnd
port 2 nsew
rlabel metal3 s 22808 6338 22906 6436 4 gnd
port 2 nsew
rlabel metal3 s 26662 7107 26760 7205 4 gnd
port 2 nsew
rlabel metal3 s 26552 6338 26650 6436 4 gnd
port 2 nsew
rlabel metal3 s 25414 7107 25512 7205 4 gnd
port 2 nsew
rlabel metal3 s 21670 7107 21768 7205 4 gnd
port 2 nsew
rlabel metal3 s 30410 5545 30508 5643 4 gnd
port 2 nsew
rlabel metal3 s 25304 6338 25402 6436 4 gnd
port 2 nsew
rlabel metal3 s 26547 7309 26645 7407 4 gnd
port 2 nsew
rlabel metal3 s 24166 7107 24264 7205 4 gnd
port 2 nsew
rlabel metal3 s 21674 5223 21772 5321 4 vdd
port 1 nsew
rlabel metal3 s 29043 7309 29141 7407 4 gnd
port 2 nsew
rlabel metal3 s 25418 5223 25516 5321 4 vdd
port 1 nsew
rlabel metal3 s 27795 7309 27893 7407 4 gnd
port 2 nsew
rlabel metal3 s 29048 6338 29146 6436 4 gnd
port 2 nsew
rlabel metal3 s 30285 6775 30383 6873 4 vdd
port 1 nsew
rlabel metal3 s 21569 7725 21667 7823 4 vdd
port 1 nsew
rlabel metal3 s 30406 7107 30504 7205 4 gnd
port 2 nsew
rlabel metal3 s 26909 1862 27007 1960 4 gnd
port 2 nsew
rlabel metal3 s 24158 4385 24256 4483 4 vdd
port 1 nsew
rlabel metal3 s 29405 1862 29503 1960 4 gnd
port 2 nsew
rlabel metal3 s 22910 4385 23008 4483 4 vdd
port 1 nsew
rlabel metal3 s 26736 3611 26834 3709 4 gnd
port 2 nsew
rlabel metal3 s 25406 4385 25504 4483 4 vdd
port 1 nsew
rlabel metal3 s 21917 1862 22015 1960 4 gnd
port 2 nsew
rlabel metal3 s 29232 3611 29330 3709 4 gnd
port 2 nsew
rlabel metal3 s 21744 3611 21842 3709 4 gnd
port 2 nsew
rlabel metal3 s 26654 4385 26752 4483 4 vdd
port 1 nsew
rlabel metal3 s 30653 1862 30751 1960 4 gnd
port 2 nsew
rlabel metal3 s 28157 1862 28255 1960 4 gnd
port 2 nsew
rlabel metal3 s 30480 3611 30578 3709 4 gnd
port 2 nsew
rlabel metal3 s 27984 3611 28082 3709 4 gnd
port 2 nsew
rlabel metal3 s 24413 1862 24511 1960 4 gnd
port 2 nsew
rlabel metal3 s 21662 4385 21760 4483 4 vdd
port 1 nsew
rlabel metal3 s 24240 3611 24338 3709 4 gnd
port 2 nsew
rlabel metal3 s 30398 4385 30496 4483 4 vdd
port 1 nsew
rlabel metal3 s 25661 1862 25759 1960 4 gnd
port 2 nsew
rlabel metal3 s 20669 1862 20767 1960 4 gnd
port 2 nsew
rlabel metal3 s 27902 4385 28000 4483 4 vdd
port 1 nsew
rlabel metal3 s 23165 1862 23263 1960 4 gnd
port 2 nsew
rlabel metal3 s 22992 3611 23090 3709 4 gnd
port 2 nsew
rlabel metal3 s 29150 4385 29248 4483 4 vdd
port 1 nsew
rlabel metal3 s 25488 3611 25586 3709 4 gnd
port 2 nsew
rlabel metal3 s 40637 1862 40735 1960 4 gnd
port 2 nsew
rlabel metal3 s 31728 3611 31826 3709 4 gnd
port 2 nsew
rlabel metal3 s 40382 4385 40480 4483 4 vdd
port 1 nsew
rlabel metal3 s 39134 4385 39232 4483 4 vdd
port 1 nsew
rlabel metal3 s 31646 4385 31744 4483 4 vdd
port 1 nsew
rlabel metal3 s 36893 1862 36991 1960 4 gnd
port 2 nsew
rlabel metal3 s 33149 1862 33247 1960 4 gnd
port 2 nsew
rlabel metal3 s 39389 1862 39487 1960 4 gnd
port 2 nsew
rlabel metal3 s 37968 3611 38066 3709 4 gnd
port 2 nsew
rlabel metal3 s 40464 3611 40562 3709 4 gnd
port 2 nsew
rlabel metal3 s 38141 1862 38239 1960 4 gnd
port 2 nsew
rlabel metal3 s 39216 3611 39314 3709 4 gnd
port 2 nsew
rlabel metal3 s 35390 4385 35488 4483 4 vdd
port 1 nsew
rlabel metal3 s 36720 3611 36818 3709 4 gnd
port 2 nsew
rlabel metal3 s 34142 4385 34240 4483 4 vdd
port 1 nsew
rlabel metal3 s 36638 4385 36736 4483 4 vdd
port 1 nsew
rlabel metal3 s 34224 3611 34322 3709 4 gnd
port 2 nsew
rlabel metal3 s 35645 1862 35743 1960 4 gnd
port 2 nsew
rlabel metal3 s 35472 3611 35570 3709 4 gnd
port 2 nsew
rlabel metal3 s 31901 1862 31999 1960 4 gnd
port 2 nsew
rlabel metal3 s 32894 4385 32992 4483 4 vdd
port 1 nsew
rlabel metal3 s 37886 4385 37984 4483 4 vdd
port 1 nsew
rlabel metal3 s 34397 1862 34495 1960 4 gnd
port 2 nsew
rlabel metal3 s 32976 3611 33074 3709 4 gnd
port 2 nsew
rlabel metal3 s 16678 7107 16776 7205 4 gnd
port 2 nsew
rlabel metal3 s 14186 5545 14284 5643 4 gnd
port 2 nsew
rlabel metal3 s 17825 7725 17923 7823 4 vdd
port 1 nsew
rlabel metal3 s 12824 6338 12922 6436 4 gnd
port 2 nsew
rlabel metal3 s 14081 7725 14179 7823 4 vdd
port 1 nsew
rlabel metal3 s 19174 7107 19272 7205 4 gnd
port 2 nsew
rlabel metal3 s 19064 6338 19162 6436 4 gnd
port 2 nsew
rlabel metal3 s 17805 6775 17903 6873 4 vdd
port 1 nsew
rlabel metal3 s 20301 6775 20399 6873 4 vdd
port 1 nsew
rlabel metal3 s 10337 7725 10435 7823 4 vdd
port 1 nsew
rlabel metal3 s 10442 5223 10540 5321 4 vdd
port 1 nsew
rlabel metal3 s 12833 7725 12931 7823 4 vdd
port 1 nsew
rlabel metal3 s 10438 7107 10536 7205 4 gnd
port 2 nsew
rlabel metal3 s 17811 7309 17909 7407 4 gnd
port 2 nsew
rlabel metal3 s 15329 7725 15427 7823 4 vdd
port 1 nsew
rlabel metal3 s 11576 6338 11674 6436 4 gnd
port 2 nsew
rlabel metal3 s 15309 6775 15407 6873 4 vdd
port 1 nsew
rlabel metal3 s 20422 7107 20520 7205 4 gnd
port 2 nsew
rlabel metal3 s 16563 7309 16661 7407 4 gnd
port 2 nsew
rlabel metal3 s 19178 5223 19276 5321 4 vdd
port 1 nsew
rlabel metal3 s 17930 5223 18028 5321 4 vdd
port 1 nsew
rlabel metal3 s 11690 5545 11788 5643 4 gnd
port 2 nsew
rlabel metal3 s 16682 5223 16780 5321 4 vdd
port 1 nsew
rlabel metal3 s 12938 5223 13036 5321 4 vdd
port 1 nsew
rlabel metal3 s 16577 7725 16675 7823 4 vdd
port 1 nsew
rlabel metal3 s 12813 6775 12911 6873 4 vdd
port 1 nsew
rlabel metal3 s 12934 7107 13032 7205 4 gnd
port 2 nsew
rlabel metal3 s 11585 7725 11683 7823 4 vdd
port 1 nsew
rlabel metal3 s 10328 6338 10426 6436 4 gnd
port 2 nsew
rlabel metal3 s 14067 7309 14165 7407 4 gnd
port 2 nsew
rlabel metal3 s 16568 6338 16666 6436 4 gnd
port 2 nsew
rlabel metal3 s 19053 6775 19151 6873 4 vdd
port 1 nsew
rlabel metal3 s 17816 6338 17914 6436 4 gnd
port 2 nsew
rlabel metal3 s 0 8789 41310 8849 4 w_en
port 3 nsew
rlabel metal3 s 20312 6338 20410 6436 4 gnd
port 2 nsew
rlabel metal3 s 20426 5223 20524 5321 4 vdd
port 1 nsew
rlabel metal3 s 11686 7107 11784 7205 4 gnd
port 2 nsew
rlabel metal3 s 10442 5545 10540 5643 4 gnd
port 2 nsew
rlabel metal3 s 10323 7309 10421 7407 4 gnd
port 2 nsew
rlabel metal3 s 12938 5545 13036 5643 4 gnd
port 2 nsew
rlabel metal3 s 11571 7309 11669 7407 4 gnd
port 2 nsew
rlabel metal3 s 15434 5223 15532 5321 4 vdd
port 1 nsew
rlabel metal3 s 14186 5223 14284 5321 4 vdd
port 1 nsew
rlabel metal3 s 19059 7309 19157 7407 4 gnd
port 2 nsew
rlabel metal3 s 17926 7107 18024 7205 4 gnd
port 2 nsew
rlabel metal3 s 14072 6338 14170 6436 4 gnd
port 2 nsew
rlabel metal3 s 14061 6775 14159 6873 4 vdd
port 1 nsew
rlabel metal3 s 14182 7107 14280 7205 4 gnd
port 2 nsew
rlabel metal3 s 12819 7309 12917 7407 4 gnd
port 2 nsew
rlabel metal3 s 19178 5545 19276 5643 4 gnd
port 2 nsew
rlabel metal3 s 11690 5223 11788 5321 4 vdd
port 1 nsew
rlabel metal3 s 15315 7309 15413 7407 4 gnd
port 2 nsew
rlabel metal3 s 20307 7309 20405 7407 4 gnd
port 2 nsew
rlabel metal3 s 20321 7725 20419 7823 4 vdd
port 1 nsew
rlabel metal3 s 16557 6775 16655 6873 4 vdd
port 1 nsew
rlabel metal3 s 15320 6338 15418 6436 4 gnd
port 2 nsew
rlabel metal3 s 20426 5545 20524 5643 4 gnd
port 2 nsew
rlabel metal3 s 10317 6775 10415 6873 4 vdd
port 1 nsew
rlabel metal3 s 15434 5545 15532 5643 4 gnd
port 2 nsew
rlabel metal3 s 15430 7107 15528 7205 4 gnd
port 2 nsew
rlabel metal3 s 11565 6775 11663 6873 4 vdd
port 1 nsew
rlabel metal3 s 16682 5545 16780 5643 4 gnd
port 2 nsew
rlabel metal3 s 19073 7725 19171 7823 4 vdd
port 1 nsew
rlabel metal3 s 17930 5545 18028 5643 4 gnd
port 2 nsew
rlabel metal3 s 2829 6775 2927 6873 4 vdd
port 1 nsew
rlabel metal3 s 2954 5223 3052 5321 4 vdd
port 1 nsew
rlabel metal3 s 5336 6338 5434 6436 4 gnd
port 2 nsew
rlabel metal3 s 1587 7309 1685 7407 4 gnd
port 2 nsew
rlabel metal3 s 5331 7309 5429 7407 4 gnd
port 2 nsew
rlabel metal3 s 1702 7107 1800 7205 4 gnd
port 2 nsew
rlabel metal3 s 9194 5223 9292 5321 4 vdd
port 1 nsew
rlabel metal3 s 6573 6775 6671 6873 4 vdd
port 1 nsew
rlabel metal3 s 5446 7107 5544 7205 4 gnd
port 2 nsew
rlabel metal3 s 1581 6775 1679 6873 4 vdd
port 1 nsew
rlabel metal3 s 9080 6338 9178 6436 4 gnd
port 2 nsew
rlabel metal3 s 6593 7725 6691 7823 4 vdd
port 1 nsew
rlabel metal3 s 1601 7725 1699 7823 4 vdd
port 1 nsew
rlabel metal3 s 4202 5545 4300 5643 4 gnd
port 2 nsew
rlabel metal3 s 4083 7309 4181 7407 4 gnd
port 2 nsew
rlabel metal3 s 1706 5223 1804 5321 4 vdd
port 1 nsew
rlabel metal3 s 7841 7725 7939 7823 4 vdd
port 1 nsew
rlabel metal3 s 4198 7107 4296 7205 4 gnd
port 2 nsew
rlabel metal3 s 5450 5223 5548 5321 4 vdd
port 1 nsew
rlabel metal3 s 7827 7309 7925 7407 4 gnd
port 2 nsew
rlabel metal3 s 5325 6775 5423 6873 4 vdd
port 1 nsew
rlabel metal3 s 9075 7309 9173 7407 4 gnd
port 2 nsew
rlabel metal3 s 2950 7107 3048 7205 4 gnd
port 2 nsew
rlabel metal3 s 7946 5545 8044 5643 4 gnd
port 2 nsew
rlabel metal3 s 4077 6775 4175 6873 4 vdd
port 1 nsew
rlabel metal3 s 5345 7725 5443 7823 4 vdd
port 1 nsew
rlabel metal3 s 1706 5545 1804 5643 4 gnd
port 2 nsew
rlabel metal3 s 2849 7725 2947 7823 4 vdd
port 1 nsew
rlabel metal3 s 6698 5545 6796 5643 4 gnd
port 2 nsew
rlabel metal3 s 7821 6775 7919 6873 4 vdd
port 1 nsew
rlabel metal3 s 2954 5545 3052 5643 4 gnd
port 2 nsew
rlabel metal3 s 6584 6338 6682 6436 4 gnd
port 2 nsew
rlabel metal3 s 7942 7107 8040 7205 4 gnd
port 2 nsew
rlabel metal3 s 9069 6775 9167 6873 4 vdd
port 1 nsew
rlabel metal3 s -49 9288 49 9386 4 gnd
port 2 nsew
rlabel metal3 s 2835 7309 2933 7407 4 gnd
port 2 nsew
rlabel metal3 s 5450 5545 5548 5643 4 gnd
port 2 nsew
rlabel metal3 s 9190 7107 9288 7205 4 gnd
port 2 nsew
rlabel metal3 s 4088 6338 4186 6436 4 gnd
port 2 nsew
rlabel metal3 s 2840 6338 2938 6436 4 gnd
port 2 nsew
rlabel metal3 s 6579 7309 6677 7407 4 gnd
port 2 nsew
rlabel metal3 s -49 8168 49 8266 4 vdd
port 1 nsew
rlabel metal3 s 6694 7107 6792 7205 4 gnd
port 2 nsew
rlabel metal3 s 9089 7725 9187 7823 4 vdd
port 1 nsew
rlabel metal3 s 6698 5223 6796 5321 4 vdd
port 1 nsew
rlabel metal3 s 9194 5545 9292 5643 4 gnd
port 2 nsew
rlabel metal3 s 4097 7725 4195 7823 4 vdd
port 1 nsew
rlabel metal3 s 1592 6338 1690 6436 4 gnd
port 2 nsew
rlabel metal3 s 7946 5223 8044 5321 4 vdd
port 1 nsew
rlabel metal3 s 4202 5223 4300 5321 4 vdd
port 1 nsew
rlabel metal3 s 7832 6338 7930 6436 4 gnd
port 2 nsew
rlabel metal3 s 5693 1862 5791 1960 4 gnd
port 2 nsew
rlabel metal3 s 4445 1862 4543 1960 4 gnd
port 2 nsew
rlabel metal3 s 1949 1862 2047 1960 4 gnd
port 2 nsew
rlabel metal3 s 6768 3611 6866 3709 4 gnd
port 2 nsew
rlabel metal3 s 8016 3611 8114 3709 4 gnd
port 2 nsew
rlabel metal3 s 8189 1862 8287 1960 4 gnd
port 2 nsew
rlabel metal3 s 5438 4385 5536 4483 4 vdd
port 1 nsew
rlabel metal3 s 1776 3611 1874 3709 4 gnd
port 2 nsew
rlabel metal3 s 9182 4385 9280 4483 4 vdd
port 1 nsew
rlabel metal3 s 6686 4385 6784 4483 4 vdd
port 1 nsew
rlabel metal3 s 3197 1862 3295 1960 4 gnd
port 2 nsew
rlabel metal3 s 9264 3611 9362 3709 4 gnd
port 2 nsew
rlabel metal3 s 9437 1862 9535 1960 4 gnd
port 2 nsew
rlabel metal3 s 5520 3611 5618 3709 4 gnd
port 2 nsew
rlabel metal3 s 7934 4385 8032 4483 4 vdd
port 1 nsew
rlabel metal3 s 4190 4385 4288 4483 4 vdd
port 1 nsew
rlabel metal3 s 4272 3611 4370 3709 4 gnd
port 2 nsew
rlabel metal3 s 1694 4385 1792 4483 4 vdd
port 1 nsew
rlabel metal3 s 2942 4385 3040 4483 4 vdd
port 1 nsew
rlabel metal3 s 3024 3611 3122 3709 4 gnd
port 2 nsew
rlabel metal3 s 6941 1862 7039 1960 4 gnd
port 2 nsew
rlabel metal3 s 19421 1862 19519 1960 4 gnd
port 2 nsew
rlabel metal3 s 11760 3611 11858 3709 4 gnd
port 2 nsew
rlabel metal3 s 15422 4385 15520 4483 4 vdd
port 1 nsew
rlabel metal3 s 16925 1862 17023 1960 4 gnd
port 2 nsew
rlabel metal3 s 20414 4385 20512 4483 4 vdd
port 1 nsew
rlabel metal3 s 0 2762 41310 2822 4 sel_0
port 4 nsew
rlabel metal3 s 0 2638 41310 2698 4 sel_1
port 5 nsew
rlabel metal3 s 14429 1862 14527 1960 4 gnd
port 2 nsew
rlabel metal3 s 0 3478 40562 3538 4 s_en
port 6 nsew
rlabel metal3 s 11933 1862 12031 1960 4 gnd
port 2 nsew
rlabel metal3 s 14256 3611 14354 3709 4 gnd
port 2 nsew
rlabel metal3 s 20496 3611 20594 3709 4 gnd
port 2 nsew
rlabel metal3 s 10430 4385 10528 4483 4 vdd
port 1 nsew
rlabel metal3 s 15504 3611 15602 3709 4 gnd
port 2 nsew
rlabel metal3 s 12926 4385 13024 4483 4 vdd
port 1 nsew
rlabel metal3 s 10685 1862 10783 1960 4 gnd
port 2 nsew
rlabel metal3 s 19248 3611 19346 3709 4 gnd
port 2 nsew
rlabel metal3 s 16752 3611 16850 3709 4 gnd
port 2 nsew
rlabel metal3 s 18173 1862 18271 1960 4 gnd
port 2 nsew
rlabel metal3 s 14174 4385 14272 4483 4 vdd
port 1 nsew
rlabel metal3 s 16670 4385 16768 4483 4 vdd
port 1 nsew
rlabel metal3 s 11678 4385 11776 4483 4 vdd
port 1 nsew
rlabel metal3 s 17918 4385 18016 4483 4 vdd
port 1 nsew
rlabel metal3 s 15677 1862 15775 1960 4 gnd
port 2 nsew
rlabel metal3 s 13008 3611 13106 3709 4 gnd
port 2 nsew
rlabel metal3 s 19166 4385 19264 4483 4 vdd
port 1 nsew
rlabel metal3 s 13181 1862 13279 1960 4 gnd
port 2 nsew
rlabel metal3 s 0 951 41310 1011 4 p_en_bar
port 7 nsew
rlabel metal3 s 18000 3611 18098 3709 4 gnd
port 2 nsew
rlabel metal3 s 10512 3611 10610 3709 4 gnd
port 2 nsew
rlabel metal3 s 12364 313 12462 411 4 vdd
port 1 nsew
rlabel metal3 s 1132 313 1230 411 4 vdd
port 1 nsew
rlabel metal3 s 12750 313 12848 411 4 vdd
port 1 nsew
rlabel metal3 s 19852 313 19950 411 4 vdd
port 1 nsew
rlabel metal3 s 6124 313 6222 411 4 vdd
port 1 nsew
rlabel metal3 s 9868 313 9966 411 4 vdd
port 1 nsew
rlabel metal3 s 18604 313 18702 411 4 vdd
port 1 nsew
rlabel metal3 s 8620 313 8718 411 4 vdd
port 1 nsew
rlabel metal3 s 7758 313 7856 411 4 vdd
port 1 nsew
rlabel metal3 s 16494 313 16592 411 4 vdd
port 1 nsew
rlabel metal3 s 20238 313 20336 411 4 vdd
port 1 nsew
rlabel metal3 s 4014 313 4112 411 4 vdd
port 1 nsew
rlabel metal3 s 4876 313 4974 411 4 vdd
port 1 nsew
rlabel metal3 s 16108 313 16206 411 4 vdd
port 1 nsew
rlabel metal3 s 17356 313 17454 411 4 vdd
port 1 nsew
rlabel metal3 s 17742 313 17840 411 4 vdd
port 1 nsew
rlabel metal3 s 5262 313 5360 411 4 vdd
port 1 nsew
rlabel metal3 s 2380 313 2478 411 4 vdd
port 1 nsew
rlabel metal3 s 10254 313 10352 411 4 vdd
port 1 nsew
rlabel metal3 s 7372 313 7470 411 4 vdd
port 1 nsew
rlabel metal3 s 18990 313 19088 411 4 vdd
port 1 nsew
rlabel metal3 s 13998 313 14096 411 4 vdd
port 1 nsew
rlabel metal3 s 6510 313 6608 411 4 vdd
port 1 nsew
rlabel metal3 s 9006 313 9104 411 4 vdd
port 1 nsew
rlabel metal3 s 3628 313 3726 411 4 vdd
port 1 nsew
rlabel metal3 s 1518 313 1616 411 4 vdd
port 1 nsew
rlabel metal3 s 11502 313 11600 411 4 vdd
port 1 nsew
rlabel metal3 s 14860 313 14958 411 4 vdd
port 1 nsew
rlabel metal3 s 2766 313 2864 411 4 vdd
port 1 nsew
rlabel metal3 s 11116 313 11214 411 4 vdd
port 1 nsew
rlabel metal3 s 15246 313 15344 411 4 vdd
port 1 nsew
rlabel metal3 s 13612 313 13710 411 4 vdd
port 1 nsew
rlabel metal3 s 32332 313 32430 411 4 vdd
port 1 nsew
rlabel metal3 s 33966 313 34064 411 4 vdd
port 1 nsew
rlabel metal3 s 26478 313 26576 411 4 vdd
port 1 nsew
rlabel metal3 s 22348 313 22446 411 4 vdd
port 1 nsew
rlabel metal3 s 36462 313 36560 411 4 vdd
port 1 nsew
rlabel metal3 s 23982 313 24080 411 4 vdd
port 1 nsew
rlabel metal3 s 24844 313 24942 411 4 vdd
port 1 nsew
rlabel metal3 s 27726 313 27824 411 4 vdd
port 1 nsew
rlabel metal3 s 30222 313 30320 411 4 vdd
port 1 nsew
rlabel metal3 s 36076 313 36174 411 4 vdd
port 1 nsew
rlabel metal3 s 22734 313 22832 411 4 vdd
port 1 nsew
rlabel metal3 s 33580 313 33678 411 4 vdd
port 1 nsew
rlabel metal3 s 39820 313 39918 411 4 vdd
port 1 nsew
rlabel metal3 s 29836 313 29934 411 4 vdd
port 1 nsew
rlabel metal3 s 21100 313 21198 411 4 vdd
port 1 nsew
rlabel metal3 s 38572 313 38670 411 4 vdd
port 1 nsew
rlabel metal3 s 41068 313 41166 411 4 vdd
port 1 nsew
rlabel metal3 s 37710 313 37808 411 4 vdd
port 1 nsew
rlabel metal3 s 35214 313 35312 411 4 vdd
port 1 nsew
rlabel metal3 s 28588 313 28686 411 4 vdd
port 1 nsew
rlabel metal3 s 23596 313 23694 411 4 vdd
port 1 nsew
rlabel metal3 s 26092 313 26190 411 4 vdd
port 1 nsew
rlabel metal3 s 37324 313 37422 411 4 vdd
port 1 nsew
rlabel metal3 s 21486 313 21584 411 4 vdd
port 1 nsew
rlabel metal3 s 34828 313 34926 411 4 vdd
port 1 nsew
rlabel metal3 s 28974 313 29072 411 4 vdd
port 1 nsew
rlabel metal3 s 38958 313 39056 411 4 vdd
port 1 nsew
rlabel metal3 s 31470 313 31568 411 4 vdd
port 1 nsew
rlabel metal3 s 25230 313 25328 411 4 vdd
port 1 nsew
rlabel metal3 s 31084 313 31182 411 4 vdd
port 1 nsew
rlabel metal3 s 32718 313 32816 411 4 vdd
port 1 nsew
rlabel metal3 s 40206 313 40304 411 4 vdd
port 1 nsew
rlabel metal3 s 27340 313 27438 411 4 vdd
port 1 nsew
rlabel metal2 s 1360 9053 1388 9081 4 bank_wmask_0
port 8 nsew
rlabel metal2 s 11344 9053 11372 9081 4 bank_wmask_1
port 9 nsew
rlabel metal2 s 21328 9053 21356 9081 4 bank_wmask_2
port 10 nsew
rlabel metal2 s 31312 9053 31340 9081 4 bank_wmask_3
port 11 nsew
rlabel metal1 s 21441 7837 30801 7871 4 wdriver_sel_2
port 12 nsew
rlabel metal1 s 31425 7837 40785 7871 4 wdriver_sel_3
port 13 nsew
rlabel metal1 s 21597 7905 21657 7961 4 din_16
port 14 nsew
rlabel metal1 s 22845 7905 22905 7961 4 din_17
port 15 nsew
rlabel metal1 s 24093 7905 24153 7961 4 din_18
port 16 nsew
rlabel metal1 s 25341 7905 25401 7961 4 din_19
port 17 nsew
rlabel metal1 s 26589 7905 26649 7961 4 din_20
port 18 nsew
rlabel metal1 s 27837 7905 27897 7961 4 din_21
port 19 nsew
rlabel metal1 s 29085 7905 29145 7961 4 din_22
port 20 nsew
rlabel metal1 s 30333 7905 30393 7961 4 din_23
port 21 nsew
rlabel metal1 s 31581 7905 31641 7961 4 din_24
port 22 nsew
rlabel metal1 s 32829 7905 32889 7961 4 din_25
port 23 nsew
rlabel metal1 s 34077 7905 34137 7961 4 din_26
port 24 nsew
rlabel metal1 s 35325 7905 35385 7961 4 din_27
port 25 nsew
rlabel metal1 s 36573 7905 36633 7961 4 din_28
port 26 nsew
rlabel metal1 s 37821 7905 37881 7961 4 din_29
port 27 nsew
rlabel metal1 s 39069 7905 39129 7961 4 din_30
port 28 nsew
rlabel metal1 s 40317 7905 40377 7961 4 din_31
port 29 nsew
rlabel metal1 s 21446 5448 21492 5702 4 dout_16
port 30 nsew
rlabel metal1 s 22694 5448 22740 5702 4 dout_17
port 31 nsew
rlabel metal1 s 23942 5448 23988 5702 4 dout_18
port 32 nsew
rlabel metal1 s 25190 5448 25236 5702 4 dout_19
port 33 nsew
rlabel metal1 s 26438 5448 26484 5702 4 dout_20
port 34 nsew
rlabel metal1 s 27686 5448 27732 5702 4 dout_21
port 35 nsew
rlabel metal1 s 28934 5448 28980 5702 4 dout_22
port 36 nsew
rlabel metal1 s 30182 5448 30228 5702 4 dout_23
port 37 nsew
rlabel metal1 s 31430 5448 31476 5702 4 dout_24
port 38 nsew
rlabel metal1 s 32678 5448 32724 5702 4 dout_25
port 39 nsew
rlabel metal1 s 33926 5448 33972 5702 4 dout_26
port 40 nsew
rlabel metal1 s 35174 5448 35220 5702 4 dout_27
port 41 nsew
rlabel metal1 s 36422 5448 36468 5702 4 dout_28
port 42 nsew
rlabel metal1 s 37670 5448 37716 5702 4 dout_29
port 43 nsew
rlabel metal1 s 38918 5448 38964 5702 4 dout_30
port 44 nsew
rlabel metal1 s 40166 5448 40212 5702 4 dout_31
port 45 nsew
rlabel metal1 s 16605 7905 16665 7961 4 din_12
port 46 nsew
rlabel metal1 s 17853 7905 17913 7961 4 din_13
port 47 nsew
rlabel metal1 s 1478 5448 1524 5702 4 dout_0
port 48 nsew
rlabel metal1 s 2726 5448 2772 5702 4 dout_1
port 49 nsew
rlabel metal1 s 3974 5448 4020 5702 4 dout_2
port 50 nsew
rlabel metal1 s 5222 5448 5268 5702 4 dout_3
port 51 nsew
rlabel metal1 s 6470 5448 6516 5702 4 dout_4
port 52 nsew
rlabel metal1 s 7718 5448 7764 5702 4 dout_5
port 53 nsew
rlabel metal1 s 8966 5448 9012 5702 4 dout_6
port 54 nsew
rlabel metal1 s 10214 5448 10260 5702 4 dout_7
port 55 nsew
rlabel metal1 s 11462 5448 11508 5702 4 dout_8
port 56 nsew
rlabel metal1 s 12710 5448 12756 5702 4 dout_9
port 57 nsew
rlabel metal1 s 13958 5448 14004 5702 4 dout_10
port 58 nsew
rlabel metal1 s 15206 5448 15252 5702 4 dout_11
port 59 nsew
rlabel metal1 s 16454 5448 16500 5702 4 dout_12
port 60 nsew
rlabel metal1 s 17702 5448 17748 5702 4 dout_13
port 61 nsew
rlabel metal1 s 18950 5448 18996 5702 4 dout_14
port 62 nsew
rlabel metal1 s 20198 5448 20244 5702 4 dout_15
port 63 nsew
rlabel metal1 s 19101 7905 19161 7961 4 din_14
port 64 nsew
rlabel metal1 s 20349 7905 20409 7961 4 din_15
port 65 nsew
rlabel metal1 s 1473 7837 10833 7871 4 wdriver_sel_0
port 66 nsew
rlabel metal1 s 11457 7837 20817 7871 4 wdriver_sel_1
port 67 nsew
rlabel metal1 s 1629 7905 1689 7961 4 din_0
port 68 nsew
rlabel metal1 s 2877 7905 2937 7961 4 din_1
port 69 nsew
rlabel metal1 s 4125 7905 4185 7961 4 din_2
port 70 nsew
rlabel metal1 s 5373 7905 5433 7961 4 din_3
port 71 nsew
rlabel metal1 s 6621 7905 6681 7961 4 din_4
port 72 nsew
rlabel metal1 s 7869 7905 7929 7961 4 din_5
port 73 nsew
rlabel metal1 s 9117 7905 9177 7961 4 din_6
port 74 nsew
rlabel metal1 s 10365 7905 10425 7961 4 din_7
port 75 nsew
rlabel metal1 s 11613 7905 11673 7961 4 din_8
port 76 nsew
rlabel metal1 s 12861 7905 12921 7961 4 din_9
port 77 nsew
rlabel metal1 s 14109 7905 14169 7961 4 din_10
port 78 nsew
rlabel metal1 s 15357 7905 15417 7961 4 din_11
port 79 nsew
rlabel metal1 s 1280 252 1308 1006 4 rbl_bl
port 80 nsew
rlabel metal1 s 816 252 844 1006 4 rbl_br
port 81 nsew
rlabel metal1 s 1440 252 1468 1006 4 bl_0
port 82 nsew
rlabel metal1 s 1904 252 1932 1006 4 br_0
port 83 nsew
rlabel metal1 s 2528 252 2556 1006 4 bl_1
port 84 nsew
rlabel metal1 s 2064 252 2092 1006 4 br_1
port 85 nsew
rlabel metal1 s 2688 252 2716 1006 4 bl_2
port 86 nsew
rlabel metal1 s 3152 252 3180 1006 4 br_2
port 87 nsew
rlabel metal1 s 3776 252 3804 1006 4 bl_3
port 88 nsew
rlabel metal1 s 3312 252 3340 1006 4 br_3
port 89 nsew
rlabel metal1 s 3936 252 3964 1006 4 bl_4
port 90 nsew
rlabel metal1 s 4400 252 4428 1006 4 br_4
port 91 nsew
rlabel metal1 s 5024 252 5052 1006 4 bl_5
port 92 nsew
rlabel metal1 s 4560 252 4588 1006 4 br_5
port 93 nsew
rlabel metal1 s 5184 252 5212 1006 4 bl_6
port 94 nsew
rlabel metal1 s 5648 252 5676 1006 4 br_6
port 95 nsew
rlabel metal1 s 6272 252 6300 1006 4 bl_7
port 96 nsew
rlabel metal1 s 5808 252 5836 1006 4 br_7
port 97 nsew
rlabel metal1 s 6432 252 6460 1006 4 bl_8
port 98 nsew
rlabel metal1 s 6896 252 6924 1006 4 br_8
port 99 nsew
rlabel metal1 s 7520 252 7548 1006 4 bl_9
port 100 nsew
rlabel metal1 s 7056 252 7084 1006 4 br_9
port 101 nsew
rlabel metal1 s 7680 252 7708 1006 4 bl_10
port 102 nsew
rlabel metal1 s 8144 252 8172 1006 4 br_10
port 103 nsew
rlabel metal1 s 8768 252 8796 1006 4 bl_11
port 104 nsew
rlabel metal1 s 8304 252 8332 1006 4 br_11
port 105 nsew
rlabel metal1 s 8928 252 8956 1006 4 bl_12
port 106 nsew
rlabel metal1 s 9392 252 9420 1006 4 br_12
port 107 nsew
rlabel metal1 s 10016 252 10044 1006 4 bl_13
port 108 nsew
rlabel metal1 s 9552 252 9580 1006 4 br_13
port 109 nsew
rlabel metal1 s 10176 252 10204 1006 4 bl_14
port 110 nsew
rlabel metal1 s 10640 252 10668 1006 4 br_14
port 111 nsew
rlabel metal1 s 11264 252 11292 1006 4 bl_15
port 112 nsew
rlabel metal1 s 10800 252 10828 1006 4 br_15
port 113 nsew
rlabel metal1 s 11424 252 11452 1006 4 bl_16
port 114 nsew
rlabel metal1 s 11888 252 11916 1006 4 br_16
port 115 nsew
rlabel metal1 s 12512 252 12540 1006 4 bl_17
port 116 nsew
rlabel metal1 s 12048 252 12076 1006 4 br_17
port 117 nsew
rlabel metal1 s 12672 252 12700 1006 4 bl_18
port 118 nsew
rlabel metal1 s 13136 252 13164 1006 4 br_18
port 119 nsew
rlabel metal1 s 13760 252 13788 1006 4 bl_19
port 120 nsew
rlabel metal1 s 13296 252 13324 1006 4 br_19
port 121 nsew
rlabel metal1 s 13920 252 13948 1006 4 bl_20
port 122 nsew
rlabel metal1 s 14384 252 14412 1006 4 br_20
port 123 nsew
rlabel metal1 s 15008 252 15036 1006 4 bl_21
port 124 nsew
rlabel metal1 s 14544 252 14572 1006 4 br_21
port 125 nsew
rlabel metal1 s 15168 252 15196 1006 4 bl_22
port 126 nsew
rlabel metal1 s 15632 252 15660 1006 4 br_22
port 127 nsew
rlabel metal1 s 16256 252 16284 1006 4 bl_23
port 128 nsew
rlabel metal1 s 15792 252 15820 1006 4 br_23
port 129 nsew
rlabel metal1 s 16416 252 16444 1006 4 bl_24
port 130 nsew
rlabel metal1 s 16880 252 16908 1006 4 br_24
port 131 nsew
rlabel metal1 s 17504 252 17532 1006 4 bl_25
port 132 nsew
rlabel metal1 s 17040 252 17068 1006 4 br_25
port 133 nsew
rlabel metal1 s 17664 252 17692 1006 4 bl_26
port 134 nsew
rlabel metal1 s 18128 252 18156 1006 4 br_26
port 135 nsew
rlabel metal1 s 18752 252 18780 1006 4 bl_27
port 136 nsew
rlabel metal1 s 18288 252 18316 1006 4 br_27
port 137 nsew
rlabel metal1 s 18912 252 18940 1006 4 bl_28
port 138 nsew
rlabel metal1 s 19376 252 19404 1006 4 br_28
port 139 nsew
rlabel metal1 s 20000 252 20028 1006 4 bl_29
port 140 nsew
rlabel metal1 s 19536 252 19564 1006 4 br_29
port 141 nsew
rlabel metal1 s 20160 252 20188 1006 4 bl_30
port 142 nsew
rlabel metal1 s 20624 252 20652 1006 4 br_30
port 143 nsew
rlabel metal1 s 20784 252 20812 1006 4 br_31
port 144 nsew
rlabel metal1 s 21248 252 21276 1006 4 bl_31
port 145 nsew
rlabel metal1 s 21408 252 21436 1006 4 bl_32
port 146 nsew
rlabel metal1 s 21872 252 21900 1006 4 br_32
port 147 nsew
rlabel metal1 s 22496 252 22524 1006 4 bl_33
port 148 nsew
rlabel metal1 s 22032 252 22060 1006 4 br_33
port 149 nsew
rlabel metal1 s 22656 252 22684 1006 4 bl_34
port 150 nsew
rlabel metal1 s 23120 252 23148 1006 4 br_34
port 151 nsew
rlabel metal1 s 23744 252 23772 1006 4 bl_35
port 152 nsew
rlabel metal1 s 23280 252 23308 1006 4 br_35
port 153 nsew
rlabel metal1 s 23904 252 23932 1006 4 bl_36
port 154 nsew
rlabel metal1 s 24368 252 24396 1006 4 br_36
port 155 nsew
rlabel metal1 s 24992 252 25020 1006 4 bl_37
port 156 nsew
rlabel metal1 s 24528 252 24556 1006 4 br_37
port 157 nsew
rlabel metal1 s 25152 252 25180 1006 4 bl_38
port 158 nsew
rlabel metal1 s 25616 252 25644 1006 4 br_38
port 159 nsew
rlabel metal1 s 26240 252 26268 1006 4 bl_39
port 160 nsew
rlabel metal1 s 25776 252 25804 1006 4 br_39
port 161 nsew
rlabel metal1 s 26400 252 26428 1006 4 bl_40
port 162 nsew
rlabel metal1 s 26864 252 26892 1006 4 br_40
port 163 nsew
rlabel metal1 s 27488 252 27516 1006 4 bl_41
port 164 nsew
rlabel metal1 s 27024 252 27052 1006 4 br_41
port 165 nsew
rlabel metal1 s 27648 252 27676 1006 4 bl_42
port 166 nsew
rlabel metal1 s 28112 252 28140 1006 4 br_42
port 167 nsew
rlabel metal1 s 28736 252 28764 1006 4 bl_43
port 168 nsew
rlabel metal1 s 28272 252 28300 1006 4 br_43
port 169 nsew
rlabel metal1 s 28896 252 28924 1006 4 bl_44
port 170 nsew
rlabel metal1 s 29360 252 29388 1006 4 br_44
port 171 nsew
rlabel metal1 s 29984 252 30012 1006 4 bl_45
port 172 nsew
rlabel metal1 s 29520 252 29548 1006 4 br_45
port 173 nsew
rlabel metal1 s 30144 252 30172 1006 4 bl_46
port 174 nsew
rlabel metal1 s 30608 252 30636 1006 4 br_46
port 175 nsew
rlabel metal1 s 31232 252 31260 1006 4 bl_47
port 176 nsew
rlabel metal1 s 30768 252 30796 1006 4 br_47
port 177 nsew
rlabel metal1 s 31392 252 31420 1006 4 bl_48
port 178 nsew
rlabel metal1 s 31856 252 31884 1006 4 br_48
port 179 nsew
rlabel metal1 s 32480 252 32508 1006 4 bl_49
port 180 nsew
rlabel metal1 s 32016 252 32044 1006 4 br_49
port 181 nsew
rlabel metal1 s 32640 252 32668 1006 4 bl_50
port 182 nsew
rlabel metal1 s 33104 252 33132 1006 4 br_50
port 183 nsew
rlabel metal1 s 33728 252 33756 1006 4 bl_51
port 184 nsew
rlabel metal1 s 33264 252 33292 1006 4 br_51
port 185 nsew
rlabel metal1 s 33888 252 33916 1006 4 bl_52
port 186 nsew
rlabel metal1 s 34352 252 34380 1006 4 br_52
port 187 nsew
rlabel metal1 s 34976 252 35004 1006 4 bl_53
port 188 nsew
rlabel metal1 s 34512 252 34540 1006 4 br_53
port 189 nsew
rlabel metal1 s 35136 252 35164 1006 4 bl_54
port 190 nsew
rlabel metal1 s 35600 252 35628 1006 4 br_54
port 191 nsew
rlabel metal1 s 36224 252 36252 1006 4 bl_55
port 192 nsew
rlabel metal1 s 35760 252 35788 1006 4 br_55
port 193 nsew
rlabel metal1 s 36384 252 36412 1006 4 bl_56
port 194 nsew
rlabel metal1 s 36848 252 36876 1006 4 br_56
port 195 nsew
rlabel metal1 s 37472 252 37500 1006 4 bl_57
port 196 nsew
rlabel metal1 s 37008 252 37036 1006 4 br_57
port 197 nsew
rlabel metal1 s 37632 252 37660 1006 4 bl_58
port 198 nsew
rlabel metal1 s 38096 252 38124 1006 4 br_58
port 199 nsew
rlabel metal1 s 38720 252 38748 1006 4 bl_59
port 200 nsew
rlabel metal1 s 38256 252 38284 1006 4 br_59
port 201 nsew
rlabel metal1 s 38880 252 38908 1006 4 bl_60
port 202 nsew
rlabel metal1 s 39344 252 39372 1006 4 br_60
port 203 nsew
rlabel metal1 s 39968 252 39996 1006 4 bl_61
port 204 nsew
rlabel metal1 s 39504 252 39532 1006 4 br_61
port 205 nsew
rlabel metal1 s 40128 252 40156 1006 4 bl_62
port 206 nsew
rlabel metal1 s 40592 252 40620 1006 4 br_62
port 207 nsew
rlabel metal1 s 41216 252 41244 1006 4 bl_63
port 208 nsew
rlabel metal1 s 40752 252 40780 1006 4 br_63
port 209 nsew
rlabel locali s 1952 8803 1952 8803 4 wdriver_sel_0
port 66 nsew
rlabel locali s 11936 8803 11936 8803 4 wdriver_sel_1
port 67 nsew
rlabel locali s 21920 8803 21920 8803 4 wdriver_sel_2
port 12 nsew
rlabel locali s 31904 8803 31904 8803 4 wdriver_sel_3
port 13 nsew
<< properties >>
string FIXED_BBOX 0 0 41310 9337
string GDS_END 6989624
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_32x256_8.gds
string GDS_START 6801110
<< end >>
