magic
tech sky130B
magscale 1 2
timestamp 1666199351
<< metal4 >>
rect 0 13600 4000 18593
rect 0 12410 4000 13300
rect 0 11240 4000 12130
rect 0 10874 4000 10940
rect 0 10218 4000 10814
rect 0 9266 4000 9862
rect 0 9140 4000 9206
rect 0 7910 4000 8840
rect 0 6940 4000 7630
rect 0 5970 4000 6660
rect 0 4760 4000 5690
rect 0 3550 4000 4480
rect 0 2580 4000 3270
rect 0 1370 4000 2300
rect 0 0 4000 1090
<< obsm4 >>
rect 0 34750 4000 39593
rect 0 13380 4000 13520
rect 0 12210 4000 12330
rect 0 11020 4000 11160
rect 0 9922 4000 10158
<< metal5 >>
rect 0 34750 4000 39593
rect 0 13600 4000 18590
rect 0 12430 4000 13280
rect 0 11260 4000 12110
rect 0 9140 4000 10940
rect 0 7930 4000 8820
rect 0 6960 4000 7610
rect 0 5990 4000 6640
rect 0 4780 4000 5670
rect 0 3570 4000 4460
rect 0 2600 4000 3250
rect 0 1390 4000 2280
rect 0 20 4000 1070
<< labels >>
rlabel metal4 s 0 10218 4000 10814 6 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel metal4 s 0 9266 4000 9862 6 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel metal5 s 0 9140 4000 10940 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 10874 4000 10940 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 9140 4000 9206 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 0 6960 4000 7610 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 6940 4000 7630 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 0 2600 4000 3250 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 0 2580 4000 3270 6 VDDA
port 4 nsew power bidirectional
rlabel metal5 s 0 5990 4000 6640 6 VSWITCH
port 5 nsew power bidirectional
rlabel metal4 s 0 5970 4000 6660 6 VSWITCH
port 5 nsew power bidirectional
rlabel metal5 s 0 12430 4000 13280 6 VDDIO_Q
port 6 nsew power bidirectional
rlabel metal4 s 0 12410 4000 13300 6 VDDIO_Q
port 6 nsew power bidirectional
rlabel metal5 s 0 20 4000 1070 6 VCCHIB
port 7 nsew power bidirectional
rlabel metal4 s 0 0 4000 1090 6 VCCHIB
port 7 nsew power bidirectional
rlabel metal5 s 0 13600 4000 18590 6 VDDIO
port 8 nsew power bidirectional
rlabel metal4 s 0 13600 4000 18593 6 VDDIO
port 8 nsew power bidirectional
rlabel metal5 s 0 3570 4000 4460 6 VDDIO
port 8 nsew power bidirectional
rlabel metal4 s 0 3550 4000 4480 6 VDDIO
port 8 nsew power bidirectional
rlabel metal5 s 0 1390 4000 2280 6 VCCD
port 9 nsew power bidirectional
rlabel metal4 s 0 1370 4000 2300 6 VCCD
port 9 nsew power bidirectional
rlabel metal5 s 0 4780 4000 5670 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 0 4760 4000 5690 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal5 s 0 34750 4000 39593 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal5 s 0 7930 4000 8820 6 VSSD
port 11 nsew ground bidirectional
rlabel metal4 s 0 7910 4000 8840 6 VSSD
port 11 nsew ground bidirectional
rlabel metal5 s 0 11260 4000 12110 6 VSSIO_Q
port 12 nsew ground bidirectional
rlabel metal4 s 0 11240 4000 12130 6 VSSIO_Q
port 12 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 4000 39593
string LEFclass PAD SPACER
string LEFview TRUE
string GDS_END 2323990
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io.gds
string GDS_START 2314726
<< end >>
