magic
tech sky130A
timestamp 1666199351
<< properties >>
string GDS_END 29662656
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 29662268
<< end >>
