magic
tech sky130A
magscale 1 2
timestamp 1666464484
<< nwell >>
rect -38 261 2062 582
<< pwell >>
rect 1 21 2000 203
rect 29 -17 63 21
<< locali >>
rect 526 289 1233 323
rect 526 255 560 289
rect 1199 255 1233 289
rect 85 215 560 255
rect 594 221 1148 255
rect 594 215 1000 221
rect 1199 215 1474 255
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 17 401 80 493
rect 114 435 164 527
rect 198 401 248 493
rect 282 435 332 527
rect 366 459 752 493
rect 366 401 416 459
rect 534 425 584 459
rect 17 357 416 401
rect 450 391 500 425
rect 618 391 668 425
rect 450 357 668 391
rect 702 359 752 459
rect 806 401 856 493
rect 890 435 940 527
rect 974 401 1024 493
rect 1058 435 1108 527
rect 1142 401 1192 493
rect 1226 435 1276 527
rect 1310 401 1360 493
rect 1394 435 1444 527
rect 1478 459 1886 493
rect 1478 401 1528 459
rect 806 357 1528 401
rect 450 323 484 357
rect 17 289 484 323
rect 1310 291 1360 357
rect 1576 333 1634 425
rect 1668 367 1718 459
rect 1752 333 1802 425
rect 1836 359 1886 459
rect 1576 325 1802 333
rect 1920 325 2007 493
rect 1452 289 1542 323
rect 1576 289 2007 325
rect 17 181 51 289
rect 1508 255 1542 289
rect 1508 221 1913 255
rect 1708 215 1913 221
rect 1030 181 1041 187
rect 17 147 676 181
rect 106 145 676 147
rect 17 17 72 113
rect 106 51 172 145
rect 206 17 240 111
rect 274 51 340 145
rect 374 17 408 111
rect 442 51 508 145
rect 542 17 576 111
rect 610 51 676 145
rect 710 17 764 179
rect 833 153 1041 181
rect 1075 153 1116 187
rect 833 129 1116 153
rect 1150 145 1536 181
rect 1570 153 1593 187
rect 1627 181 1661 187
rect 1947 181 2007 289
rect 1627 153 2007 181
rect 1570 147 2007 153
rect 1570 145 1726 147
rect 1150 95 1200 145
rect 798 51 1200 95
rect 1234 17 1268 111
rect 1302 51 1368 145
rect 1402 17 1436 111
rect 1470 51 1536 145
rect 1592 17 1626 111
rect 1660 51 1726 145
rect 1760 17 1794 111
rect 1828 51 1894 147
rect 1928 17 1962 111
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 1041 153 1075 187
rect 1593 153 1627 187
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
<< metal1 >>
rect 0 561 2024 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 0 496 2024 527
rect 1029 187 1087 193
rect 1029 153 1041 187
rect 1075 184 1087 187
rect 1581 187 1639 193
rect 1581 184 1593 187
rect 1075 156 1593 184
rect 1075 153 1087 156
rect 1029 147 1087 153
rect 1581 153 1593 156
rect 1627 153 1639 187
rect 1581 147 1639 153
rect 0 17 2024 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
rect 0 -48 2024 -17
<< obsm1 >>
rect 385 320 443 329
rect 1489 320 1547 329
rect 385 292 1547 320
rect 385 283 443 292
rect 1489 283 1547 292
<< labels >>
rlabel locali s 1199 215 1474 255 6 A
port 1 nsew signal input
rlabel locali s 1199 255 1233 289 6 A
port 1 nsew signal input
rlabel locali s 85 215 560 255 6 A
port 1 nsew signal input
rlabel locali s 526 255 560 289 6 A
port 1 nsew signal input
rlabel locali s 526 289 1233 323 6 A
port 1 nsew signal input
rlabel locali s 594 215 1000 221 6 B
port 2 nsew signal input
rlabel locali s 594 221 1148 255 6 B
port 2 nsew signal input
rlabel metal1 s 0 -48 2024 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 1 21 2000 203 6 VNB
port 4 nsew ground bidirectional
rlabel nwell s -38 261 2062 582 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 496 2024 592 6 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 1581 147 1639 156 6 X
port 7 nsew signal output
rlabel metal1 s 1029 147 1087 156 6 X
port 7 nsew signal output
rlabel metal1 s 1029 156 1639 184 6 X
port 7 nsew signal output
rlabel metal1 s 1581 184 1639 193 6 X
port 7 nsew signal output
rlabel metal1 s 1029 184 1087 193 6 X
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2024 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 661364
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 646958
<< end >>
