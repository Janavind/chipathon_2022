magic
tech sky130B
magscale 1 2
timestamp 1666199351
<< locali >>
rect 310 1322 402 1368
<< metal1 >>
rect 2496 8314 2549 8360
rect 13310 7954 13365 8287
rect 451 932 1620 1077
rect 11799 737 11831 795
rect 761 681 794 713
rect 6540 685 6596 718
rect 4107 173 5276 318
rect 14167 280 14252 332
rect 13921 168 14073 220
rect 14164 88 14240 140
rect 47 -1145 84 -1010
rect 166 -1151 207 -1005
rect 256 -1157 316 -1019
rect 374 -1157 415 -1015
<< metal2 >>
rect 4692 12367 7591 13421
rect 11116 10856 12657 11949
rect 11116 4023 12657 5116
rect 5376 3624 6558 3626
rect 5376 3568 5385 3624
rect 5441 3568 5471 3624
rect 5527 3568 5557 3624
rect 5613 3568 5643 3624
rect 5699 3568 5728 3624
rect 5784 3568 5813 3624
rect 5869 3568 5898 3624
rect 5954 3568 5983 3624
rect 6039 3568 6068 3624
rect 6124 3568 6153 3624
rect 6209 3568 6238 3624
rect 6294 3568 6323 3624
rect 6379 3568 6408 3624
rect 6464 3568 6493 3624
rect 6549 3568 6558 3624
rect 5376 3538 6558 3568
rect 5376 3482 5385 3538
rect 5441 3482 5471 3538
rect 5527 3482 5557 3538
rect 5613 3482 5643 3538
rect 5699 3482 5728 3538
rect 5784 3482 5813 3538
rect 5869 3482 5898 3538
rect 5954 3482 5983 3538
rect 6039 3482 6068 3538
rect 6124 3482 6153 3538
rect 6209 3482 6238 3538
rect 6294 3482 6323 3538
rect 6379 3482 6408 3538
rect 6464 3482 6493 3538
rect 6549 3482 6558 3538
rect 5376 3452 6558 3482
rect 5376 3396 5385 3452
rect 5441 3396 5471 3452
rect 5527 3396 5557 3452
rect 5613 3396 5643 3452
rect 5699 3396 5728 3452
rect 5784 3396 5813 3452
rect 5869 3396 5898 3452
rect 5954 3396 5983 3452
rect 6039 3396 6068 3452
rect 6124 3396 6153 3452
rect 6209 3396 6238 3452
rect 6294 3396 6323 3452
rect 6379 3396 6408 3452
rect 6464 3396 6493 3452
rect 6549 3396 6558 3452
rect 5376 3366 6558 3396
rect 5376 3310 5385 3366
rect 5441 3310 5471 3366
rect 5527 3310 5557 3366
rect 5613 3310 5643 3366
rect 5699 3310 5728 3366
rect 5784 3310 5813 3366
rect 5869 3310 5898 3366
rect 5954 3310 5983 3366
rect 6039 3310 6068 3366
rect 6124 3310 6153 3366
rect 6209 3310 6238 3366
rect 6294 3310 6323 3366
rect 6379 3310 6408 3366
rect 6464 3310 6493 3366
rect 6549 3310 6558 3366
rect 5376 3280 6558 3310
rect 5376 3224 5385 3280
rect 5441 3224 5471 3280
rect 5527 3224 5557 3280
rect 5613 3224 5643 3280
rect 5699 3224 5728 3280
rect 5784 3224 5813 3280
rect 5869 3224 5898 3280
rect 5954 3224 5983 3280
rect 6039 3224 6068 3280
rect 6124 3224 6153 3280
rect 6209 3224 6238 3280
rect 6294 3224 6323 3280
rect 6379 3224 6408 3280
rect 6464 3224 6493 3280
rect 6549 3224 6558 3280
rect 5376 3194 6558 3224
rect 5376 3138 5385 3194
rect 5441 3138 5471 3194
rect 5527 3138 5557 3194
rect 5613 3138 5643 3194
rect 5699 3138 5728 3194
rect 5784 3138 5813 3194
rect 5869 3138 5898 3194
rect 5954 3138 5983 3194
rect 6039 3138 6068 3194
rect 6124 3138 6153 3194
rect 6209 3138 6238 3194
rect 6294 3138 6323 3194
rect 6379 3138 6408 3194
rect 6464 3138 6493 3194
rect 6549 3138 6558 3194
rect 5376 3108 6558 3138
rect 5376 3052 5385 3108
rect 5441 3052 5471 3108
rect 5527 3052 5557 3108
rect 5613 3052 5643 3108
rect 5699 3052 5728 3108
rect 5784 3052 5813 3108
rect 5869 3052 5898 3108
rect 5954 3052 5983 3108
rect 6039 3052 6068 3108
rect 6124 3052 6153 3108
rect 6209 3052 6238 3108
rect 6294 3052 6323 3108
rect 6379 3052 6408 3108
rect 6464 3052 6493 3108
rect 6549 3052 6558 3108
rect 5376 3022 6558 3052
rect 5376 2966 5385 3022
rect 5441 2966 5471 3022
rect 5527 2966 5557 3022
rect 5613 2966 5643 3022
rect 5699 2966 5728 3022
rect 5784 2966 5813 3022
rect 5869 2966 5898 3022
rect 5954 2966 5983 3022
rect 6039 2966 6068 3022
rect 6124 2966 6153 3022
rect 6209 2966 6238 3022
rect 6294 2966 6323 3022
rect 6379 2966 6408 3022
rect 6464 2966 6493 3022
rect 6549 2966 6558 3022
rect 5376 2936 6558 2966
rect 5376 2880 5385 2936
rect 5441 2880 5471 2936
rect 5527 2880 5557 2936
rect 5613 2880 5643 2936
rect 5699 2880 5728 2936
rect 5784 2880 5813 2936
rect 5869 2880 5898 2936
rect 5954 2880 5983 2936
rect 6039 2880 6068 2936
rect 6124 2880 6153 2936
rect 6209 2880 6238 2936
rect 6294 2880 6323 2936
rect 6379 2880 6408 2936
rect 6464 2880 6493 2936
rect 6549 2880 6558 2936
rect 5376 2850 6558 2880
rect 5376 2794 5385 2850
rect 5441 2794 5471 2850
rect 5527 2794 5557 2850
rect 5613 2794 5643 2850
rect 5699 2794 5728 2850
rect 5784 2794 5813 2850
rect 5869 2794 5898 2850
rect 5954 2794 5983 2850
rect 6039 2794 6068 2850
rect 6124 2794 6153 2850
rect 6209 2794 6238 2850
rect 6294 2794 6323 2850
rect 6379 2794 6408 2850
rect 6464 2794 6493 2850
rect 6549 2794 6558 2850
rect 5376 2764 6558 2794
rect 5376 2708 5385 2764
rect 5441 2708 5471 2764
rect 5527 2708 5557 2764
rect 5613 2708 5643 2764
rect 5699 2708 5728 2764
rect 5784 2708 5813 2764
rect 5869 2708 5898 2764
rect 5954 2708 5983 2764
rect 6039 2708 6068 2764
rect 6124 2708 6153 2764
rect 6209 2708 6238 2764
rect 6294 2708 6323 2764
rect 6379 2708 6408 2764
rect 6464 2708 6493 2764
rect 6549 2708 6558 2764
rect 5376 2678 6558 2708
rect 5376 2622 5385 2678
rect 5441 2622 5471 2678
rect 5527 2622 5557 2678
rect 5613 2622 5643 2678
rect 5699 2622 5728 2678
rect 5784 2622 5813 2678
rect 5869 2622 5898 2678
rect 5954 2622 5983 2678
rect 6039 2622 6068 2678
rect 6124 2622 6153 2678
rect 6209 2622 6238 2678
rect 6294 2622 6323 2678
rect 6379 2622 6408 2678
rect 6464 2622 6493 2678
rect 6549 2622 6558 2678
rect 5376 2592 6558 2622
rect 5376 2536 5385 2592
rect 5441 2536 5471 2592
rect 5527 2536 5557 2592
rect 5613 2536 5643 2592
rect 5699 2536 5728 2592
rect 5784 2536 5813 2592
rect 5869 2536 5898 2592
rect 5954 2536 5983 2592
rect 6039 2536 6068 2592
rect 6124 2536 6153 2592
rect 6209 2536 6238 2592
rect 6294 2536 6323 2592
rect 6379 2536 6408 2592
rect 6464 2536 6493 2592
rect 6549 2536 6558 2592
rect 5376 2534 6558 2536
rect 6987 3624 8169 3626
rect 6987 3568 6996 3624
rect 7052 3568 7082 3624
rect 7138 3568 7168 3624
rect 7224 3568 7254 3624
rect 7310 3568 7339 3624
rect 7395 3568 7424 3624
rect 7480 3568 7509 3624
rect 7565 3568 7594 3624
rect 7650 3568 7679 3624
rect 7735 3568 7764 3624
rect 7820 3568 7849 3624
rect 7905 3568 7934 3624
rect 7990 3568 8019 3624
rect 8075 3568 8104 3624
rect 8160 3568 8169 3624
rect 6987 3538 8169 3568
rect 6987 3482 6996 3538
rect 7052 3482 7082 3538
rect 7138 3482 7168 3538
rect 7224 3482 7254 3538
rect 7310 3482 7339 3538
rect 7395 3482 7424 3538
rect 7480 3482 7509 3538
rect 7565 3482 7594 3538
rect 7650 3482 7679 3538
rect 7735 3482 7764 3538
rect 7820 3482 7849 3538
rect 7905 3482 7934 3538
rect 7990 3482 8019 3538
rect 8075 3482 8104 3538
rect 8160 3482 8169 3538
rect 6987 3452 8169 3482
rect 6987 3396 6996 3452
rect 7052 3396 7082 3452
rect 7138 3396 7168 3452
rect 7224 3396 7254 3452
rect 7310 3396 7339 3452
rect 7395 3396 7424 3452
rect 7480 3396 7509 3452
rect 7565 3396 7594 3452
rect 7650 3396 7679 3452
rect 7735 3396 7764 3452
rect 7820 3396 7849 3452
rect 7905 3396 7934 3452
rect 7990 3396 8019 3452
rect 8075 3396 8104 3452
rect 8160 3396 8169 3452
rect 6987 3366 8169 3396
rect 6987 3310 6996 3366
rect 7052 3310 7082 3366
rect 7138 3310 7168 3366
rect 7224 3310 7254 3366
rect 7310 3310 7339 3366
rect 7395 3310 7424 3366
rect 7480 3310 7509 3366
rect 7565 3310 7594 3366
rect 7650 3310 7679 3366
rect 7735 3310 7764 3366
rect 7820 3310 7849 3366
rect 7905 3310 7934 3366
rect 7990 3310 8019 3366
rect 8075 3310 8104 3366
rect 8160 3310 8169 3366
rect 6987 3280 8169 3310
rect 6987 3224 6996 3280
rect 7052 3224 7082 3280
rect 7138 3224 7168 3280
rect 7224 3224 7254 3280
rect 7310 3224 7339 3280
rect 7395 3224 7424 3280
rect 7480 3224 7509 3280
rect 7565 3224 7594 3280
rect 7650 3224 7679 3280
rect 7735 3224 7764 3280
rect 7820 3224 7849 3280
rect 7905 3224 7934 3280
rect 7990 3224 8019 3280
rect 8075 3224 8104 3280
rect 8160 3224 8169 3280
rect 6987 3194 8169 3224
rect 6987 3138 6996 3194
rect 7052 3138 7082 3194
rect 7138 3138 7168 3194
rect 7224 3138 7254 3194
rect 7310 3138 7339 3194
rect 7395 3138 7424 3194
rect 7480 3138 7509 3194
rect 7565 3138 7594 3194
rect 7650 3138 7679 3194
rect 7735 3138 7764 3194
rect 7820 3138 7849 3194
rect 7905 3138 7934 3194
rect 7990 3138 8019 3194
rect 8075 3138 8104 3194
rect 8160 3138 8169 3194
rect 6987 3108 8169 3138
rect 6987 3052 6996 3108
rect 7052 3052 7082 3108
rect 7138 3052 7168 3108
rect 7224 3052 7254 3108
rect 7310 3052 7339 3108
rect 7395 3052 7424 3108
rect 7480 3052 7509 3108
rect 7565 3052 7594 3108
rect 7650 3052 7679 3108
rect 7735 3052 7764 3108
rect 7820 3052 7849 3108
rect 7905 3052 7934 3108
rect 7990 3052 8019 3108
rect 8075 3052 8104 3108
rect 8160 3052 8169 3108
rect 6987 3022 8169 3052
rect 6987 2966 6996 3022
rect 7052 2966 7082 3022
rect 7138 2966 7168 3022
rect 7224 2966 7254 3022
rect 7310 2966 7339 3022
rect 7395 2966 7424 3022
rect 7480 2966 7509 3022
rect 7565 2966 7594 3022
rect 7650 2966 7679 3022
rect 7735 2966 7764 3022
rect 7820 2966 7849 3022
rect 7905 2966 7934 3022
rect 7990 2966 8019 3022
rect 8075 2966 8104 3022
rect 8160 2966 8169 3022
rect 6987 2936 8169 2966
rect 6987 2880 6996 2936
rect 7052 2880 7082 2936
rect 7138 2880 7168 2936
rect 7224 2880 7254 2936
rect 7310 2880 7339 2936
rect 7395 2880 7424 2936
rect 7480 2880 7509 2936
rect 7565 2880 7594 2936
rect 7650 2880 7679 2936
rect 7735 2880 7764 2936
rect 7820 2880 7849 2936
rect 7905 2880 7934 2936
rect 7990 2880 8019 2936
rect 8075 2880 8104 2936
rect 8160 2880 8169 2936
rect 6987 2850 8169 2880
rect 6987 2794 6996 2850
rect 7052 2794 7082 2850
rect 7138 2794 7168 2850
rect 7224 2794 7254 2850
rect 7310 2794 7339 2850
rect 7395 2794 7424 2850
rect 7480 2794 7509 2850
rect 7565 2794 7594 2850
rect 7650 2794 7679 2850
rect 7735 2794 7764 2850
rect 7820 2794 7849 2850
rect 7905 2794 7934 2850
rect 7990 2794 8019 2850
rect 8075 2794 8104 2850
rect 8160 2794 8169 2850
rect 6987 2764 8169 2794
rect 6987 2708 6996 2764
rect 7052 2708 7082 2764
rect 7138 2708 7168 2764
rect 7224 2708 7254 2764
rect 7310 2708 7339 2764
rect 7395 2708 7424 2764
rect 7480 2708 7509 2764
rect 7565 2708 7594 2764
rect 7650 2708 7679 2764
rect 7735 2708 7764 2764
rect 7820 2708 7849 2764
rect 7905 2708 7934 2764
rect 7990 2708 8019 2764
rect 8075 2708 8104 2764
rect 8160 2708 8169 2764
rect 6987 2678 8169 2708
rect 6987 2622 6996 2678
rect 7052 2622 7082 2678
rect 7138 2622 7168 2678
rect 7224 2622 7254 2678
rect 7310 2622 7339 2678
rect 7395 2622 7424 2678
rect 7480 2622 7509 2678
rect 7565 2622 7594 2678
rect 7650 2622 7679 2678
rect 7735 2622 7764 2678
rect 7820 2622 7849 2678
rect 7905 2622 7934 2678
rect 7990 2622 8019 2678
rect 8075 2622 8104 2678
rect 8160 2622 8169 2678
rect 6987 2592 8169 2622
rect 6987 2536 6996 2592
rect 7052 2536 7082 2592
rect 7138 2536 7168 2592
rect 7224 2536 7254 2592
rect 7310 2536 7339 2592
rect 7395 2536 7424 2592
rect 7480 2536 7509 2592
rect 7565 2536 7594 2592
rect 7650 2536 7679 2592
rect 7735 2536 7764 2592
rect 7820 2536 7849 2592
rect 7905 2536 7934 2592
rect 7990 2536 8019 2592
rect 8075 2536 8104 2592
rect 8160 2536 8169 2592
rect 6987 2534 8169 2536
rect 9167 3623 10359 3626
rect 9167 3567 9176 3623
rect 9232 3567 9262 3623
rect 9318 3567 9348 3623
rect 9404 3567 9434 3623
rect 9490 3567 9520 3623
rect 9576 3567 9606 3623
rect 9662 3567 9692 3623
rect 9748 3567 9778 3623
rect 9834 3567 9864 3623
rect 9920 3567 9950 3623
rect 10006 3567 10036 3623
rect 10092 3567 10122 3623
rect 10178 3567 10208 3623
rect 10264 3567 10294 3623
rect 10350 3567 10359 3623
rect 9167 3537 10359 3567
rect 9167 3481 9176 3537
rect 9232 3481 9262 3537
rect 9318 3481 9348 3537
rect 9404 3481 9434 3537
rect 9490 3481 9520 3537
rect 9576 3481 9606 3537
rect 9662 3481 9692 3537
rect 9748 3481 9778 3537
rect 9834 3481 9864 3537
rect 9920 3481 9950 3537
rect 10006 3481 10036 3537
rect 10092 3481 10122 3537
rect 10178 3481 10208 3537
rect 10264 3481 10294 3537
rect 10350 3481 10359 3537
rect 9167 3451 10359 3481
rect 9167 3395 9176 3451
rect 9232 3395 9262 3451
rect 9318 3395 9348 3451
rect 9404 3395 9434 3451
rect 9490 3395 9520 3451
rect 9576 3395 9606 3451
rect 9662 3395 9692 3451
rect 9748 3395 9778 3451
rect 9834 3395 9864 3451
rect 9920 3395 9950 3451
rect 10006 3395 10036 3451
rect 10092 3395 10122 3451
rect 10178 3395 10208 3451
rect 10264 3395 10294 3451
rect 10350 3395 10359 3451
rect 9167 3365 10359 3395
rect 9167 3309 9176 3365
rect 9232 3309 9262 3365
rect 9318 3309 9348 3365
rect 9404 3309 9434 3365
rect 9490 3309 9520 3365
rect 9576 3309 9606 3365
rect 9662 3309 9692 3365
rect 9748 3309 9778 3365
rect 9834 3309 9864 3365
rect 9920 3309 9950 3365
rect 10006 3309 10036 3365
rect 10092 3309 10122 3365
rect 10178 3309 10208 3365
rect 10264 3309 10294 3365
rect 10350 3309 10359 3365
rect 9167 3279 10359 3309
rect 9167 3223 9176 3279
rect 9232 3223 9262 3279
rect 9318 3223 9348 3279
rect 9404 3223 9434 3279
rect 9490 3223 9520 3279
rect 9576 3223 9606 3279
rect 9662 3223 9692 3279
rect 9748 3223 9778 3279
rect 9834 3223 9864 3279
rect 9920 3223 9950 3279
rect 10006 3223 10036 3279
rect 10092 3223 10122 3279
rect 10178 3223 10208 3279
rect 10264 3223 10294 3279
rect 10350 3223 10359 3279
rect 9167 3193 10359 3223
rect 9167 3137 9176 3193
rect 9232 3137 9262 3193
rect 9318 3137 9348 3193
rect 9404 3137 9434 3193
rect 9490 3137 9520 3193
rect 9576 3137 9606 3193
rect 9662 3137 9692 3193
rect 9748 3137 9778 3193
rect 9834 3137 9864 3193
rect 9920 3137 9950 3193
rect 10006 3137 10036 3193
rect 10092 3137 10122 3193
rect 10178 3137 10208 3193
rect 10264 3137 10294 3193
rect 10350 3137 10359 3193
rect 9167 3107 10359 3137
rect 9167 3051 9176 3107
rect 9232 3051 9262 3107
rect 9318 3051 9348 3107
rect 9404 3051 9434 3107
rect 9490 3051 9520 3107
rect 9576 3051 9606 3107
rect 9662 3051 9692 3107
rect 9748 3051 9778 3107
rect 9834 3051 9864 3107
rect 9920 3051 9950 3107
rect 10006 3051 10036 3107
rect 10092 3051 10122 3107
rect 10178 3051 10208 3107
rect 10264 3051 10294 3107
rect 10350 3051 10359 3107
rect 9167 3021 10359 3051
rect 9167 2965 9176 3021
rect 9232 2965 9262 3021
rect 9318 2965 9348 3021
rect 9404 2965 9434 3021
rect 9490 2965 9520 3021
rect 9576 2965 9606 3021
rect 9662 2965 9692 3021
rect 9748 2965 9778 3021
rect 9834 2965 9864 3021
rect 9920 2965 9950 3021
rect 10006 2965 10036 3021
rect 10092 2965 10122 3021
rect 10178 2965 10208 3021
rect 10264 2965 10294 3021
rect 10350 2965 10359 3021
rect 9167 2935 10359 2965
rect 9167 2879 9176 2935
rect 9232 2879 9262 2935
rect 9318 2879 9348 2935
rect 9404 2879 9434 2935
rect 9490 2879 9520 2935
rect 9576 2879 9606 2935
rect 9662 2879 9692 2935
rect 9748 2879 9778 2935
rect 9834 2879 9864 2935
rect 9920 2879 9950 2935
rect 10006 2879 10036 2935
rect 10092 2879 10122 2935
rect 10178 2879 10208 2935
rect 10264 2879 10294 2935
rect 10350 2879 10359 2935
rect 9167 2849 10359 2879
rect 9167 2793 9176 2849
rect 9232 2793 9262 2849
rect 9318 2793 9348 2849
rect 9404 2793 9434 2849
rect 9490 2793 9520 2849
rect 9576 2793 9606 2849
rect 9662 2793 9692 2849
rect 9748 2793 9778 2849
rect 9834 2793 9864 2849
rect 9920 2793 9950 2849
rect 10006 2793 10036 2849
rect 10092 2793 10122 2849
rect 10178 2793 10208 2849
rect 10264 2793 10294 2849
rect 10350 2793 10359 2849
rect 9167 2763 10359 2793
rect 9167 2707 9176 2763
rect 9232 2707 9262 2763
rect 9318 2707 9348 2763
rect 9404 2707 9434 2763
rect 9490 2707 9520 2763
rect 9576 2707 9606 2763
rect 9662 2707 9692 2763
rect 9748 2707 9778 2763
rect 9834 2707 9864 2763
rect 9920 2707 9950 2763
rect 10006 2707 10036 2763
rect 10092 2707 10122 2763
rect 10178 2707 10208 2763
rect 10264 2707 10294 2763
rect 10350 2707 10359 2763
rect 9167 2677 10359 2707
rect 9167 2621 9176 2677
rect 9232 2621 9262 2677
rect 9318 2621 9348 2677
rect 9404 2621 9434 2677
rect 9490 2621 9520 2677
rect 9576 2621 9606 2677
rect 9662 2621 9692 2677
rect 9748 2621 9778 2677
rect 9834 2621 9864 2677
rect 9920 2621 9950 2677
rect 10006 2621 10036 2677
rect 10092 2621 10122 2677
rect 10178 2621 10208 2677
rect 10264 2621 10294 2677
rect 10350 2621 10359 2677
rect 9167 2591 10359 2621
rect 9167 2535 9176 2591
rect 9232 2535 9262 2591
rect 9318 2535 9348 2591
rect 9404 2535 9434 2591
rect 9490 2535 9520 2591
rect 9576 2535 9606 2591
rect 9662 2535 9692 2591
rect 9748 2535 9778 2591
rect 9834 2535 9864 2591
rect 9920 2535 9950 2591
rect 10006 2535 10036 2591
rect 10092 2535 10122 2591
rect 10178 2535 10208 2591
rect 10264 2535 10294 2591
rect 10350 2535 10359 2591
rect 9167 2532 10359 2535
rect 10659 3623 11854 3626
rect 10659 3567 10668 3623
rect 10724 3567 10749 3623
rect 10805 3567 10829 3623
rect 10885 3567 10909 3623
rect 10965 3567 10989 3623
rect 11045 3567 11069 3623
rect 11125 3567 11149 3623
rect 11205 3567 11229 3623
rect 11285 3567 11309 3623
rect 11365 3567 11389 3623
rect 11445 3567 11469 3623
rect 11525 3567 11549 3623
rect 11605 3567 11629 3623
rect 11685 3567 11709 3623
rect 11765 3567 11789 3623
rect 11845 3567 11854 3623
rect 10659 3537 11854 3567
rect 10659 3481 10668 3537
rect 10724 3481 10749 3537
rect 10805 3481 10829 3537
rect 10885 3481 10909 3537
rect 10965 3481 10989 3537
rect 11045 3481 11069 3537
rect 11125 3481 11149 3537
rect 11205 3481 11229 3537
rect 11285 3481 11309 3537
rect 11365 3481 11389 3537
rect 11445 3481 11469 3537
rect 11525 3481 11549 3537
rect 11605 3481 11629 3537
rect 11685 3481 11709 3537
rect 11765 3481 11789 3537
rect 11845 3481 11854 3537
rect 10659 3451 11854 3481
rect 10659 3395 10668 3451
rect 10724 3395 10749 3451
rect 10805 3395 10829 3451
rect 10885 3395 10909 3451
rect 10965 3395 10989 3451
rect 11045 3395 11069 3451
rect 11125 3395 11149 3451
rect 11205 3395 11229 3451
rect 11285 3395 11309 3451
rect 11365 3395 11389 3451
rect 11445 3395 11469 3451
rect 11525 3395 11549 3451
rect 11605 3395 11629 3451
rect 11685 3395 11709 3451
rect 11765 3395 11789 3451
rect 11845 3395 11854 3451
rect 10659 3365 11854 3395
rect 10659 3309 10668 3365
rect 10724 3309 10749 3365
rect 10805 3309 10829 3365
rect 10885 3309 10909 3365
rect 10965 3309 10989 3365
rect 11045 3309 11069 3365
rect 11125 3309 11149 3365
rect 11205 3309 11229 3365
rect 11285 3309 11309 3365
rect 11365 3309 11389 3365
rect 11445 3309 11469 3365
rect 11525 3309 11549 3365
rect 11605 3309 11629 3365
rect 11685 3309 11709 3365
rect 11765 3309 11789 3365
rect 11845 3309 11854 3365
rect 10659 3279 11854 3309
rect 10659 3223 10668 3279
rect 10724 3223 10749 3279
rect 10805 3223 10829 3279
rect 10885 3223 10909 3279
rect 10965 3223 10989 3279
rect 11045 3223 11069 3279
rect 11125 3223 11149 3279
rect 11205 3223 11229 3279
rect 11285 3223 11309 3279
rect 11365 3223 11389 3279
rect 11445 3223 11469 3279
rect 11525 3223 11549 3279
rect 11605 3223 11629 3279
rect 11685 3223 11709 3279
rect 11765 3223 11789 3279
rect 11845 3223 11854 3279
rect 10659 3193 11854 3223
rect 10659 3137 10668 3193
rect 10724 3137 10749 3193
rect 10805 3137 10829 3193
rect 10885 3137 10909 3193
rect 10965 3137 10989 3193
rect 11045 3137 11069 3193
rect 11125 3137 11149 3193
rect 11205 3137 11229 3193
rect 11285 3137 11309 3193
rect 11365 3137 11389 3193
rect 11445 3137 11469 3193
rect 11525 3137 11549 3193
rect 11605 3137 11629 3193
rect 11685 3137 11709 3193
rect 11765 3137 11789 3193
rect 11845 3137 11854 3193
rect 10659 3107 11854 3137
rect 10659 3051 10668 3107
rect 10724 3051 10749 3107
rect 10805 3051 10829 3107
rect 10885 3051 10909 3107
rect 10965 3051 10989 3107
rect 11045 3051 11069 3107
rect 11125 3051 11149 3107
rect 11205 3051 11229 3107
rect 11285 3051 11309 3107
rect 11365 3051 11389 3107
rect 11445 3051 11469 3107
rect 11525 3051 11549 3107
rect 11605 3051 11629 3107
rect 11685 3051 11709 3107
rect 11765 3051 11789 3107
rect 11845 3051 11854 3107
rect 10659 3021 11854 3051
rect 10659 2965 10668 3021
rect 10724 2965 10749 3021
rect 10805 2965 10829 3021
rect 10885 2965 10909 3021
rect 10965 2965 10989 3021
rect 11045 2965 11069 3021
rect 11125 2965 11149 3021
rect 11205 2965 11229 3021
rect 11285 2965 11309 3021
rect 11365 2965 11389 3021
rect 11445 2965 11469 3021
rect 11525 2965 11549 3021
rect 11605 2965 11629 3021
rect 11685 2965 11709 3021
rect 11765 2965 11789 3021
rect 11845 2965 11854 3021
rect 10659 2935 11854 2965
rect 10659 2879 10668 2935
rect 10724 2879 10749 2935
rect 10805 2879 10829 2935
rect 10885 2879 10909 2935
rect 10965 2879 10989 2935
rect 11045 2879 11069 2935
rect 11125 2879 11149 2935
rect 11205 2879 11229 2935
rect 11285 2879 11309 2935
rect 11365 2879 11389 2935
rect 11445 2879 11469 2935
rect 11525 2879 11549 2935
rect 11605 2879 11629 2935
rect 11685 2879 11709 2935
rect 11765 2879 11789 2935
rect 11845 2879 11854 2935
rect 10659 2849 11854 2879
rect 10659 2793 10668 2849
rect 10724 2793 10749 2849
rect 10805 2793 10829 2849
rect 10885 2793 10909 2849
rect 10965 2793 10989 2849
rect 11045 2793 11069 2849
rect 11125 2793 11149 2849
rect 11205 2793 11229 2849
rect 11285 2793 11309 2849
rect 11365 2793 11389 2849
rect 11445 2793 11469 2849
rect 11525 2793 11549 2849
rect 11605 2793 11629 2849
rect 11685 2793 11709 2849
rect 11765 2793 11789 2849
rect 11845 2793 11854 2849
rect 10659 2763 11854 2793
rect 10659 2707 10668 2763
rect 10724 2707 10749 2763
rect 10805 2707 10829 2763
rect 10885 2707 10909 2763
rect 10965 2707 10989 2763
rect 11045 2707 11069 2763
rect 11125 2707 11149 2763
rect 11205 2707 11229 2763
rect 11285 2707 11309 2763
rect 11365 2707 11389 2763
rect 11445 2707 11469 2763
rect 11525 2707 11549 2763
rect 11605 2707 11629 2763
rect 11685 2707 11709 2763
rect 11765 2707 11789 2763
rect 11845 2707 11854 2763
rect 10659 2677 11854 2707
rect 10659 2621 10668 2677
rect 10724 2621 10749 2677
rect 10805 2621 10829 2677
rect 10885 2621 10909 2677
rect 10965 2621 10989 2677
rect 11045 2621 11069 2677
rect 11125 2621 11149 2677
rect 11205 2621 11229 2677
rect 11285 2621 11309 2677
rect 11365 2621 11389 2677
rect 11445 2621 11469 2677
rect 11525 2621 11549 2677
rect 11605 2621 11629 2677
rect 11685 2621 11709 2677
rect 11765 2621 11789 2677
rect 11845 2621 11854 2677
rect 10659 2591 11854 2621
rect 10659 2535 10668 2591
rect 10724 2535 10749 2591
rect 10805 2535 10829 2591
rect 10885 2535 10909 2591
rect 10965 2535 10989 2591
rect 11045 2535 11069 2591
rect 11125 2535 11149 2591
rect 11205 2535 11229 2591
rect 11285 2535 11309 2591
rect 11365 2535 11389 2591
rect 11445 2535 11469 2591
rect 11525 2535 11549 2591
rect 11605 2535 11629 2591
rect 11685 2535 11709 2591
rect 11765 2535 11789 2591
rect 11845 2535 11854 2591
rect 13327 2545 14496 3616
rect 10659 2532 11854 2535
rect 14708 -6 14748 186
rect 14788 -6 14828 186
rect 14868 -6 14908 186
rect 14948 -6 14988 186
rect 15028 -6 15068 186
<< via2 >>
rect 5385 3568 5441 3624
rect 5471 3568 5527 3624
rect 5557 3568 5613 3624
rect 5643 3568 5699 3624
rect 5728 3568 5784 3624
rect 5813 3568 5869 3624
rect 5898 3568 5954 3624
rect 5983 3568 6039 3624
rect 6068 3568 6124 3624
rect 6153 3568 6209 3624
rect 6238 3568 6294 3624
rect 6323 3568 6379 3624
rect 6408 3568 6464 3624
rect 6493 3568 6549 3624
rect 5385 3482 5441 3538
rect 5471 3482 5527 3538
rect 5557 3482 5613 3538
rect 5643 3482 5699 3538
rect 5728 3482 5784 3538
rect 5813 3482 5869 3538
rect 5898 3482 5954 3538
rect 5983 3482 6039 3538
rect 6068 3482 6124 3538
rect 6153 3482 6209 3538
rect 6238 3482 6294 3538
rect 6323 3482 6379 3538
rect 6408 3482 6464 3538
rect 6493 3482 6549 3538
rect 5385 3396 5441 3452
rect 5471 3396 5527 3452
rect 5557 3396 5613 3452
rect 5643 3396 5699 3452
rect 5728 3396 5784 3452
rect 5813 3396 5869 3452
rect 5898 3396 5954 3452
rect 5983 3396 6039 3452
rect 6068 3396 6124 3452
rect 6153 3396 6209 3452
rect 6238 3396 6294 3452
rect 6323 3396 6379 3452
rect 6408 3396 6464 3452
rect 6493 3396 6549 3452
rect 5385 3310 5441 3366
rect 5471 3310 5527 3366
rect 5557 3310 5613 3366
rect 5643 3310 5699 3366
rect 5728 3310 5784 3366
rect 5813 3310 5869 3366
rect 5898 3310 5954 3366
rect 5983 3310 6039 3366
rect 6068 3310 6124 3366
rect 6153 3310 6209 3366
rect 6238 3310 6294 3366
rect 6323 3310 6379 3366
rect 6408 3310 6464 3366
rect 6493 3310 6549 3366
rect 5385 3224 5441 3280
rect 5471 3224 5527 3280
rect 5557 3224 5613 3280
rect 5643 3224 5699 3280
rect 5728 3224 5784 3280
rect 5813 3224 5869 3280
rect 5898 3224 5954 3280
rect 5983 3224 6039 3280
rect 6068 3224 6124 3280
rect 6153 3224 6209 3280
rect 6238 3224 6294 3280
rect 6323 3224 6379 3280
rect 6408 3224 6464 3280
rect 6493 3224 6549 3280
rect 5385 3138 5441 3194
rect 5471 3138 5527 3194
rect 5557 3138 5613 3194
rect 5643 3138 5699 3194
rect 5728 3138 5784 3194
rect 5813 3138 5869 3194
rect 5898 3138 5954 3194
rect 5983 3138 6039 3194
rect 6068 3138 6124 3194
rect 6153 3138 6209 3194
rect 6238 3138 6294 3194
rect 6323 3138 6379 3194
rect 6408 3138 6464 3194
rect 6493 3138 6549 3194
rect 5385 3052 5441 3108
rect 5471 3052 5527 3108
rect 5557 3052 5613 3108
rect 5643 3052 5699 3108
rect 5728 3052 5784 3108
rect 5813 3052 5869 3108
rect 5898 3052 5954 3108
rect 5983 3052 6039 3108
rect 6068 3052 6124 3108
rect 6153 3052 6209 3108
rect 6238 3052 6294 3108
rect 6323 3052 6379 3108
rect 6408 3052 6464 3108
rect 6493 3052 6549 3108
rect 5385 2966 5441 3022
rect 5471 2966 5527 3022
rect 5557 2966 5613 3022
rect 5643 2966 5699 3022
rect 5728 2966 5784 3022
rect 5813 2966 5869 3022
rect 5898 2966 5954 3022
rect 5983 2966 6039 3022
rect 6068 2966 6124 3022
rect 6153 2966 6209 3022
rect 6238 2966 6294 3022
rect 6323 2966 6379 3022
rect 6408 2966 6464 3022
rect 6493 2966 6549 3022
rect 5385 2880 5441 2936
rect 5471 2880 5527 2936
rect 5557 2880 5613 2936
rect 5643 2880 5699 2936
rect 5728 2880 5784 2936
rect 5813 2880 5869 2936
rect 5898 2880 5954 2936
rect 5983 2880 6039 2936
rect 6068 2880 6124 2936
rect 6153 2880 6209 2936
rect 6238 2880 6294 2936
rect 6323 2880 6379 2936
rect 6408 2880 6464 2936
rect 6493 2880 6549 2936
rect 5385 2794 5441 2850
rect 5471 2794 5527 2850
rect 5557 2794 5613 2850
rect 5643 2794 5699 2850
rect 5728 2794 5784 2850
rect 5813 2794 5869 2850
rect 5898 2794 5954 2850
rect 5983 2794 6039 2850
rect 6068 2794 6124 2850
rect 6153 2794 6209 2850
rect 6238 2794 6294 2850
rect 6323 2794 6379 2850
rect 6408 2794 6464 2850
rect 6493 2794 6549 2850
rect 5385 2708 5441 2764
rect 5471 2708 5527 2764
rect 5557 2708 5613 2764
rect 5643 2708 5699 2764
rect 5728 2708 5784 2764
rect 5813 2708 5869 2764
rect 5898 2708 5954 2764
rect 5983 2708 6039 2764
rect 6068 2708 6124 2764
rect 6153 2708 6209 2764
rect 6238 2708 6294 2764
rect 6323 2708 6379 2764
rect 6408 2708 6464 2764
rect 6493 2708 6549 2764
rect 5385 2622 5441 2678
rect 5471 2622 5527 2678
rect 5557 2622 5613 2678
rect 5643 2622 5699 2678
rect 5728 2622 5784 2678
rect 5813 2622 5869 2678
rect 5898 2622 5954 2678
rect 5983 2622 6039 2678
rect 6068 2622 6124 2678
rect 6153 2622 6209 2678
rect 6238 2622 6294 2678
rect 6323 2622 6379 2678
rect 6408 2622 6464 2678
rect 6493 2622 6549 2678
rect 5385 2536 5441 2592
rect 5471 2536 5527 2592
rect 5557 2536 5613 2592
rect 5643 2536 5699 2592
rect 5728 2536 5784 2592
rect 5813 2536 5869 2592
rect 5898 2536 5954 2592
rect 5983 2536 6039 2592
rect 6068 2536 6124 2592
rect 6153 2536 6209 2592
rect 6238 2536 6294 2592
rect 6323 2536 6379 2592
rect 6408 2536 6464 2592
rect 6493 2536 6549 2592
rect 6996 3568 7052 3624
rect 7082 3568 7138 3624
rect 7168 3568 7224 3624
rect 7254 3568 7310 3624
rect 7339 3568 7395 3624
rect 7424 3568 7480 3624
rect 7509 3568 7565 3624
rect 7594 3568 7650 3624
rect 7679 3568 7735 3624
rect 7764 3568 7820 3624
rect 7849 3568 7905 3624
rect 7934 3568 7990 3624
rect 8019 3568 8075 3624
rect 8104 3568 8160 3624
rect 6996 3482 7052 3538
rect 7082 3482 7138 3538
rect 7168 3482 7224 3538
rect 7254 3482 7310 3538
rect 7339 3482 7395 3538
rect 7424 3482 7480 3538
rect 7509 3482 7565 3538
rect 7594 3482 7650 3538
rect 7679 3482 7735 3538
rect 7764 3482 7820 3538
rect 7849 3482 7905 3538
rect 7934 3482 7990 3538
rect 8019 3482 8075 3538
rect 8104 3482 8160 3538
rect 6996 3396 7052 3452
rect 7082 3396 7138 3452
rect 7168 3396 7224 3452
rect 7254 3396 7310 3452
rect 7339 3396 7395 3452
rect 7424 3396 7480 3452
rect 7509 3396 7565 3452
rect 7594 3396 7650 3452
rect 7679 3396 7735 3452
rect 7764 3396 7820 3452
rect 7849 3396 7905 3452
rect 7934 3396 7990 3452
rect 8019 3396 8075 3452
rect 8104 3396 8160 3452
rect 6996 3310 7052 3366
rect 7082 3310 7138 3366
rect 7168 3310 7224 3366
rect 7254 3310 7310 3366
rect 7339 3310 7395 3366
rect 7424 3310 7480 3366
rect 7509 3310 7565 3366
rect 7594 3310 7650 3366
rect 7679 3310 7735 3366
rect 7764 3310 7820 3366
rect 7849 3310 7905 3366
rect 7934 3310 7990 3366
rect 8019 3310 8075 3366
rect 8104 3310 8160 3366
rect 6996 3224 7052 3280
rect 7082 3224 7138 3280
rect 7168 3224 7224 3280
rect 7254 3224 7310 3280
rect 7339 3224 7395 3280
rect 7424 3224 7480 3280
rect 7509 3224 7565 3280
rect 7594 3224 7650 3280
rect 7679 3224 7735 3280
rect 7764 3224 7820 3280
rect 7849 3224 7905 3280
rect 7934 3224 7990 3280
rect 8019 3224 8075 3280
rect 8104 3224 8160 3280
rect 6996 3138 7052 3194
rect 7082 3138 7138 3194
rect 7168 3138 7224 3194
rect 7254 3138 7310 3194
rect 7339 3138 7395 3194
rect 7424 3138 7480 3194
rect 7509 3138 7565 3194
rect 7594 3138 7650 3194
rect 7679 3138 7735 3194
rect 7764 3138 7820 3194
rect 7849 3138 7905 3194
rect 7934 3138 7990 3194
rect 8019 3138 8075 3194
rect 8104 3138 8160 3194
rect 6996 3052 7052 3108
rect 7082 3052 7138 3108
rect 7168 3052 7224 3108
rect 7254 3052 7310 3108
rect 7339 3052 7395 3108
rect 7424 3052 7480 3108
rect 7509 3052 7565 3108
rect 7594 3052 7650 3108
rect 7679 3052 7735 3108
rect 7764 3052 7820 3108
rect 7849 3052 7905 3108
rect 7934 3052 7990 3108
rect 8019 3052 8075 3108
rect 8104 3052 8160 3108
rect 6996 2966 7052 3022
rect 7082 2966 7138 3022
rect 7168 2966 7224 3022
rect 7254 2966 7310 3022
rect 7339 2966 7395 3022
rect 7424 2966 7480 3022
rect 7509 2966 7565 3022
rect 7594 2966 7650 3022
rect 7679 2966 7735 3022
rect 7764 2966 7820 3022
rect 7849 2966 7905 3022
rect 7934 2966 7990 3022
rect 8019 2966 8075 3022
rect 8104 2966 8160 3022
rect 6996 2880 7052 2936
rect 7082 2880 7138 2936
rect 7168 2880 7224 2936
rect 7254 2880 7310 2936
rect 7339 2880 7395 2936
rect 7424 2880 7480 2936
rect 7509 2880 7565 2936
rect 7594 2880 7650 2936
rect 7679 2880 7735 2936
rect 7764 2880 7820 2936
rect 7849 2880 7905 2936
rect 7934 2880 7990 2936
rect 8019 2880 8075 2936
rect 8104 2880 8160 2936
rect 6996 2794 7052 2850
rect 7082 2794 7138 2850
rect 7168 2794 7224 2850
rect 7254 2794 7310 2850
rect 7339 2794 7395 2850
rect 7424 2794 7480 2850
rect 7509 2794 7565 2850
rect 7594 2794 7650 2850
rect 7679 2794 7735 2850
rect 7764 2794 7820 2850
rect 7849 2794 7905 2850
rect 7934 2794 7990 2850
rect 8019 2794 8075 2850
rect 8104 2794 8160 2850
rect 6996 2708 7052 2764
rect 7082 2708 7138 2764
rect 7168 2708 7224 2764
rect 7254 2708 7310 2764
rect 7339 2708 7395 2764
rect 7424 2708 7480 2764
rect 7509 2708 7565 2764
rect 7594 2708 7650 2764
rect 7679 2708 7735 2764
rect 7764 2708 7820 2764
rect 7849 2708 7905 2764
rect 7934 2708 7990 2764
rect 8019 2708 8075 2764
rect 8104 2708 8160 2764
rect 6996 2622 7052 2678
rect 7082 2622 7138 2678
rect 7168 2622 7224 2678
rect 7254 2622 7310 2678
rect 7339 2622 7395 2678
rect 7424 2622 7480 2678
rect 7509 2622 7565 2678
rect 7594 2622 7650 2678
rect 7679 2622 7735 2678
rect 7764 2622 7820 2678
rect 7849 2622 7905 2678
rect 7934 2622 7990 2678
rect 8019 2622 8075 2678
rect 8104 2622 8160 2678
rect 6996 2536 7052 2592
rect 7082 2536 7138 2592
rect 7168 2536 7224 2592
rect 7254 2536 7310 2592
rect 7339 2536 7395 2592
rect 7424 2536 7480 2592
rect 7509 2536 7565 2592
rect 7594 2536 7650 2592
rect 7679 2536 7735 2592
rect 7764 2536 7820 2592
rect 7849 2536 7905 2592
rect 7934 2536 7990 2592
rect 8019 2536 8075 2592
rect 8104 2536 8160 2592
rect 9176 3567 9232 3623
rect 9262 3567 9318 3623
rect 9348 3567 9404 3623
rect 9434 3567 9490 3623
rect 9520 3567 9576 3623
rect 9606 3567 9662 3623
rect 9692 3567 9748 3623
rect 9778 3567 9834 3623
rect 9864 3567 9920 3623
rect 9950 3567 10006 3623
rect 10036 3567 10092 3623
rect 10122 3567 10178 3623
rect 10208 3567 10264 3623
rect 10294 3567 10350 3623
rect 9176 3481 9232 3537
rect 9262 3481 9318 3537
rect 9348 3481 9404 3537
rect 9434 3481 9490 3537
rect 9520 3481 9576 3537
rect 9606 3481 9662 3537
rect 9692 3481 9748 3537
rect 9778 3481 9834 3537
rect 9864 3481 9920 3537
rect 9950 3481 10006 3537
rect 10036 3481 10092 3537
rect 10122 3481 10178 3537
rect 10208 3481 10264 3537
rect 10294 3481 10350 3537
rect 9176 3395 9232 3451
rect 9262 3395 9318 3451
rect 9348 3395 9404 3451
rect 9434 3395 9490 3451
rect 9520 3395 9576 3451
rect 9606 3395 9662 3451
rect 9692 3395 9748 3451
rect 9778 3395 9834 3451
rect 9864 3395 9920 3451
rect 9950 3395 10006 3451
rect 10036 3395 10092 3451
rect 10122 3395 10178 3451
rect 10208 3395 10264 3451
rect 10294 3395 10350 3451
rect 9176 3309 9232 3365
rect 9262 3309 9318 3365
rect 9348 3309 9404 3365
rect 9434 3309 9490 3365
rect 9520 3309 9576 3365
rect 9606 3309 9662 3365
rect 9692 3309 9748 3365
rect 9778 3309 9834 3365
rect 9864 3309 9920 3365
rect 9950 3309 10006 3365
rect 10036 3309 10092 3365
rect 10122 3309 10178 3365
rect 10208 3309 10264 3365
rect 10294 3309 10350 3365
rect 9176 3223 9232 3279
rect 9262 3223 9318 3279
rect 9348 3223 9404 3279
rect 9434 3223 9490 3279
rect 9520 3223 9576 3279
rect 9606 3223 9662 3279
rect 9692 3223 9748 3279
rect 9778 3223 9834 3279
rect 9864 3223 9920 3279
rect 9950 3223 10006 3279
rect 10036 3223 10092 3279
rect 10122 3223 10178 3279
rect 10208 3223 10264 3279
rect 10294 3223 10350 3279
rect 9176 3137 9232 3193
rect 9262 3137 9318 3193
rect 9348 3137 9404 3193
rect 9434 3137 9490 3193
rect 9520 3137 9576 3193
rect 9606 3137 9662 3193
rect 9692 3137 9748 3193
rect 9778 3137 9834 3193
rect 9864 3137 9920 3193
rect 9950 3137 10006 3193
rect 10036 3137 10092 3193
rect 10122 3137 10178 3193
rect 10208 3137 10264 3193
rect 10294 3137 10350 3193
rect 9176 3051 9232 3107
rect 9262 3051 9318 3107
rect 9348 3051 9404 3107
rect 9434 3051 9490 3107
rect 9520 3051 9576 3107
rect 9606 3051 9662 3107
rect 9692 3051 9748 3107
rect 9778 3051 9834 3107
rect 9864 3051 9920 3107
rect 9950 3051 10006 3107
rect 10036 3051 10092 3107
rect 10122 3051 10178 3107
rect 10208 3051 10264 3107
rect 10294 3051 10350 3107
rect 9176 2965 9232 3021
rect 9262 2965 9318 3021
rect 9348 2965 9404 3021
rect 9434 2965 9490 3021
rect 9520 2965 9576 3021
rect 9606 2965 9662 3021
rect 9692 2965 9748 3021
rect 9778 2965 9834 3021
rect 9864 2965 9920 3021
rect 9950 2965 10006 3021
rect 10036 2965 10092 3021
rect 10122 2965 10178 3021
rect 10208 2965 10264 3021
rect 10294 2965 10350 3021
rect 9176 2879 9232 2935
rect 9262 2879 9318 2935
rect 9348 2879 9404 2935
rect 9434 2879 9490 2935
rect 9520 2879 9576 2935
rect 9606 2879 9662 2935
rect 9692 2879 9748 2935
rect 9778 2879 9834 2935
rect 9864 2879 9920 2935
rect 9950 2879 10006 2935
rect 10036 2879 10092 2935
rect 10122 2879 10178 2935
rect 10208 2879 10264 2935
rect 10294 2879 10350 2935
rect 9176 2793 9232 2849
rect 9262 2793 9318 2849
rect 9348 2793 9404 2849
rect 9434 2793 9490 2849
rect 9520 2793 9576 2849
rect 9606 2793 9662 2849
rect 9692 2793 9748 2849
rect 9778 2793 9834 2849
rect 9864 2793 9920 2849
rect 9950 2793 10006 2849
rect 10036 2793 10092 2849
rect 10122 2793 10178 2849
rect 10208 2793 10264 2849
rect 10294 2793 10350 2849
rect 9176 2707 9232 2763
rect 9262 2707 9318 2763
rect 9348 2707 9404 2763
rect 9434 2707 9490 2763
rect 9520 2707 9576 2763
rect 9606 2707 9662 2763
rect 9692 2707 9748 2763
rect 9778 2707 9834 2763
rect 9864 2707 9920 2763
rect 9950 2707 10006 2763
rect 10036 2707 10092 2763
rect 10122 2707 10178 2763
rect 10208 2707 10264 2763
rect 10294 2707 10350 2763
rect 9176 2621 9232 2677
rect 9262 2621 9318 2677
rect 9348 2621 9404 2677
rect 9434 2621 9490 2677
rect 9520 2621 9576 2677
rect 9606 2621 9662 2677
rect 9692 2621 9748 2677
rect 9778 2621 9834 2677
rect 9864 2621 9920 2677
rect 9950 2621 10006 2677
rect 10036 2621 10092 2677
rect 10122 2621 10178 2677
rect 10208 2621 10264 2677
rect 10294 2621 10350 2677
rect 9176 2535 9232 2591
rect 9262 2535 9318 2591
rect 9348 2535 9404 2591
rect 9434 2535 9490 2591
rect 9520 2535 9576 2591
rect 9606 2535 9662 2591
rect 9692 2535 9748 2591
rect 9778 2535 9834 2591
rect 9864 2535 9920 2591
rect 9950 2535 10006 2591
rect 10036 2535 10092 2591
rect 10122 2535 10178 2591
rect 10208 2535 10264 2591
rect 10294 2535 10350 2591
rect 10668 3567 10724 3623
rect 10749 3567 10805 3623
rect 10829 3567 10885 3623
rect 10909 3567 10965 3623
rect 10989 3567 11045 3623
rect 11069 3567 11125 3623
rect 11149 3567 11205 3623
rect 11229 3567 11285 3623
rect 11309 3567 11365 3623
rect 11389 3567 11445 3623
rect 11469 3567 11525 3623
rect 11549 3567 11605 3623
rect 11629 3567 11685 3623
rect 11709 3567 11765 3623
rect 11789 3567 11845 3623
rect 10668 3481 10724 3537
rect 10749 3481 10805 3537
rect 10829 3481 10885 3537
rect 10909 3481 10965 3537
rect 10989 3481 11045 3537
rect 11069 3481 11125 3537
rect 11149 3481 11205 3537
rect 11229 3481 11285 3537
rect 11309 3481 11365 3537
rect 11389 3481 11445 3537
rect 11469 3481 11525 3537
rect 11549 3481 11605 3537
rect 11629 3481 11685 3537
rect 11709 3481 11765 3537
rect 11789 3481 11845 3537
rect 10668 3395 10724 3451
rect 10749 3395 10805 3451
rect 10829 3395 10885 3451
rect 10909 3395 10965 3451
rect 10989 3395 11045 3451
rect 11069 3395 11125 3451
rect 11149 3395 11205 3451
rect 11229 3395 11285 3451
rect 11309 3395 11365 3451
rect 11389 3395 11445 3451
rect 11469 3395 11525 3451
rect 11549 3395 11605 3451
rect 11629 3395 11685 3451
rect 11709 3395 11765 3451
rect 11789 3395 11845 3451
rect 10668 3309 10724 3365
rect 10749 3309 10805 3365
rect 10829 3309 10885 3365
rect 10909 3309 10965 3365
rect 10989 3309 11045 3365
rect 11069 3309 11125 3365
rect 11149 3309 11205 3365
rect 11229 3309 11285 3365
rect 11309 3309 11365 3365
rect 11389 3309 11445 3365
rect 11469 3309 11525 3365
rect 11549 3309 11605 3365
rect 11629 3309 11685 3365
rect 11709 3309 11765 3365
rect 11789 3309 11845 3365
rect 10668 3223 10724 3279
rect 10749 3223 10805 3279
rect 10829 3223 10885 3279
rect 10909 3223 10965 3279
rect 10989 3223 11045 3279
rect 11069 3223 11125 3279
rect 11149 3223 11205 3279
rect 11229 3223 11285 3279
rect 11309 3223 11365 3279
rect 11389 3223 11445 3279
rect 11469 3223 11525 3279
rect 11549 3223 11605 3279
rect 11629 3223 11685 3279
rect 11709 3223 11765 3279
rect 11789 3223 11845 3279
rect 10668 3137 10724 3193
rect 10749 3137 10805 3193
rect 10829 3137 10885 3193
rect 10909 3137 10965 3193
rect 10989 3137 11045 3193
rect 11069 3137 11125 3193
rect 11149 3137 11205 3193
rect 11229 3137 11285 3193
rect 11309 3137 11365 3193
rect 11389 3137 11445 3193
rect 11469 3137 11525 3193
rect 11549 3137 11605 3193
rect 11629 3137 11685 3193
rect 11709 3137 11765 3193
rect 11789 3137 11845 3193
rect 10668 3051 10724 3107
rect 10749 3051 10805 3107
rect 10829 3051 10885 3107
rect 10909 3051 10965 3107
rect 10989 3051 11045 3107
rect 11069 3051 11125 3107
rect 11149 3051 11205 3107
rect 11229 3051 11285 3107
rect 11309 3051 11365 3107
rect 11389 3051 11445 3107
rect 11469 3051 11525 3107
rect 11549 3051 11605 3107
rect 11629 3051 11685 3107
rect 11709 3051 11765 3107
rect 11789 3051 11845 3107
rect 10668 2965 10724 3021
rect 10749 2965 10805 3021
rect 10829 2965 10885 3021
rect 10909 2965 10965 3021
rect 10989 2965 11045 3021
rect 11069 2965 11125 3021
rect 11149 2965 11205 3021
rect 11229 2965 11285 3021
rect 11309 2965 11365 3021
rect 11389 2965 11445 3021
rect 11469 2965 11525 3021
rect 11549 2965 11605 3021
rect 11629 2965 11685 3021
rect 11709 2965 11765 3021
rect 11789 2965 11845 3021
rect 10668 2879 10724 2935
rect 10749 2879 10805 2935
rect 10829 2879 10885 2935
rect 10909 2879 10965 2935
rect 10989 2879 11045 2935
rect 11069 2879 11125 2935
rect 11149 2879 11205 2935
rect 11229 2879 11285 2935
rect 11309 2879 11365 2935
rect 11389 2879 11445 2935
rect 11469 2879 11525 2935
rect 11549 2879 11605 2935
rect 11629 2879 11685 2935
rect 11709 2879 11765 2935
rect 11789 2879 11845 2935
rect 10668 2793 10724 2849
rect 10749 2793 10805 2849
rect 10829 2793 10885 2849
rect 10909 2793 10965 2849
rect 10989 2793 11045 2849
rect 11069 2793 11125 2849
rect 11149 2793 11205 2849
rect 11229 2793 11285 2849
rect 11309 2793 11365 2849
rect 11389 2793 11445 2849
rect 11469 2793 11525 2849
rect 11549 2793 11605 2849
rect 11629 2793 11685 2849
rect 11709 2793 11765 2849
rect 11789 2793 11845 2849
rect 10668 2707 10724 2763
rect 10749 2707 10805 2763
rect 10829 2707 10885 2763
rect 10909 2707 10965 2763
rect 10989 2707 11045 2763
rect 11069 2707 11125 2763
rect 11149 2707 11205 2763
rect 11229 2707 11285 2763
rect 11309 2707 11365 2763
rect 11389 2707 11445 2763
rect 11469 2707 11525 2763
rect 11549 2707 11605 2763
rect 11629 2707 11685 2763
rect 11709 2707 11765 2763
rect 11789 2707 11845 2763
rect 10668 2621 10724 2677
rect 10749 2621 10805 2677
rect 10829 2621 10885 2677
rect 10909 2621 10965 2677
rect 10989 2621 11045 2677
rect 11069 2621 11125 2677
rect 11149 2621 11205 2677
rect 11229 2621 11285 2677
rect 11309 2621 11365 2677
rect 11389 2621 11445 2677
rect 11469 2621 11525 2677
rect 11549 2621 11605 2677
rect 11629 2621 11685 2677
rect 11709 2621 11765 2677
rect 11789 2621 11845 2677
rect 10668 2535 10724 2591
rect 10749 2535 10805 2591
rect 10829 2535 10885 2591
rect 10909 2535 10965 2591
rect 10989 2535 11045 2591
rect 11069 2535 11125 2591
rect 11149 2535 11205 2591
rect 11229 2535 11285 2591
rect 11309 2535 11365 2591
rect 11389 2535 11445 2591
rect 11469 2535 11525 2591
rect 11549 2535 11605 2591
rect 11629 2535 11685 2591
rect 11709 2535 11765 2591
rect 11789 2535 11845 2591
<< metal3 >>
rect 5376 3624 6571 3631
rect 5376 3568 5385 3624
rect 5441 3568 5471 3624
rect 5527 3568 5557 3624
rect 5613 3568 5643 3624
rect 5699 3568 5728 3624
rect 5784 3568 5813 3624
rect 5869 3568 5898 3624
rect 5954 3568 5983 3624
rect 6039 3568 6068 3624
rect 6124 3568 6153 3624
rect 6209 3568 6238 3624
rect 6294 3568 6323 3624
rect 6379 3568 6408 3624
rect 6464 3568 6493 3624
rect 6549 3568 6571 3624
rect 5376 3538 6571 3568
rect 5376 3482 5385 3538
rect 5441 3482 5471 3538
rect 5527 3482 5557 3538
rect 5613 3482 5643 3538
rect 5699 3482 5728 3538
rect 5784 3482 5813 3538
rect 5869 3482 5898 3538
rect 5954 3482 5983 3538
rect 6039 3482 6068 3538
rect 6124 3482 6153 3538
rect 6209 3482 6238 3538
rect 6294 3482 6323 3538
rect 6379 3482 6408 3538
rect 6464 3482 6493 3538
rect 6549 3482 6571 3538
rect 5376 3452 6571 3482
rect 5376 3396 5385 3452
rect 5441 3396 5471 3452
rect 5527 3396 5557 3452
rect 5613 3396 5643 3452
rect 5699 3396 5728 3452
rect 5784 3396 5813 3452
rect 5869 3396 5898 3452
rect 5954 3396 5983 3452
rect 6039 3396 6068 3452
rect 6124 3396 6153 3452
rect 6209 3396 6238 3452
rect 6294 3396 6323 3452
rect 6379 3396 6408 3452
rect 6464 3396 6493 3452
rect 6549 3396 6571 3452
rect 5376 3366 6571 3396
rect 5376 3310 5385 3366
rect 5441 3310 5471 3366
rect 5527 3310 5557 3366
rect 5613 3310 5643 3366
rect 5699 3310 5728 3366
rect 5784 3310 5813 3366
rect 5869 3310 5898 3366
rect 5954 3310 5983 3366
rect 6039 3310 6068 3366
rect 6124 3310 6153 3366
rect 6209 3310 6238 3366
rect 6294 3310 6323 3366
rect 6379 3310 6408 3366
rect 6464 3310 6493 3366
rect 6549 3310 6571 3366
rect 5376 3280 6571 3310
rect 5376 3224 5385 3280
rect 5441 3224 5471 3280
rect 5527 3224 5557 3280
rect 5613 3224 5643 3280
rect 5699 3224 5728 3280
rect 5784 3224 5813 3280
rect 5869 3224 5898 3280
rect 5954 3224 5983 3280
rect 6039 3224 6068 3280
rect 6124 3224 6153 3280
rect 6209 3224 6238 3280
rect 6294 3224 6323 3280
rect 6379 3224 6408 3280
rect 6464 3224 6493 3280
rect 6549 3224 6571 3280
rect 5376 3194 6571 3224
rect 5376 3138 5385 3194
rect 5441 3138 5471 3194
rect 5527 3138 5557 3194
rect 5613 3138 5643 3194
rect 5699 3138 5728 3194
rect 5784 3138 5813 3194
rect 5869 3138 5898 3194
rect 5954 3138 5983 3194
rect 6039 3138 6068 3194
rect 6124 3138 6153 3194
rect 6209 3138 6238 3194
rect 6294 3138 6323 3194
rect 6379 3138 6408 3194
rect 6464 3138 6493 3194
rect 6549 3138 6571 3194
rect 5376 3108 6571 3138
rect 5376 3052 5385 3108
rect 5441 3052 5471 3108
rect 5527 3052 5557 3108
rect 5613 3052 5643 3108
rect 5699 3052 5728 3108
rect 5784 3052 5813 3108
rect 5869 3052 5898 3108
rect 5954 3052 5983 3108
rect 6039 3052 6068 3108
rect 6124 3052 6153 3108
rect 6209 3052 6238 3108
rect 6294 3052 6323 3108
rect 6379 3052 6408 3108
rect 6464 3052 6493 3108
rect 6549 3052 6571 3108
rect 5376 3022 6571 3052
rect 5376 2966 5385 3022
rect 5441 2966 5471 3022
rect 5527 2966 5557 3022
rect 5613 2966 5643 3022
rect 5699 2966 5728 3022
rect 5784 2966 5813 3022
rect 5869 2966 5898 3022
rect 5954 2966 5983 3022
rect 6039 2966 6068 3022
rect 6124 2966 6153 3022
rect 6209 2966 6238 3022
rect 6294 2966 6323 3022
rect 6379 2966 6408 3022
rect 6464 2966 6493 3022
rect 6549 2966 6571 3022
rect 5376 2936 6571 2966
rect 5376 2880 5385 2936
rect 5441 2880 5471 2936
rect 5527 2880 5557 2936
rect 5613 2880 5643 2936
rect 5699 2880 5728 2936
rect 5784 2880 5813 2936
rect 5869 2880 5898 2936
rect 5954 2880 5983 2936
rect 6039 2880 6068 2936
rect 6124 2880 6153 2936
rect 6209 2880 6238 2936
rect 6294 2880 6323 2936
rect 6379 2880 6408 2936
rect 6464 2880 6493 2936
rect 6549 2880 6571 2936
rect 5376 2850 6571 2880
rect 5376 2794 5385 2850
rect 5441 2794 5471 2850
rect 5527 2794 5557 2850
rect 5613 2794 5643 2850
rect 5699 2794 5728 2850
rect 5784 2794 5813 2850
rect 5869 2794 5898 2850
rect 5954 2794 5983 2850
rect 6039 2794 6068 2850
rect 6124 2794 6153 2850
rect 6209 2794 6238 2850
rect 6294 2794 6323 2850
rect 6379 2794 6408 2850
rect 6464 2794 6493 2850
rect 6549 2794 6571 2850
rect 5376 2764 6571 2794
rect 5376 2708 5385 2764
rect 5441 2708 5471 2764
rect 5527 2708 5557 2764
rect 5613 2708 5643 2764
rect 5699 2708 5728 2764
rect 5784 2708 5813 2764
rect 5869 2708 5898 2764
rect 5954 2708 5983 2764
rect 6039 2708 6068 2764
rect 6124 2708 6153 2764
rect 6209 2708 6238 2764
rect 6294 2708 6323 2764
rect 6379 2708 6408 2764
rect 6464 2708 6493 2764
rect 6549 2708 6571 2764
rect 5376 2678 6571 2708
rect 5376 2622 5385 2678
rect 5441 2622 5471 2678
rect 5527 2622 5557 2678
rect 5613 2622 5643 2678
rect 5699 2622 5728 2678
rect 5784 2622 5813 2678
rect 5869 2622 5898 2678
rect 5954 2622 5983 2678
rect 6039 2622 6068 2678
rect 6124 2622 6153 2678
rect 6209 2622 6238 2678
rect 6294 2622 6323 2678
rect 6379 2622 6408 2678
rect 6464 2622 6493 2678
rect 6549 2622 6571 2678
rect 5376 2592 6571 2622
rect 5376 2536 5385 2592
rect 5441 2536 5471 2592
rect 5527 2536 5557 2592
rect 5613 2536 5643 2592
rect 5699 2536 5728 2592
rect 5784 2536 5813 2592
rect 5869 2536 5898 2592
rect 5954 2536 5983 2592
rect 6039 2536 6068 2592
rect 6124 2536 6153 2592
rect 6209 2536 6238 2592
rect 6294 2536 6323 2592
rect 6379 2536 6408 2592
rect 6464 2536 6493 2592
rect 6549 2536 6571 2592
rect 5376 -205 6571 2536
rect 5376 -269 5403 -205
rect 5467 -269 5485 -205
rect 5549 -269 5567 -205
rect 5631 -269 5649 -205
rect 5713 -269 5731 -205
rect 5795 -269 5813 -205
rect 5877 -269 5895 -205
rect 5959 -269 5976 -205
rect 6040 -269 6057 -205
rect 6121 -269 6138 -205
rect 6202 -269 6219 -205
rect 6283 -269 6300 -205
rect 6364 -269 6381 -205
rect 6445 -269 6462 -205
rect 6526 -269 6571 -205
rect 5376 -285 6571 -269
rect 5376 -349 5403 -285
rect 5467 -349 5485 -285
rect 5549 -349 5567 -285
rect 5631 -349 5649 -285
rect 5713 -349 5731 -285
rect 5795 -349 5813 -285
rect 5877 -349 5895 -285
rect 5959 -349 5976 -285
rect 6040 -349 6057 -285
rect 6121 -349 6138 -285
rect 6202 -349 6219 -285
rect 6283 -349 6300 -285
rect 6364 -349 6381 -285
rect 6445 -349 6462 -285
rect 6526 -349 6571 -285
rect 5376 -365 6571 -349
rect 5376 -429 5403 -365
rect 5467 -429 5485 -365
rect 5549 -429 5567 -365
rect 5631 -429 5649 -365
rect 5713 -429 5731 -365
rect 5795 -429 5813 -365
rect 5877 -429 5895 -365
rect 5959 -429 5976 -365
rect 6040 -429 6057 -365
rect 6121 -429 6138 -365
rect 6202 -429 6219 -365
rect 6283 -429 6300 -365
rect 6364 -429 6381 -365
rect 6445 -429 6462 -365
rect 6526 -429 6571 -365
rect 5376 -445 6571 -429
rect 5376 -509 5403 -445
rect 5467 -509 5485 -445
rect 5549 -509 5567 -445
rect 5631 -509 5649 -445
rect 5713 -509 5731 -445
rect 5795 -509 5813 -445
rect 5877 -509 5895 -445
rect 5959 -509 5976 -445
rect 6040 -509 6057 -445
rect 6121 -509 6138 -445
rect 6202 -509 6219 -445
rect 6283 -509 6300 -445
rect 6364 -509 6381 -445
rect 6445 -509 6462 -445
rect 6526 -509 6571 -445
rect 5376 -525 6571 -509
rect 5376 -589 5403 -525
rect 5467 -589 5485 -525
rect 5549 -589 5567 -525
rect 5631 -589 5649 -525
rect 5713 -589 5731 -525
rect 5795 -589 5813 -525
rect 5877 -589 5895 -525
rect 5959 -589 5976 -525
rect 6040 -589 6057 -525
rect 6121 -589 6138 -525
rect 6202 -589 6219 -525
rect 6283 -589 6300 -525
rect 6364 -589 6381 -525
rect 6445 -589 6462 -525
rect 6526 -589 6571 -525
rect 5376 -605 6571 -589
rect 5376 -669 5403 -605
rect 5467 -669 5485 -605
rect 5549 -669 5567 -605
rect 5631 -669 5649 -605
rect 5713 -669 5731 -605
rect 5795 -669 5813 -605
rect 5877 -669 5895 -605
rect 5959 -669 5976 -605
rect 6040 -669 6057 -605
rect 6121 -669 6138 -605
rect 6202 -669 6219 -605
rect 6283 -669 6300 -605
rect 6364 -669 6381 -605
rect 6445 -669 6462 -605
rect 6526 -669 6571 -605
rect 5376 -685 6571 -669
rect 5376 -749 5403 -685
rect 5467 -749 5485 -685
rect 5549 -749 5567 -685
rect 5631 -749 5649 -685
rect 5713 -749 5731 -685
rect 5795 -749 5813 -685
rect 5877 -749 5895 -685
rect 5959 -749 5976 -685
rect 6040 -749 6057 -685
rect 6121 -749 6138 -685
rect 6202 -749 6219 -685
rect 6283 -749 6300 -685
rect 6364 -749 6381 -685
rect 6445 -749 6462 -685
rect 6526 -749 6571 -685
rect 5376 -765 6571 -749
rect 5376 -829 5403 -765
rect 5467 -829 5485 -765
rect 5549 -829 5567 -765
rect 5631 -829 5649 -765
rect 5713 -829 5731 -765
rect 5795 -829 5813 -765
rect 5877 -829 5895 -765
rect 5959 -829 5976 -765
rect 6040 -829 6057 -765
rect 6121 -829 6138 -765
rect 6202 -829 6219 -765
rect 6283 -829 6300 -765
rect 6364 -829 6381 -765
rect 6445 -829 6462 -765
rect 6526 -829 6571 -765
rect 5376 -845 6571 -829
rect 5376 -909 5403 -845
rect 5467 -909 5485 -845
rect 5549 -909 5567 -845
rect 5631 -909 5649 -845
rect 5713 -909 5731 -845
rect 5795 -909 5813 -845
rect 5877 -909 5895 -845
rect 5959 -909 5976 -845
rect 6040 -909 6057 -845
rect 6121 -909 6138 -845
rect 6202 -909 6219 -845
rect 6283 -909 6300 -845
rect 6364 -909 6381 -845
rect 6445 -909 6462 -845
rect 6526 -909 6571 -845
rect 5376 -925 6571 -909
rect 5376 -989 5403 -925
rect 5467 -989 5485 -925
rect 5549 -989 5567 -925
rect 5631 -989 5649 -925
rect 5713 -989 5731 -925
rect 5795 -989 5813 -925
rect 5877 -989 5895 -925
rect 5959 -989 5976 -925
rect 6040 -989 6057 -925
rect 6121 -989 6138 -925
rect 6202 -989 6219 -925
rect 6283 -989 6300 -925
rect 6364 -989 6381 -925
rect 6445 -989 6462 -925
rect 6526 -989 6571 -925
rect 5376 -991 6571 -989
rect 6987 3624 8182 3631
rect 6987 3568 6996 3624
rect 7052 3568 7082 3624
rect 7138 3568 7168 3624
rect 7224 3568 7254 3624
rect 7310 3568 7339 3624
rect 7395 3568 7424 3624
rect 7480 3568 7509 3624
rect 7565 3568 7594 3624
rect 7650 3568 7679 3624
rect 7735 3568 7764 3624
rect 7820 3568 7849 3624
rect 7905 3568 7934 3624
rect 7990 3568 8019 3624
rect 8075 3568 8104 3624
rect 8160 3568 8182 3624
rect 6987 3538 8182 3568
rect 6987 3482 6996 3538
rect 7052 3482 7082 3538
rect 7138 3482 7168 3538
rect 7224 3482 7254 3538
rect 7310 3482 7339 3538
rect 7395 3482 7424 3538
rect 7480 3482 7509 3538
rect 7565 3482 7594 3538
rect 7650 3482 7679 3538
rect 7735 3482 7764 3538
rect 7820 3482 7849 3538
rect 7905 3482 7934 3538
rect 7990 3482 8019 3538
rect 8075 3482 8104 3538
rect 8160 3482 8182 3538
rect 6987 3452 8182 3482
rect 6987 3396 6996 3452
rect 7052 3396 7082 3452
rect 7138 3396 7168 3452
rect 7224 3396 7254 3452
rect 7310 3396 7339 3452
rect 7395 3396 7424 3452
rect 7480 3396 7509 3452
rect 7565 3396 7594 3452
rect 7650 3396 7679 3452
rect 7735 3396 7764 3452
rect 7820 3396 7849 3452
rect 7905 3396 7934 3452
rect 7990 3396 8019 3452
rect 8075 3396 8104 3452
rect 8160 3396 8182 3452
rect 6987 3366 8182 3396
rect 6987 3310 6996 3366
rect 7052 3310 7082 3366
rect 7138 3310 7168 3366
rect 7224 3310 7254 3366
rect 7310 3310 7339 3366
rect 7395 3310 7424 3366
rect 7480 3310 7509 3366
rect 7565 3310 7594 3366
rect 7650 3310 7679 3366
rect 7735 3310 7764 3366
rect 7820 3310 7849 3366
rect 7905 3310 7934 3366
rect 7990 3310 8019 3366
rect 8075 3310 8104 3366
rect 8160 3310 8182 3366
rect 6987 3280 8182 3310
rect 6987 3224 6996 3280
rect 7052 3224 7082 3280
rect 7138 3224 7168 3280
rect 7224 3224 7254 3280
rect 7310 3224 7339 3280
rect 7395 3224 7424 3280
rect 7480 3224 7509 3280
rect 7565 3224 7594 3280
rect 7650 3224 7679 3280
rect 7735 3224 7764 3280
rect 7820 3224 7849 3280
rect 7905 3224 7934 3280
rect 7990 3224 8019 3280
rect 8075 3224 8104 3280
rect 8160 3224 8182 3280
rect 6987 3194 8182 3224
rect 6987 3138 6996 3194
rect 7052 3138 7082 3194
rect 7138 3138 7168 3194
rect 7224 3138 7254 3194
rect 7310 3138 7339 3194
rect 7395 3138 7424 3194
rect 7480 3138 7509 3194
rect 7565 3138 7594 3194
rect 7650 3138 7679 3194
rect 7735 3138 7764 3194
rect 7820 3138 7849 3194
rect 7905 3138 7934 3194
rect 7990 3138 8019 3194
rect 8075 3138 8104 3194
rect 8160 3138 8182 3194
rect 6987 3108 8182 3138
rect 6987 3052 6996 3108
rect 7052 3052 7082 3108
rect 7138 3052 7168 3108
rect 7224 3052 7254 3108
rect 7310 3052 7339 3108
rect 7395 3052 7424 3108
rect 7480 3052 7509 3108
rect 7565 3052 7594 3108
rect 7650 3052 7679 3108
rect 7735 3052 7764 3108
rect 7820 3052 7849 3108
rect 7905 3052 7934 3108
rect 7990 3052 8019 3108
rect 8075 3052 8104 3108
rect 8160 3052 8182 3108
rect 6987 3022 8182 3052
rect 6987 2966 6996 3022
rect 7052 2966 7082 3022
rect 7138 2966 7168 3022
rect 7224 2966 7254 3022
rect 7310 2966 7339 3022
rect 7395 2966 7424 3022
rect 7480 2966 7509 3022
rect 7565 2966 7594 3022
rect 7650 2966 7679 3022
rect 7735 2966 7764 3022
rect 7820 2966 7849 3022
rect 7905 2966 7934 3022
rect 7990 2966 8019 3022
rect 8075 2966 8104 3022
rect 8160 2966 8182 3022
rect 6987 2936 8182 2966
rect 6987 2880 6996 2936
rect 7052 2880 7082 2936
rect 7138 2880 7168 2936
rect 7224 2880 7254 2936
rect 7310 2880 7339 2936
rect 7395 2880 7424 2936
rect 7480 2880 7509 2936
rect 7565 2880 7594 2936
rect 7650 2880 7679 2936
rect 7735 2880 7764 2936
rect 7820 2880 7849 2936
rect 7905 2880 7934 2936
rect 7990 2880 8019 2936
rect 8075 2880 8104 2936
rect 8160 2880 8182 2936
rect 6987 2850 8182 2880
rect 6987 2794 6996 2850
rect 7052 2794 7082 2850
rect 7138 2794 7168 2850
rect 7224 2794 7254 2850
rect 7310 2794 7339 2850
rect 7395 2794 7424 2850
rect 7480 2794 7509 2850
rect 7565 2794 7594 2850
rect 7650 2794 7679 2850
rect 7735 2794 7764 2850
rect 7820 2794 7849 2850
rect 7905 2794 7934 2850
rect 7990 2794 8019 2850
rect 8075 2794 8104 2850
rect 8160 2794 8182 2850
rect 6987 2764 8182 2794
rect 6987 2708 6996 2764
rect 7052 2708 7082 2764
rect 7138 2708 7168 2764
rect 7224 2708 7254 2764
rect 7310 2708 7339 2764
rect 7395 2708 7424 2764
rect 7480 2708 7509 2764
rect 7565 2708 7594 2764
rect 7650 2708 7679 2764
rect 7735 2708 7764 2764
rect 7820 2708 7849 2764
rect 7905 2708 7934 2764
rect 7990 2708 8019 2764
rect 8075 2708 8104 2764
rect 8160 2708 8182 2764
rect 6987 2678 8182 2708
rect 6987 2622 6996 2678
rect 7052 2622 7082 2678
rect 7138 2622 7168 2678
rect 7224 2622 7254 2678
rect 7310 2622 7339 2678
rect 7395 2622 7424 2678
rect 7480 2622 7509 2678
rect 7565 2622 7594 2678
rect 7650 2622 7679 2678
rect 7735 2622 7764 2678
rect 7820 2622 7849 2678
rect 7905 2622 7934 2678
rect 7990 2622 8019 2678
rect 8075 2622 8104 2678
rect 8160 2622 8182 2678
rect 6987 2592 8182 2622
rect 6987 2536 6996 2592
rect 7052 2536 7082 2592
rect 7138 2536 7168 2592
rect 7224 2536 7254 2592
rect 7310 2536 7339 2592
rect 7395 2536 7424 2592
rect 7480 2536 7509 2592
rect 7565 2536 7594 2592
rect 7650 2536 7679 2592
rect 7735 2536 7764 2592
rect 7820 2536 7849 2592
rect 7905 2536 7934 2592
rect 7990 2536 8019 2592
rect 8075 2536 8104 2592
rect 8160 2536 8182 2592
rect 6987 -205 8182 2536
rect 6987 -269 7014 -205
rect 7078 -269 7096 -205
rect 7160 -269 7178 -205
rect 7242 -269 7260 -205
rect 7324 -269 7342 -205
rect 7406 -269 7424 -205
rect 7488 -269 7506 -205
rect 7570 -269 7587 -205
rect 7651 -269 7668 -205
rect 7732 -269 7749 -205
rect 7813 -269 7830 -205
rect 7894 -269 7911 -205
rect 7975 -269 7992 -205
rect 8056 -269 8073 -205
rect 8137 -269 8182 -205
rect 6987 -285 8182 -269
rect 6987 -349 7014 -285
rect 7078 -349 7096 -285
rect 7160 -349 7178 -285
rect 7242 -349 7260 -285
rect 7324 -349 7342 -285
rect 7406 -349 7424 -285
rect 7488 -349 7506 -285
rect 7570 -349 7587 -285
rect 7651 -349 7668 -285
rect 7732 -349 7749 -285
rect 7813 -349 7830 -285
rect 7894 -349 7911 -285
rect 7975 -349 7992 -285
rect 8056 -349 8073 -285
rect 8137 -349 8182 -285
rect 9164 3623 10359 3631
rect 9164 3567 9176 3623
rect 9232 3567 9262 3623
rect 9318 3567 9348 3623
rect 9404 3567 9434 3623
rect 9490 3567 9520 3623
rect 9576 3567 9606 3623
rect 9662 3567 9692 3623
rect 9748 3567 9778 3623
rect 9834 3567 9864 3623
rect 9920 3567 9950 3623
rect 10006 3567 10036 3623
rect 10092 3567 10122 3623
rect 10178 3567 10208 3623
rect 10264 3567 10294 3623
rect 10350 3567 10359 3623
rect 9164 3537 10359 3567
rect 9164 3481 9176 3537
rect 9232 3481 9262 3537
rect 9318 3481 9348 3537
rect 9404 3481 9434 3537
rect 9490 3481 9520 3537
rect 9576 3481 9606 3537
rect 9662 3481 9692 3537
rect 9748 3481 9778 3537
rect 9834 3481 9864 3537
rect 9920 3481 9950 3537
rect 10006 3481 10036 3537
rect 10092 3481 10122 3537
rect 10178 3481 10208 3537
rect 10264 3481 10294 3537
rect 10350 3481 10359 3537
rect 9164 3451 10359 3481
rect 9164 3395 9176 3451
rect 9232 3395 9262 3451
rect 9318 3395 9348 3451
rect 9404 3395 9434 3451
rect 9490 3395 9520 3451
rect 9576 3395 9606 3451
rect 9662 3395 9692 3451
rect 9748 3395 9778 3451
rect 9834 3395 9864 3451
rect 9920 3395 9950 3451
rect 10006 3395 10036 3451
rect 10092 3395 10122 3451
rect 10178 3395 10208 3451
rect 10264 3395 10294 3451
rect 10350 3395 10359 3451
rect 9164 3365 10359 3395
rect 9164 3309 9176 3365
rect 9232 3309 9262 3365
rect 9318 3309 9348 3365
rect 9404 3309 9434 3365
rect 9490 3309 9520 3365
rect 9576 3309 9606 3365
rect 9662 3309 9692 3365
rect 9748 3309 9778 3365
rect 9834 3309 9864 3365
rect 9920 3309 9950 3365
rect 10006 3309 10036 3365
rect 10092 3309 10122 3365
rect 10178 3309 10208 3365
rect 10264 3309 10294 3365
rect 10350 3309 10359 3365
rect 9164 3279 10359 3309
rect 9164 3223 9176 3279
rect 9232 3223 9262 3279
rect 9318 3223 9348 3279
rect 9404 3223 9434 3279
rect 9490 3223 9520 3279
rect 9576 3223 9606 3279
rect 9662 3223 9692 3279
rect 9748 3223 9778 3279
rect 9834 3223 9864 3279
rect 9920 3223 9950 3279
rect 10006 3223 10036 3279
rect 10092 3223 10122 3279
rect 10178 3223 10208 3279
rect 10264 3223 10294 3279
rect 10350 3223 10359 3279
rect 9164 3193 10359 3223
rect 9164 3137 9176 3193
rect 9232 3137 9262 3193
rect 9318 3137 9348 3193
rect 9404 3137 9434 3193
rect 9490 3137 9520 3193
rect 9576 3137 9606 3193
rect 9662 3137 9692 3193
rect 9748 3137 9778 3193
rect 9834 3137 9864 3193
rect 9920 3137 9950 3193
rect 10006 3137 10036 3193
rect 10092 3137 10122 3193
rect 10178 3137 10208 3193
rect 10264 3137 10294 3193
rect 10350 3137 10359 3193
rect 9164 3107 10359 3137
rect 9164 3051 9176 3107
rect 9232 3051 9262 3107
rect 9318 3051 9348 3107
rect 9404 3051 9434 3107
rect 9490 3051 9520 3107
rect 9576 3051 9606 3107
rect 9662 3051 9692 3107
rect 9748 3051 9778 3107
rect 9834 3051 9864 3107
rect 9920 3051 9950 3107
rect 10006 3051 10036 3107
rect 10092 3051 10122 3107
rect 10178 3051 10208 3107
rect 10264 3051 10294 3107
rect 10350 3051 10359 3107
rect 9164 3021 10359 3051
rect 9164 2965 9176 3021
rect 9232 2965 9262 3021
rect 9318 2965 9348 3021
rect 9404 2965 9434 3021
rect 9490 2965 9520 3021
rect 9576 2965 9606 3021
rect 9662 2965 9692 3021
rect 9748 2965 9778 3021
rect 9834 2965 9864 3021
rect 9920 2965 9950 3021
rect 10006 2965 10036 3021
rect 10092 2965 10122 3021
rect 10178 2965 10208 3021
rect 10264 2965 10294 3021
rect 10350 2965 10359 3021
rect 9164 2935 10359 2965
rect 9164 2879 9176 2935
rect 9232 2879 9262 2935
rect 9318 2879 9348 2935
rect 9404 2879 9434 2935
rect 9490 2879 9520 2935
rect 9576 2879 9606 2935
rect 9662 2879 9692 2935
rect 9748 2879 9778 2935
rect 9834 2879 9864 2935
rect 9920 2879 9950 2935
rect 10006 2879 10036 2935
rect 10092 2879 10122 2935
rect 10178 2879 10208 2935
rect 10264 2879 10294 2935
rect 10350 2879 10359 2935
rect 9164 2849 10359 2879
rect 9164 2793 9176 2849
rect 9232 2793 9262 2849
rect 9318 2793 9348 2849
rect 9404 2793 9434 2849
rect 9490 2793 9520 2849
rect 9576 2793 9606 2849
rect 9662 2793 9692 2849
rect 9748 2793 9778 2849
rect 9834 2793 9864 2849
rect 9920 2793 9950 2849
rect 10006 2793 10036 2849
rect 10092 2793 10122 2849
rect 10178 2793 10208 2849
rect 10264 2793 10294 2849
rect 10350 2793 10359 2849
rect 9164 2763 10359 2793
rect 9164 2707 9176 2763
rect 9232 2707 9262 2763
rect 9318 2707 9348 2763
rect 9404 2707 9434 2763
rect 9490 2707 9520 2763
rect 9576 2707 9606 2763
rect 9662 2707 9692 2763
rect 9748 2707 9778 2763
rect 9834 2707 9864 2763
rect 9920 2707 9950 2763
rect 10006 2707 10036 2763
rect 10092 2707 10122 2763
rect 10178 2707 10208 2763
rect 10264 2707 10294 2763
rect 10350 2707 10359 2763
rect 9164 2677 10359 2707
rect 9164 2621 9176 2677
rect 9232 2621 9262 2677
rect 9318 2621 9348 2677
rect 9404 2621 9434 2677
rect 9490 2621 9520 2677
rect 9576 2621 9606 2677
rect 9662 2621 9692 2677
rect 9748 2621 9778 2677
rect 9834 2621 9864 2677
rect 9920 2621 9950 2677
rect 10006 2621 10036 2677
rect 10092 2621 10122 2677
rect 10178 2621 10208 2677
rect 10264 2621 10294 2677
rect 10350 2621 10359 2677
rect 9164 2591 10359 2621
rect 9164 2535 9176 2591
rect 9232 2535 9262 2591
rect 9318 2535 9348 2591
rect 9404 2535 9434 2591
rect 9490 2535 9520 2591
rect 9576 2535 9606 2591
rect 9662 2535 9692 2591
rect 9748 2535 9778 2591
rect 9834 2535 9864 2591
rect 9920 2535 9950 2591
rect 10006 2535 10036 2591
rect 10092 2535 10122 2591
rect 10178 2535 10208 2591
rect 10264 2535 10294 2591
rect 10350 2535 10359 2591
rect 9164 -28 10359 2535
rect 10659 3623 11854 3631
rect 10659 3567 10668 3623
rect 10724 3567 10749 3623
rect 10805 3567 10829 3623
rect 10885 3567 10909 3623
rect 10965 3567 10989 3623
rect 11045 3567 11069 3623
rect 11125 3567 11149 3623
rect 11205 3567 11229 3623
rect 11285 3567 11309 3623
rect 11365 3567 11389 3623
rect 11445 3567 11469 3623
rect 11525 3567 11549 3623
rect 11605 3567 11629 3623
rect 11685 3567 11709 3623
rect 11765 3567 11789 3623
rect 11845 3567 11854 3623
rect 10659 3537 11854 3567
rect 10659 3481 10668 3537
rect 10724 3481 10749 3537
rect 10805 3481 10829 3537
rect 10885 3481 10909 3537
rect 10965 3481 10989 3537
rect 11045 3481 11069 3537
rect 11125 3481 11149 3537
rect 11205 3481 11229 3537
rect 11285 3481 11309 3537
rect 11365 3481 11389 3537
rect 11445 3481 11469 3537
rect 11525 3481 11549 3537
rect 11605 3481 11629 3537
rect 11685 3481 11709 3537
rect 11765 3481 11789 3537
rect 11845 3481 11854 3537
rect 10659 3451 11854 3481
rect 10659 3395 10668 3451
rect 10724 3395 10749 3451
rect 10805 3395 10829 3451
rect 10885 3395 10909 3451
rect 10965 3395 10989 3451
rect 11045 3395 11069 3451
rect 11125 3395 11149 3451
rect 11205 3395 11229 3451
rect 11285 3395 11309 3451
rect 11365 3395 11389 3451
rect 11445 3395 11469 3451
rect 11525 3395 11549 3451
rect 11605 3395 11629 3451
rect 11685 3395 11709 3451
rect 11765 3395 11789 3451
rect 11845 3395 11854 3451
rect 10659 3365 11854 3395
rect 10659 3309 10668 3365
rect 10724 3309 10749 3365
rect 10805 3309 10829 3365
rect 10885 3309 10909 3365
rect 10965 3309 10989 3365
rect 11045 3309 11069 3365
rect 11125 3309 11149 3365
rect 11205 3309 11229 3365
rect 11285 3309 11309 3365
rect 11365 3309 11389 3365
rect 11445 3309 11469 3365
rect 11525 3309 11549 3365
rect 11605 3309 11629 3365
rect 11685 3309 11709 3365
rect 11765 3309 11789 3365
rect 11845 3309 11854 3365
rect 10659 3279 11854 3309
rect 10659 3223 10668 3279
rect 10724 3223 10749 3279
rect 10805 3223 10829 3279
rect 10885 3223 10909 3279
rect 10965 3223 10989 3279
rect 11045 3223 11069 3279
rect 11125 3223 11149 3279
rect 11205 3223 11229 3279
rect 11285 3223 11309 3279
rect 11365 3223 11389 3279
rect 11445 3223 11469 3279
rect 11525 3223 11549 3279
rect 11605 3223 11629 3279
rect 11685 3223 11709 3279
rect 11765 3223 11789 3279
rect 11845 3223 11854 3279
rect 10659 3193 11854 3223
rect 10659 3137 10668 3193
rect 10724 3137 10749 3193
rect 10805 3137 10829 3193
rect 10885 3137 10909 3193
rect 10965 3137 10989 3193
rect 11045 3137 11069 3193
rect 11125 3137 11149 3193
rect 11205 3137 11229 3193
rect 11285 3137 11309 3193
rect 11365 3137 11389 3193
rect 11445 3137 11469 3193
rect 11525 3137 11549 3193
rect 11605 3137 11629 3193
rect 11685 3137 11709 3193
rect 11765 3137 11789 3193
rect 11845 3137 11854 3193
rect 10659 3107 11854 3137
rect 10659 3051 10668 3107
rect 10724 3051 10749 3107
rect 10805 3051 10829 3107
rect 10885 3051 10909 3107
rect 10965 3051 10989 3107
rect 11045 3051 11069 3107
rect 11125 3051 11149 3107
rect 11205 3051 11229 3107
rect 11285 3051 11309 3107
rect 11365 3051 11389 3107
rect 11445 3051 11469 3107
rect 11525 3051 11549 3107
rect 11605 3051 11629 3107
rect 11685 3051 11709 3107
rect 11765 3051 11789 3107
rect 11845 3051 11854 3107
rect 10659 3021 11854 3051
rect 10659 2965 10668 3021
rect 10724 2965 10749 3021
rect 10805 2965 10829 3021
rect 10885 2965 10909 3021
rect 10965 2965 10989 3021
rect 11045 2965 11069 3021
rect 11125 2965 11149 3021
rect 11205 2965 11229 3021
rect 11285 2965 11309 3021
rect 11365 2965 11389 3021
rect 11445 2965 11469 3021
rect 11525 2965 11549 3021
rect 11605 2965 11629 3021
rect 11685 2965 11709 3021
rect 11765 2965 11789 3021
rect 11845 2965 11854 3021
rect 10659 2935 11854 2965
rect 10659 2879 10668 2935
rect 10724 2879 10749 2935
rect 10805 2879 10829 2935
rect 10885 2879 10909 2935
rect 10965 2879 10989 2935
rect 11045 2879 11069 2935
rect 11125 2879 11149 2935
rect 11205 2879 11229 2935
rect 11285 2879 11309 2935
rect 11365 2879 11389 2935
rect 11445 2879 11469 2935
rect 11525 2879 11549 2935
rect 11605 2879 11629 2935
rect 11685 2879 11709 2935
rect 11765 2879 11789 2935
rect 11845 2879 11854 2935
rect 10659 2849 11854 2879
rect 10659 2793 10668 2849
rect 10724 2793 10749 2849
rect 10805 2793 10829 2849
rect 10885 2793 10909 2849
rect 10965 2793 10989 2849
rect 11045 2793 11069 2849
rect 11125 2793 11149 2849
rect 11205 2793 11229 2849
rect 11285 2793 11309 2849
rect 11365 2793 11389 2849
rect 11445 2793 11469 2849
rect 11525 2793 11549 2849
rect 11605 2793 11629 2849
rect 11685 2793 11709 2849
rect 11765 2793 11789 2849
rect 11845 2793 11854 2849
rect 10659 2763 11854 2793
rect 10659 2707 10668 2763
rect 10724 2707 10749 2763
rect 10805 2707 10829 2763
rect 10885 2707 10909 2763
rect 10965 2707 10989 2763
rect 11045 2707 11069 2763
rect 11125 2707 11149 2763
rect 11205 2707 11229 2763
rect 11285 2707 11309 2763
rect 11365 2707 11389 2763
rect 11445 2707 11469 2763
rect 11525 2707 11549 2763
rect 11605 2707 11629 2763
rect 11685 2707 11709 2763
rect 11765 2707 11789 2763
rect 11845 2707 11854 2763
rect 10659 2677 11854 2707
rect 10659 2621 10668 2677
rect 10724 2621 10749 2677
rect 10805 2621 10829 2677
rect 10885 2621 10909 2677
rect 10965 2621 10989 2677
rect 11045 2621 11069 2677
rect 11125 2621 11149 2677
rect 11205 2621 11229 2677
rect 11285 2621 11309 2677
rect 11365 2621 11389 2677
rect 11445 2621 11469 2677
rect 11525 2621 11549 2677
rect 11605 2621 11629 2677
rect 11685 2621 11709 2677
rect 11765 2621 11789 2677
rect 11845 2621 11854 2677
rect 10659 2591 11854 2621
rect 10659 2535 10668 2591
rect 10724 2535 10749 2591
rect 10805 2535 10829 2591
rect 10885 2535 10909 2591
rect 10965 2535 10989 2591
rect 11045 2535 11069 2591
rect 11125 2535 11149 2591
rect 11205 2535 11229 2591
rect 11285 2535 11309 2591
rect 11365 2535 11389 2591
rect 11445 2535 11469 2591
rect 11525 2535 11549 2591
rect 11605 2535 11629 2591
rect 11685 2535 11709 2591
rect 11765 2535 11789 2591
rect 11845 2535 11854 2591
rect 10659 321 11854 2535
tri 10659 193 10787 321 ne
rect 10787 193 11854 321
tri 10359 -28 10580 193 sw
tri 10787 -28 11008 193 ne
rect 11008 -28 11854 193
tri 11854 -28 12698 816 sw
rect 9164 -198 10580 -28
tri 10580 -198 10750 -28 sw
tri 11008 -198 11178 -28 ne
rect 11178 -198 12698 -28
rect 9164 -203 10750 -198
tri 10750 -203 10755 -198 sw
tri 11178 -203 11183 -198 ne
rect 11183 -203 12698 -198
rect 9164 -204 10755 -203
rect 9164 -260 9528 -204
rect 9164 -302 9194 -260
tri 9164 -330 9192 -302 ne
rect 9192 -324 9194 -302
rect 9258 -324 9304 -260
rect 9368 -324 9414 -260
rect 9478 -268 9528 -260
rect 9592 -268 9609 -204
rect 9673 -268 9690 -204
rect 9754 -268 9770 -204
rect 9834 -268 9850 -204
rect 9914 -268 9930 -204
rect 9994 -268 10010 -204
rect 10074 -268 10090 -204
rect 10154 -268 10170 -204
rect 10234 -268 10250 -204
rect 10314 -268 10330 -204
rect 10394 -268 10410 -204
rect 10474 -268 10490 -204
rect 10554 -223 10755 -204
tri 10755 -223 10775 -203 sw
tri 11183 -223 11203 -203 ne
rect 11203 -218 12698 -203
rect 11203 -223 11507 -218
rect 10554 -268 10775 -223
rect 9478 -298 10775 -268
rect 9478 -324 9528 -298
rect 9192 -330 9528 -324
rect 6987 -365 8182 -349
rect 6987 -429 7014 -365
rect 7078 -429 7096 -365
rect 7160 -429 7178 -365
rect 7242 -429 7260 -365
rect 7324 -429 7342 -365
rect 7406 -429 7424 -365
rect 7488 -429 7506 -365
rect 7570 -429 7587 -365
rect 7651 -429 7668 -365
rect 7732 -429 7749 -365
rect 7813 -429 7830 -365
rect 7894 -429 7911 -365
rect 7975 -429 7992 -365
rect 8056 -429 8073 -365
rect 8137 -429 8182 -365
rect 6987 -445 8182 -429
rect 6987 -509 7014 -445
rect 7078 -509 7096 -445
rect 7160 -509 7178 -445
rect 7242 -509 7260 -445
rect 7324 -509 7342 -445
rect 7406 -509 7424 -445
rect 7488 -509 7506 -445
rect 7570 -509 7587 -445
rect 7651 -509 7668 -445
rect 7732 -509 7749 -445
rect 7813 -509 7830 -445
rect 7894 -509 7911 -445
rect 7975 -509 7992 -445
rect 8056 -509 8073 -445
rect 8137 -509 8182 -445
rect 6987 -525 8182 -509
rect 6987 -589 7014 -525
rect 7078 -589 7096 -525
rect 7160 -589 7178 -525
rect 7242 -589 7260 -525
rect 7324 -589 7342 -525
rect 7406 -589 7424 -525
rect 7488 -589 7506 -525
rect 7570 -589 7587 -525
rect 7651 -589 7668 -525
rect 7732 -589 7749 -525
rect 7813 -589 7830 -525
rect 7894 -589 7911 -525
rect 7975 -589 7992 -525
rect 8056 -589 8073 -525
rect 8137 -589 8182 -525
rect 6987 -605 8182 -589
rect 6987 -669 7014 -605
rect 7078 -669 7096 -605
rect 7160 -669 7178 -605
rect 7242 -669 7260 -605
rect 7324 -669 7342 -605
rect 7406 -669 7424 -605
rect 7488 -669 7506 -605
rect 7570 -669 7587 -605
rect 7651 -669 7668 -605
rect 7732 -669 7749 -605
rect 7813 -669 7830 -605
rect 7894 -669 7911 -605
rect 7975 -669 7992 -605
rect 8056 -669 8073 -605
rect 8137 -669 8182 -605
tri 9192 -645 9507 -330 ne
rect 9507 -362 9528 -330
rect 9592 -362 9609 -298
rect 9673 -362 9690 -298
rect 9754 -362 9770 -298
rect 9834 -362 9850 -298
rect 9914 -362 9930 -298
rect 9994 -362 10010 -298
rect 10074 -362 10090 -298
rect 10154 -362 10170 -298
rect 10234 -362 10250 -298
rect 10314 -362 10330 -298
rect 10394 -362 10410 -298
rect 10474 -362 10490 -298
rect 10554 -328 10775 -298
tri 10775 -328 10880 -223 sw
tri 11203 -328 11308 -223 ne
rect 11308 -328 11507 -223
rect 10554 -334 10880 -328
rect 10554 -362 10585 -334
rect 9507 -392 10585 -362
rect 9507 -456 9528 -392
rect 9592 -456 9609 -392
rect 9673 -456 9690 -392
rect 9754 -456 9770 -392
rect 9834 -456 9850 -392
rect 9914 -456 9930 -392
rect 9994 -456 10010 -392
rect 10074 -456 10090 -392
rect 10154 -456 10170 -392
rect 10234 -456 10250 -392
rect 10314 -456 10330 -392
rect 10394 -456 10410 -392
rect 10474 -456 10490 -392
rect 10554 -398 10585 -392
rect 10649 -398 10695 -334
rect 10759 -398 10805 -334
rect 10869 -398 10880 -334
rect 10554 -416 10880 -398
rect 10554 -456 10585 -416
rect 9507 -480 10585 -456
rect 10649 -480 10695 -416
rect 10759 -480 10805 -416
rect 10869 -480 10880 -416
rect 9507 -486 10880 -480
rect 9507 -550 9528 -486
rect 9592 -550 9609 -486
rect 9673 -550 9690 -486
rect 9754 -550 9770 -486
rect 9834 -550 9850 -486
rect 9914 -550 9930 -486
rect 9994 -550 10010 -486
rect 10074 -550 10090 -486
rect 10154 -550 10170 -486
rect 10234 -550 10250 -486
rect 10314 -550 10330 -486
rect 10394 -550 10410 -486
rect 10474 -550 10490 -486
rect 10554 -498 10880 -486
rect 10554 -550 10585 -498
rect 9507 -562 10585 -550
rect 10649 -562 10695 -498
rect 10759 -562 10805 -498
rect 10869 -524 10880 -498
tri 10880 -524 11076 -328 sw
tri 11308 -524 11504 -328 ne
rect 11504 -442 11507 -328
rect 12691 -442 12698 -218
rect 11504 -459 12698 -442
rect 11504 -523 11507 -459
rect 11571 -523 11587 -459
rect 11651 -523 11667 -459
rect 11731 -523 11747 -459
rect 11811 -523 11827 -459
rect 11891 -523 11907 -459
rect 11971 -523 11987 -459
rect 12051 -523 12067 -459
rect 12131 -523 12147 -459
rect 12211 -523 12227 -459
rect 12291 -523 12307 -459
rect 12371 -523 12387 -459
rect 12451 -523 12467 -459
rect 12531 -523 12547 -459
rect 12611 -523 12627 -459
rect 12691 -523 12698 -459
rect 10869 -562 11076 -524
rect 9507 -580 11076 -562
rect 9507 -644 9528 -580
rect 9592 -644 9609 -580
rect 9673 -644 9690 -580
rect 9754 -644 9770 -580
rect 9834 -644 9850 -580
rect 9914 -644 9930 -580
rect 9994 -644 10010 -580
rect 10074 -644 10090 -580
rect 10154 -644 10170 -580
rect 10234 -644 10250 -580
rect 10314 -644 10330 -580
rect 10394 -644 10410 -580
rect 10474 -644 10490 -580
rect 10554 -644 10585 -580
rect 10649 -644 10695 -580
rect 10759 -644 10805 -580
rect 10869 -644 11076 -580
rect 9507 -645 11076 -644
tri 9507 -651 9513 -645 ne
rect 9513 -650 11076 -645
tri 11076 -650 11202 -524 sw
rect 11504 -540 12698 -523
rect 11504 -604 11507 -540
rect 11571 -604 11587 -540
rect 11651 -604 11667 -540
rect 11731 -604 11747 -540
rect 11811 -604 11827 -540
rect 11891 -604 11907 -540
rect 11971 -604 11987 -540
rect 12051 -604 12067 -540
rect 12131 -604 12147 -540
rect 12211 -604 12227 -540
rect 12291 -604 12307 -540
rect 12371 -604 12387 -540
rect 12451 -604 12467 -540
rect 12531 -604 12547 -540
rect 12611 -604 12627 -540
rect 12691 -604 12698 -540
rect 11504 -621 12698 -604
rect 9513 -651 11202 -650
tri 11202 -651 11203 -650 sw
rect 6987 -685 8182 -669
tri 9513 -673 9535 -651 ne
rect 9535 -673 11203 -651
rect 6987 -749 7014 -685
rect 7078 -749 7096 -685
rect 7160 -749 7178 -685
rect 7242 -749 7260 -685
rect 7324 -749 7342 -685
rect 7406 -749 7424 -685
rect 7488 -749 7506 -685
rect 7570 -749 7587 -685
rect 7651 -749 7668 -685
rect 7732 -749 7749 -685
rect 7813 -749 7830 -685
rect 7894 -749 7911 -685
rect 7975 -749 7992 -685
rect 8056 -749 8073 -685
rect 8137 -749 8182 -685
rect 6987 -765 8182 -749
rect 6987 -829 7014 -765
rect 7078 -829 7096 -765
rect 7160 -829 7178 -765
rect 7242 -829 7260 -765
rect 7324 -829 7342 -765
rect 7406 -829 7424 -765
rect 7488 -829 7506 -765
rect 7570 -829 7587 -765
rect 7651 -829 7668 -765
rect 7732 -829 7749 -765
rect 7813 -829 7830 -765
rect 7894 -829 7911 -765
rect 7975 -829 7992 -765
rect 8056 -829 8073 -765
rect 8137 -829 8182 -765
rect 6987 -845 8182 -829
rect 6987 -909 7014 -845
rect 7078 -909 7096 -845
rect 7160 -909 7178 -845
rect 7242 -909 7260 -845
rect 7324 -909 7342 -845
rect 7406 -909 7424 -845
rect 7488 -909 7506 -845
rect 7570 -909 7587 -845
rect 7651 -909 7668 -845
rect 7732 -909 7749 -845
rect 7813 -909 7830 -845
rect 7894 -909 7911 -845
rect 7975 -909 7992 -845
rect 8056 -909 8073 -845
rect 8137 -909 8182 -845
tri 9535 -886 9748 -673 ne
rect 9748 -679 11203 -673
rect 9748 -743 9771 -679
rect 9835 -743 9905 -679
rect 9969 -743 10016 -679
rect 9748 -816 10016 -743
rect 9748 -880 9771 -816
rect 9835 -880 9905 -816
rect 9969 -880 10016 -816
rect 9748 -886 10016 -880
rect 6987 -925 8182 -909
rect 6987 -989 7014 -925
rect 7078 -989 7096 -925
rect 7160 -989 7178 -925
rect 7242 -989 7260 -925
rect 7324 -989 7342 -925
rect 7406 -989 7424 -925
rect 7488 -989 7506 -925
rect 7570 -989 7587 -925
rect 7651 -989 7668 -925
rect 7732 -989 7749 -925
rect 7813 -989 7830 -925
rect 7894 -989 7911 -925
rect 7975 -989 7992 -925
rect 8056 -989 8073 -925
rect 8137 -989 8182 -925
rect 6987 -991 8182 -989
tri 9748 -991 9853 -886 ne
rect 9853 -903 10016 -886
rect 11200 -903 11203 -679
rect 9853 -920 11203 -903
rect 9853 -984 10016 -920
rect 10080 -984 10096 -920
rect 10160 -984 10176 -920
rect 10240 -984 10256 -920
rect 10320 -984 10336 -920
rect 10400 -984 10416 -920
rect 10480 -984 10496 -920
rect 10560 -984 10576 -920
rect 10640 -984 10656 -920
rect 10720 -984 10736 -920
rect 10800 -984 10816 -920
rect 10880 -984 10896 -920
rect 10960 -984 10976 -920
rect 11040 -984 11056 -920
rect 11120 -984 11136 -920
rect 11200 -984 11203 -920
rect 9853 -991 11203 -984
tri 9853 -1152 10014 -991 ne
rect 10014 -1001 11203 -991
rect 10014 -1065 10016 -1001
rect 10080 -1065 10096 -1001
rect 10160 -1065 10176 -1001
rect 10240 -1065 10256 -1001
rect 10320 -1065 10336 -1001
rect 10400 -1065 10416 -1001
rect 10480 -1065 10496 -1001
rect 10560 -1065 10576 -1001
rect 10640 -1065 10656 -1001
rect 10720 -1065 10736 -1001
rect 10800 -1065 10816 -1001
rect 10880 -1065 10896 -1001
rect 10960 -1065 10976 -1001
rect 11040 -1065 11056 -1001
rect 11120 -1065 11136 -1001
rect 11200 -1065 11203 -1001
rect 10014 -1082 11203 -1065
rect 10014 -1146 10016 -1082
rect 10080 -1146 10096 -1082
rect 10160 -1146 10176 -1082
rect 10240 -1146 10256 -1082
rect 10320 -1146 10336 -1082
rect 10400 -1146 10416 -1082
rect 10480 -1146 10496 -1082
rect 10560 -1146 10576 -1082
rect 10640 -1146 10656 -1082
rect 10720 -1146 10736 -1082
rect 10800 -1146 10816 -1082
rect 10880 -1146 10896 -1082
rect 10960 -1146 10976 -1082
rect 11040 -1146 11056 -1082
rect 11120 -1146 11136 -1082
rect 11200 -1146 11203 -1082
rect 10014 -1163 11203 -1146
rect 10014 -1227 10016 -1163
rect 10080 -1227 10096 -1163
rect 10160 -1227 10176 -1163
rect 10240 -1227 10256 -1163
rect 10320 -1227 10336 -1163
rect 10400 -1227 10416 -1163
rect 10480 -1227 10496 -1163
rect 10560 -1227 10576 -1163
rect 10640 -1227 10656 -1163
rect 10720 -1227 10736 -1163
rect 10800 -1227 10816 -1163
rect 10880 -1227 10896 -1163
rect 10960 -1227 10976 -1163
rect 11040 -1227 11056 -1163
rect 11120 -1227 11136 -1163
rect 11200 -1227 11203 -1163
rect 10014 -1244 11203 -1227
rect 10014 -1308 10016 -1244
rect 10080 -1308 10096 -1244
rect 10160 -1308 10176 -1244
rect 10240 -1308 10256 -1244
rect 10320 -1308 10336 -1244
rect 10400 -1308 10416 -1244
rect 10480 -1308 10496 -1244
rect 10560 -1308 10576 -1244
rect 10640 -1308 10656 -1244
rect 10720 -1308 10736 -1244
rect 10800 -1308 10816 -1244
rect 10880 -1308 10896 -1244
rect 10960 -1308 10976 -1244
rect 11040 -1308 11056 -1244
rect 11120 -1308 11136 -1244
rect 11200 -1308 11203 -1244
rect 10014 -1325 11203 -1308
rect 10014 -1389 10016 -1325
rect 10080 -1389 10096 -1325
rect 10160 -1389 10176 -1325
rect 10240 -1389 10256 -1325
rect 10320 -1389 10336 -1325
rect 10400 -1389 10416 -1325
rect 10480 -1389 10496 -1325
rect 10560 -1389 10576 -1325
rect 10640 -1389 10656 -1325
rect 10720 -1389 10736 -1325
rect 10800 -1389 10816 -1325
rect 10880 -1389 10896 -1325
rect 10960 -1389 10976 -1325
rect 11040 -1389 11056 -1325
rect 11120 -1389 11136 -1325
rect 11200 -1389 11203 -1325
rect 10014 -1406 11203 -1389
rect 10014 -1470 10016 -1406
rect 10080 -1470 10096 -1406
rect 10160 -1470 10176 -1406
rect 10240 -1470 10256 -1406
rect 10320 -1470 10336 -1406
rect 10400 -1470 10416 -1406
rect 10480 -1470 10496 -1406
rect 10560 -1470 10576 -1406
rect 10640 -1470 10656 -1406
rect 10720 -1470 10736 -1406
rect 10800 -1470 10816 -1406
rect 10880 -1470 10896 -1406
rect 10960 -1470 10976 -1406
rect 11040 -1470 11056 -1406
rect 11120 -1470 11136 -1406
rect 11200 -1470 11203 -1406
rect 10014 -1487 11203 -1470
rect 10014 -1551 10016 -1487
rect 10080 -1551 10096 -1487
rect 10160 -1551 10176 -1487
rect 10240 -1551 10256 -1487
rect 10320 -1551 10336 -1487
rect 10400 -1551 10416 -1487
rect 10480 -1551 10496 -1487
rect 10560 -1551 10576 -1487
rect 10640 -1551 10656 -1487
rect 10720 -1551 10736 -1487
rect 10800 -1551 10816 -1487
rect 10880 -1551 10896 -1487
rect 10960 -1551 10976 -1487
rect 11040 -1551 11056 -1487
rect 11120 -1551 11136 -1487
rect 11200 -1551 11203 -1487
rect 10014 -1568 11203 -1551
rect 10014 -1632 10016 -1568
rect 10080 -1632 10096 -1568
rect 10160 -1632 10176 -1568
rect 10240 -1632 10256 -1568
rect 10320 -1632 10336 -1568
rect 10400 -1632 10416 -1568
rect 10480 -1632 10496 -1568
rect 10560 -1632 10576 -1568
rect 10640 -1632 10656 -1568
rect 10720 -1632 10736 -1568
rect 10800 -1632 10816 -1568
rect 10880 -1632 10896 -1568
rect 10960 -1632 10976 -1568
rect 11040 -1632 11056 -1568
rect 11120 -1632 11136 -1568
rect 11200 -1632 11203 -1568
rect 10014 -1649 11203 -1632
rect 10014 -1713 10016 -1649
rect 10080 -1713 10096 -1649
rect 10160 -1713 10176 -1649
rect 10240 -1713 10256 -1649
rect 10320 -1713 10336 -1649
rect 10400 -1713 10416 -1649
rect 10480 -1713 10496 -1649
rect 10560 -1713 10576 -1649
rect 10640 -1713 10656 -1649
rect 10720 -1713 10736 -1649
rect 10800 -1713 10816 -1649
rect 10880 -1713 10896 -1649
rect 10960 -1713 10976 -1649
rect 11040 -1713 11056 -1649
rect 11120 -1713 11136 -1649
rect 11200 -1713 11203 -1649
rect 10014 -1730 11203 -1713
rect 10014 -1794 10016 -1730
rect 10080 -1794 10096 -1730
rect 10160 -1794 10176 -1730
rect 10240 -1794 10256 -1730
rect 10320 -1794 10336 -1730
rect 10400 -1794 10416 -1730
rect 10480 -1794 10496 -1730
rect 10560 -1794 10576 -1730
rect 10640 -1794 10656 -1730
rect 10720 -1794 10736 -1730
rect 10800 -1794 10816 -1730
rect 10880 -1794 10896 -1730
rect 10960 -1794 10976 -1730
rect 11040 -1794 11056 -1730
rect 11120 -1794 11136 -1730
rect 11200 -1794 11203 -1730
rect 10014 -1811 11203 -1794
rect 10014 -1875 10016 -1811
rect 10080 -1875 10096 -1811
rect 10160 -1875 10176 -1811
rect 10240 -1875 10256 -1811
rect 10320 -1875 10336 -1811
rect 10400 -1875 10416 -1811
rect 10480 -1875 10496 -1811
rect 10560 -1875 10576 -1811
rect 10640 -1875 10656 -1811
rect 10720 -1875 10736 -1811
rect 10800 -1875 10816 -1811
rect 10880 -1875 10896 -1811
rect 10960 -1875 10976 -1811
rect 11040 -1875 11056 -1811
rect 11120 -1875 11136 -1811
rect 11200 -1875 11203 -1811
rect 10014 -1892 11203 -1875
rect 10014 -1956 10016 -1892
rect 10080 -1956 10096 -1892
rect 10160 -1956 10176 -1892
rect 10240 -1956 10256 -1892
rect 10320 -1956 10336 -1892
rect 10400 -1956 10416 -1892
rect 10480 -1956 10496 -1892
rect 10560 -1956 10576 -1892
rect 10640 -1956 10656 -1892
rect 10720 -1956 10736 -1892
rect 10800 -1956 10816 -1892
rect 10880 -1956 10896 -1892
rect 10960 -1956 10976 -1892
rect 11040 -1956 11056 -1892
rect 11120 -1956 11136 -1892
rect 11200 -1956 11203 -1892
rect 10014 -1973 11203 -1956
rect 10014 -2037 10016 -1973
rect 10080 -2037 10096 -1973
rect 10160 -2037 10176 -1973
rect 10240 -2037 10256 -1973
rect 10320 -2037 10336 -1973
rect 10400 -2037 10416 -1973
rect 10480 -2037 10496 -1973
rect 10560 -2037 10576 -1973
rect 10640 -2037 10656 -1973
rect 10720 -2037 10736 -1973
rect 10800 -2037 10816 -1973
rect 10880 -2037 10896 -1973
rect 10960 -2037 10976 -1973
rect 11040 -2037 11056 -1973
rect 11120 -2037 11136 -1973
rect 11200 -2037 11203 -1973
rect 10014 -2054 11203 -2037
rect 10014 -2118 10016 -2054
rect 10080 -2118 10096 -2054
rect 10160 -2118 10176 -2054
rect 10240 -2118 10256 -2054
rect 10320 -2118 10336 -2054
rect 10400 -2118 10416 -2054
rect 10480 -2118 10496 -2054
rect 10560 -2118 10576 -2054
rect 10640 -2118 10656 -2054
rect 10720 -2118 10736 -2054
rect 10800 -2118 10816 -2054
rect 10880 -2118 10896 -2054
rect 10960 -2118 10976 -2054
rect 11040 -2118 11056 -2054
rect 11120 -2118 11136 -2054
rect 11200 -2118 11203 -2054
rect 10014 -2135 11203 -2118
rect 10014 -2199 10016 -2135
rect 10080 -2199 10096 -2135
rect 10160 -2199 10176 -2135
rect 10240 -2199 10256 -2135
rect 10320 -2199 10336 -2135
rect 10400 -2199 10416 -2135
rect 10480 -2199 10496 -2135
rect 10560 -2199 10576 -2135
rect 10640 -2199 10656 -2135
rect 10720 -2199 10736 -2135
rect 10800 -2199 10816 -2135
rect 10880 -2199 10896 -2135
rect 10960 -2199 10976 -2135
rect 11040 -2199 11056 -2135
rect 11120 -2199 11136 -2135
rect 11200 -2199 11203 -2135
rect 10014 -2216 11203 -2199
rect 10014 -2280 10016 -2216
rect 10080 -2280 10096 -2216
rect 10160 -2280 10176 -2216
rect 10240 -2280 10256 -2216
rect 10320 -2280 10336 -2216
rect 10400 -2280 10416 -2216
rect 10480 -2280 10496 -2216
rect 10560 -2280 10576 -2216
rect 10640 -2280 10656 -2216
rect 10720 -2280 10736 -2216
rect 10800 -2280 10816 -2216
rect 10880 -2280 10896 -2216
rect 10960 -2280 10976 -2216
rect 11040 -2280 11056 -2216
rect 11120 -2280 11136 -2216
rect 11200 -2280 11203 -2216
rect 10014 -2297 11203 -2280
rect 10014 -2361 10016 -2297
rect 10080 -2361 10096 -2297
rect 10160 -2361 10176 -2297
rect 10240 -2361 10256 -2297
rect 10320 -2361 10336 -2297
rect 10400 -2361 10416 -2297
rect 10480 -2361 10496 -2297
rect 10560 -2361 10576 -2297
rect 10640 -2361 10656 -2297
rect 10720 -2361 10736 -2297
rect 10800 -2361 10816 -2297
rect 10880 -2361 10896 -2297
rect 10960 -2361 10976 -2297
rect 11040 -2361 11056 -2297
rect 11120 -2361 11136 -2297
rect 11200 -2361 11203 -2297
rect 10014 -2378 11203 -2361
rect 10014 -2442 10016 -2378
rect 10080 -2442 10096 -2378
rect 10160 -2442 10176 -2378
rect 10240 -2442 10256 -2378
rect 10320 -2442 10336 -2378
rect 10400 -2442 10416 -2378
rect 10480 -2442 10496 -2378
rect 10560 -2442 10576 -2378
rect 10640 -2442 10656 -2378
rect 10720 -2442 10736 -2378
rect 10800 -2442 10816 -2378
rect 10880 -2442 10896 -2378
rect 10960 -2442 10976 -2378
rect 11040 -2442 11056 -2378
rect 11120 -2442 11136 -2378
rect 11200 -2442 11203 -2378
rect 10014 -2459 11203 -2442
rect 10014 -2523 10016 -2459
rect 10080 -2523 10096 -2459
rect 10160 -2523 10176 -2459
rect 10240 -2523 10256 -2459
rect 10320 -2523 10336 -2459
rect 10400 -2523 10416 -2459
rect 10480 -2523 10496 -2459
rect 10560 -2523 10576 -2459
rect 10640 -2523 10656 -2459
rect 10720 -2523 10736 -2459
rect 10800 -2523 10816 -2459
rect 10880 -2523 10896 -2459
rect 10960 -2523 10976 -2459
rect 11040 -2523 11056 -2459
rect 11120 -2523 11136 -2459
rect 11200 -2523 11203 -2459
rect 10014 -2540 11203 -2523
rect 10014 -2604 10016 -2540
rect 10080 -2604 10096 -2540
rect 10160 -2604 10176 -2540
rect 10240 -2604 10256 -2540
rect 10320 -2604 10336 -2540
rect 10400 -2604 10416 -2540
rect 10480 -2604 10496 -2540
rect 10560 -2604 10576 -2540
rect 10640 -2604 10656 -2540
rect 10720 -2604 10736 -2540
rect 10800 -2604 10816 -2540
rect 10880 -2604 10896 -2540
rect 10960 -2604 10976 -2540
rect 11040 -2604 11056 -2540
rect 11120 -2604 11136 -2540
rect 11200 -2604 11203 -2540
rect 10014 -2621 11203 -2604
rect 10014 -2685 10016 -2621
rect 10080 -2685 10096 -2621
rect 10160 -2685 10176 -2621
rect 10240 -2685 10256 -2621
rect 10320 -2685 10336 -2621
rect 10400 -2685 10416 -2621
rect 10480 -2685 10496 -2621
rect 10560 -2685 10576 -2621
rect 10640 -2685 10656 -2621
rect 10720 -2685 10736 -2621
rect 10800 -2685 10816 -2621
rect 10880 -2685 10896 -2621
rect 10960 -2685 10976 -2621
rect 11040 -2685 11056 -2621
rect 11120 -2685 11136 -2621
rect 11200 -2685 11203 -2621
rect 10014 -2702 11203 -2685
rect 10014 -2766 10016 -2702
rect 10080 -2766 10096 -2702
rect 10160 -2766 10176 -2702
rect 10240 -2766 10256 -2702
rect 10320 -2766 10336 -2702
rect 10400 -2766 10416 -2702
rect 10480 -2766 10496 -2702
rect 10560 -2766 10576 -2702
rect 10640 -2766 10656 -2702
rect 10720 -2766 10736 -2702
rect 10800 -2766 10816 -2702
rect 10880 -2766 10896 -2702
rect 10960 -2766 10976 -2702
rect 11040 -2766 11056 -2702
rect 11120 -2766 11136 -2702
rect 11200 -2766 11203 -2702
rect 10014 -2783 11203 -2766
rect 10014 -2847 10016 -2783
rect 10080 -2847 10096 -2783
rect 10160 -2847 10176 -2783
rect 10240 -2847 10256 -2783
rect 10320 -2847 10336 -2783
rect 10400 -2847 10416 -2783
rect 10480 -2847 10496 -2783
rect 10560 -2847 10576 -2783
rect 10640 -2847 10656 -2783
rect 10720 -2847 10736 -2783
rect 10800 -2847 10816 -2783
rect 10880 -2847 10896 -2783
rect 10960 -2847 10976 -2783
rect 11040 -2847 11056 -2783
rect 11120 -2847 11136 -2783
rect 11200 -2847 11203 -2783
rect 10014 -2864 11203 -2847
rect 10014 -2928 10016 -2864
rect 10080 -2928 10096 -2864
rect 10160 -2928 10176 -2864
rect 10240 -2928 10256 -2864
rect 10320 -2928 10336 -2864
rect 10400 -2928 10416 -2864
rect 10480 -2928 10496 -2864
rect 10560 -2928 10576 -2864
rect 10640 -2928 10656 -2864
rect 10720 -2928 10736 -2864
rect 10800 -2928 10816 -2864
rect 10880 -2928 10896 -2864
rect 10960 -2928 10976 -2864
rect 11040 -2928 11056 -2864
rect 11120 -2928 11136 -2864
rect 11200 -2928 11203 -2864
rect 10014 -2945 11203 -2928
rect 10014 -3009 10016 -2945
rect 10080 -3009 10096 -2945
rect 10160 -3009 10176 -2945
rect 10240 -3009 10256 -2945
rect 10320 -3009 10336 -2945
rect 10400 -3009 10416 -2945
rect 10480 -3009 10496 -2945
rect 10560 -3009 10576 -2945
rect 10640 -3009 10656 -2945
rect 10720 -3009 10736 -2945
rect 10800 -3009 10816 -2945
rect 10880 -3009 10896 -2945
rect 10960 -3009 10976 -2945
rect 11040 -3009 11056 -2945
rect 11120 -3009 11136 -2945
rect 11200 -3009 11203 -2945
rect 10014 -3026 11203 -3009
rect 10014 -3090 10016 -3026
rect 10080 -3090 10096 -3026
rect 10160 -3090 10176 -3026
rect 10240 -3090 10256 -3026
rect 10320 -3090 10336 -3026
rect 10400 -3090 10416 -3026
rect 10480 -3090 10496 -3026
rect 10560 -3090 10576 -3026
rect 10640 -3090 10656 -3026
rect 10720 -3090 10736 -3026
rect 10800 -3090 10816 -3026
rect 10880 -3090 10896 -3026
rect 10960 -3090 10976 -3026
rect 11040 -3090 11056 -3026
rect 11120 -3090 11136 -3026
rect 11200 -3090 11203 -3026
rect 10014 -3107 11203 -3090
rect 10014 -3171 10016 -3107
rect 10080 -3171 10096 -3107
rect 10160 -3171 10176 -3107
rect 10240 -3171 10256 -3107
rect 10320 -3171 10336 -3107
rect 10400 -3171 10416 -3107
rect 10480 -3171 10496 -3107
rect 10560 -3171 10576 -3107
rect 10640 -3171 10656 -3107
rect 10720 -3171 10736 -3107
rect 10800 -3171 10816 -3107
rect 10880 -3171 10896 -3107
rect 10960 -3171 10976 -3107
rect 11040 -3171 11056 -3107
rect 11120 -3171 11136 -3107
rect 11200 -3171 11203 -3107
rect 10014 -3188 11203 -3171
rect 10014 -3252 10016 -3188
rect 10080 -3252 10096 -3188
rect 10160 -3252 10176 -3188
rect 10240 -3252 10256 -3188
rect 10320 -3252 10336 -3188
rect 10400 -3252 10416 -3188
rect 10480 -3252 10496 -3188
rect 10560 -3252 10576 -3188
rect 10640 -3252 10656 -3188
rect 10720 -3252 10736 -3188
rect 10800 -3252 10816 -3188
rect 10880 -3252 10896 -3188
rect 10960 -3252 10976 -3188
rect 11040 -3252 11056 -3188
rect 11120 -3252 11136 -3188
rect 11200 -3252 11203 -3188
rect 10014 -3269 11203 -3252
rect 10014 -3333 10016 -3269
rect 10080 -3333 10096 -3269
rect 10160 -3333 10176 -3269
rect 10240 -3333 10256 -3269
rect 10320 -3333 10336 -3269
rect 10400 -3333 10416 -3269
rect 10480 -3333 10496 -3269
rect 10560 -3333 10576 -3269
rect 10640 -3333 10656 -3269
rect 10720 -3333 10736 -3269
rect 10800 -3333 10816 -3269
rect 10880 -3333 10896 -3269
rect 10960 -3333 10976 -3269
rect 11040 -3333 11056 -3269
rect 11120 -3333 11136 -3269
rect 11200 -3333 11203 -3269
rect 10014 -3350 11203 -3333
rect 10014 -3414 10016 -3350
rect 10080 -3414 10096 -3350
rect 10160 -3414 10176 -3350
rect 10240 -3414 10256 -3350
rect 10320 -3414 10336 -3350
rect 10400 -3414 10416 -3350
rect 10480 -3414 10496 -3350
rect 10560 -3414 10576 -3350
rect 10640 -3414 10656 -3350
rect 10720 -3414 10736 -3350
rect 10800 -3414 10816 -3350
rect 10880 -3414 10896 -3350
rect 10960 -3414 10976 -3350
rect 11040 -3414 11056 -3350
rect 11120 -3414 11136 -3350
rect 11200 -3414 11203 -3350
rect 10014 -3426 11203 -3414
rect 11504 -685 11507 -621
rect 11571 -685 11587 -621
rect 11651 -685 11667 -621
rect 11731 -685 11747 -621
rect 11811 -685 11827 -621
rect 11891 -685 11907 -621
rect 11971 -685 11987 -621
rect 12051 -685 12067 -621
rect 12131 -685 12147 -621
rect 12211 -685 12227 -621
rect 12291 -685 12307 -621
rect 12371 -685 12387 -621
rect 12451 -685 12467 -621
rect 12531 -685 12547 -621
rect 12611 -685 12627 -621
rect 12691 -685 12698 -621
rect 11504 -702 12698 -685
rect 11504 -766 11507 -702
rect 11571 -766 11587 -702
rect 11651 -766 11667 -702
rect 11731 -766 11747 -702
rect 11811 -766 11827 -702
rect 11891 -766 11907 -702
rect 11971 -766 11987 -702
rect 12051 -766 12067 -702
rect 12131 -766 12147 -702
rect 12211 -766 12227 -702
rect 12291 -766 12307 -702
rect 12371 -766 12387 -702
rect 12451 -766 12467 -702
rect 12531 -766 12547 -702
rect 12611 -766 12627 -702
rect 12691 -766 12698 -702
rect 11504 -783 12698 -766
rect 11504 -847 11507 -783
rect 11571 -847 11587 -783
rect 11651 -847 11667 -783
rect 11731 -847 11747 -783
rect 11811 -847 11827 -783
rect 11891 -847 11907 -783
rect 11971 -847 11987 -783
rect 12051 -847 12067 -783
rect 12131 -847 12147 -783
rect 12211 -847 12227 -783
rect 12291 -847 12307 -783
rect 12371 -847 12387 -783
rect 12451 -847 12467 -783
rect 12531 -847 12547 -783
rect 12611 -847 12627 -783
rect 12691 -847 12698 -783
rect 11504 -864 12698 -847
rect 11504 -928 11507 -864
rect 11571 -928 11587 -864
rect 11651 -928 11667 -864
rect 11731 -928 11747 -864
rect 11811 -928 11827 -864
rect 11891 -928 11907 -864
rect 11971 -928 11987 -864
rect 12051 -928 12067 -864
rect 12131 -928 12147 -864
rect 12211 -928 12227 -864
rect 12291 -928 12307 -864
rect 12371 -928 12387 -864
rect 12451 -928 12467 -864
rect 12531 -928 12547 -864
rect 12611 -928 12627 -864
rect 12691 -928 12698 -864
rect 11504 -945 12698 -928
rect 11504 -1009 11507 -945
rect 11571 -1009 11587 -945
rect 11651 -1009 11667 -945
rect 11731 -1009 11747 -945
rect 11811 -1009 11827 -945
rect 11891 -1009 11907 -945
rect 11971 -1009 11987 -945
rect 12051 -1009 12067 -945
rect 12131 -1009 12147 -945
rect 12211 -1009 12227 -945
rect 12291 -1009 12307 -945
rect 12371 -1009 12387 -945
rect 12451 -1009 12467 -945
rect 12531 -1009 12547 -945
rect 12611 -1009 12627 -945
rect 12691 -1009 12698 -945
rect 11504 -1026 12698 -1009
rect 11504 -1090 11507 -1026
rect 11571 -1090 11587 -1026
rect 11651 -1090 11667 -1026
rect 11731 -1090 11747 -1026
rect 11811 -1090 11827 -1026
rect 11891 -1090 11907 -1026
rect 11971 -1090 11987 -1026
rect 12051 -1090 12067 -1026
rect 12131 -1090 12147 -1026
rect 12211 -1090 12227 -1026
rect 12291 -1090 12307 -1026
rect 12371 -1090 12387 -1026
rect 12451 -1090 12467 -1026
rect 12531 -1090 12547 -1026
rect 12611 -1090 12627 -1026
rect 12691 -1090 12698 -1026
rect 11504 -1107 12698 -1090
rect 11504 -1171 11507 -1107
rect 11571 -1171 11587 -1107
rect 11651 -1171 11667 -1107
rect 11731 -1171 11747 -1107
rect 11811 -1171 11827 -1107
rect 11891 -1171 11907 -1107
rect 11971 -1171 11987 -1107
rect 12051 -1171 12067 -1107
rect 12131 -1171 12147 -1107
rect 12211 -1171 12227 -1107
rect 12291 -1171 12307 -1107
rect 12371 -1171 12387 -1107
rect 12451 -1171 12467 -1107
rect 12531 -1171 12547 -1107
rect 12611 -1171 12627 -1107
rect 12691 -1171 12698 -1107
rect 11504 -1188 12698 -1171
rect 11504 -1252 11507 -1188
rect 11571 -1252 11587 -1188
rect 11651 -1252 11667 -1188
rect 11731 -1252 11747 -1188
rect 11811 -1252 11827 -1188
rect 11891 -1252 11907 -1188
rect 11971 -1252 11987 -1188
rect 12051 -1252 12067 -1188
rect 12131 -1252 12147 -1188
rect 12211 -1252 12227 -1188
rect 12291 -1252 12307 -1188
rect 12371 -1252 12387 -1188
rect 12451 -1252 12467 -1188
rect 12531 -1252 12547 -1188
rect 12611 -1252 12627 -1188
rect 12691 -1252 12698 -1188
rect 11504 -1269 12698 -1252
rect 11504 -1333 11507 -1269
rect 11571 -1333 11587 -1269
rect 11651 -1333 11667 -1269
rect 11731 -1333 11747 -1269
rect 11811 -1333 11827 -1269
rect 11891 -1333 11907 -1269
rect 11971 -1333 11987 -1269
rect 12051 -1333 12067 -1269
rect 12131 -1333 12147 -1269
rect 12211 -1333 12227 -1269
rect 12291 -1333 12307 -1269
rect 12371 -1333 12387 -1269
rect 12451 -1333 12467 -1269
rect 12531 -1333 12547 -1269
rect 12611 -1333 12627 -1269
rect 12691 -1333 12698 -1269
rect 11504 -1350 12698 -1333
rect 11504 -1414 11507 -1350
rect 11571 -1414 11587 -1350
rect 11651 -1414 11667 -1350
rect 11731 -1414 11747 -1350
rect 11811 -1414 11827 -1350
rect 11891 -1414 11907 -1350
rect 11971 -1414 11987 -1350
rect 12051 -1414 12067 -1350
rect 12131 -1414 12147 -1350
rect 12211 -1414 12227 -1350
rect 12291 -1414 12307 -1350
rect 12371 -1414 12387 -1350
rect 12451 -1414 12467 -1350
rect 12531 -1414 12547 -1350
rect 12611 -1414 12627 -1350
rect 12691 -1414 12698 -1350
rect 11504 -1431 12698 -1414
rect 11504 -1495 11507 -1431
rect 11571 -1495 11587 -1431
rect 11651 -1495 11667 -1431
rect 11731 -1495 11747 -1431
rect 11811 -1495 11827 -1431
rect 11891 -1495 11907 -1431
rect 11971 -1495 11987 -1431
rect 12051 -1495 12067 -1431
rect 12131 -1495 12147 -1431
rect 12211 -1495 12227 -1431
rect 12291 -1495 12307 -1431
rect 12371 -1495 12387 -1431
rect 12451 -1495 12467 -1431
rect 12531 -1495 12547 -1431
rect 12611 -1495 12627 -1431
rect 12691 -1495 12698 -1431
rect 11504 -1512 12698 -1495
rect 11504 -1576 11507 -1512
rect 11571 -1576 11587 -1512
rect 11651 -1576 11667 -1512
rect 11731 -1576 11747 -1512
rect 11811 -1576 11827 -1512
rect 11891 -1576 11907 -1512
rect 11971 -1576 11987 -1512
rect 12051 -1576 12067 -1512
rect 12131 -1576 12147 -1512
rect 12211 -1576 12227 -1512
rect 12291 -1576 12307 -1512
rect 12371 -1576 12387 -1512
rect 12451 -1576 12467 -1512
rect 12531 -1576 12547 -1512
rect 12611 -1576 12627 -1512
rect 12691 -1576 12698 -1512
rect 11504 -1593 12698 -1576
rect 11504 -1657 11507 -1593
rect 11571 -1657 11587 -1593
rect 11651 -1657 11667 -1593
rect 11731 -1657 11747 -1593
rect 11811 -1657 11827 -1593
rect 11891 -1657 11907 -1593
rect 11971 -1657 11987 -1593
rect 12051 -1657 12067 -1593
rect 12131 -1657 12147 -1593
rect 12211 -1657 12227 -1593
rect 12291 -1657 12307 -1593
rect 12371 -1657 12387 -1593
rect 12451 -1657 12467 -1593
rect 12531 -1657 12547 -1593
rect 12611 -1657 12627 -1593
rect 12691 -1657 12698 -1593
rect 11504 -1674 12698 -1657
rect 11504 -1738 11507 -1674
rect 11571 -1738 11587 -1674
rect 11651 -1738 11667 -1674
rect 11731 -1738 11747 -1674
rect 11811 -1738 11827 -1674
rect 11891 -1738 11907 -1674
rect 11971 -1738 11987 -1674
rect 12051 -1738 12067 -1674
rect 12131 -1738 12147 -1674
rect 12211 -1738 12227 -1674
rect 12291 -1738 12307 -1674
rect 12371 -1738 12387 -1674
rect 12451 -1738 12467 -1674
rect 12531 -1738 12547 -1674
rect 12611 -1738 12627 -1674
rect 12691 -1738 12698 -1674
rect 11504 -1755 12698 -1738
rect 11504 -1819 11507 -1755
rect 11571 -1819 11587 -1755
rect 11651 -1819 11667 -1755
rect 11731 -1819 11747 -1755
rect 11811 -1819 11827 -1755
rect 11891 -1819 11907 -1755
rect 11971 -1819 11987 -1755
rect 12051 -1819 12067 -1755
rect 12131 -1819 12147 -1755
rect 12211 -1819 12227 -1755
rect 12291 -1819 12307 -1755
rect 12371 -1819 12387 -1755
rect 12451 -1819 12467 -1755
rect 12531 -1819 12547 -1755
rect 12611 -1819 12627 -1755
rect 12691 -1819 12698 -1755
rect 11504 -1836 12698 -1819
rect 11504 -1900 11507 -1836
rect 11571 -1900 11587 -1836
rect 11651 -1900 11667 -1836
rect 11731 -1900 11747 -1836
rect 11811 -1900 11827 -1836
rect 11891 -1900 11907 -1836
rect 11971 -1900 11987 -1836
rect 12051 -1900 12067 -1836
rect 12131 -1900 12147 -1836
rect 12211 -1900 12227 -1836
rect 12291 -1900 12307 -1836
rect 12371 -1900 12387 -1836
rect 12451 -1900 12467 -1836
rect 12531 -1900 12547 -1836
rect 12611 -1900 12627 -1836
rect 12691 -1900 12698 -1836
rect 11504 -1917 12698 -1900
rect 11504 -1981 11507 -1917
rect 11571 -1981 11587 -1917
rect 11651 -1981 11667 -1917
rect 11731 -1981 11747 -1917
rect 11811 -1981 11827 -1917
rect 11891 -1981 11907 -1917
rect 11971 -1981 11987 -1917
rect 12051 -1981 12067 -1917
rect 12131 -1981 12147 -1917
rect 12211 -1981 12227 -1917
rect 12291 -1981 12307 -1917
rect 12371 -1981 12387 -1917
rect 12451 -1981 12467 -1917
rect 12531 -1981 12547 -1917
rect 12611 -1981 12627 -1917
rect 12691 -1981 12698 -1917
rect 11504 -1998 12698 -1981
rect 11504 -2062 11507 -1998
rect 11571 -2062 11587 -1998
rect 11651 -2062 11667 -1998
rect 11731 -2062 11747 -1998
rect 11811 -2062 11827 -1998
rect 11891 -2062 11907 -1998
rect 11971 -2062 11987 -1998
rect 12051 -2062 12067 -1998
rect 12131 -2062 12147 -1998
rect 12211 -2062 12227 -1998
rect 12291 -2062 12307 -1998
rect 12371 -2062 12387 -1998
rect 12451 -2062 12467 -1998
rect 12531 -2062 12547 -1998
rect 12611 -2062 12627 -1998
rect 12691 -2062 12698 -1998
rect 11504 -2079 12698 -2062
rect 11504 -2143 11507 -2079
rect 11571 -2143 11587 -2079
rect 11651 -2143 11667 -2079
rect 11731 -2143 11747 -2079
rect 11811 -2143 11827 -2079
rect 11891 -2143 11907 -2079
rect 11971 -2143 11987 -2079
rect 12051 -2143 12067 -2079
rect 12131 -2143 12147 -2079
rect 12211 -2143 12227 -2079
rect 12291 -2143 12307 -2079
rect 12371 -2143 12387 -2079
rect 12451 -2143 12467 -2079
rect 12531 -2143 12547 -2079
rect 12611 -2143 12627 -2079
rect 12691 -2143 12698 -2079
rect 11504 -2160 12698 -2143
rect 11504 -2224 11507 -2160
rect 11571 -2224 11587 -2160
rect 11651 -2224 11667 -2160
rect 11731 -2224 11747 -2160
rect 11811 -2224 11827 -2160
rect 11891 -2224 11907 -2160
rect 11971 -2224 11987 -2160
rect 12051 -2224 12067 -2160
rect 12131 -2224 12147 -2160
rect 12211 -2224 12227 -2160
rect 12291 -2224 12307 -2160
rect 12371 -2224 12387 -2160
rect 12451 -2224 12467 -2160
rect 12531 -2224 12547 -2160
rect 12611 -2224 12627 -2160
rect 12691 -2224 12698 -2160
rect 11504 -2241 12698 -2224
rect 11504 -2305 11507 -2241
rect 11571 -2305 11587 -2241
rect 11651 -2305 11667 -2241
rect 11731 -2305 11747 -2241
rect 11811 -2305 11827 -2241
rect 11891 -2305 11907 -2241
rect 11971 -2305 11987 -2241
rect 12051 -2305 12067 -2241
rect 12131 -2305 12147 -2241
rect 12211 -2305 12227 -2241
rect 12291 -2305 12307 -2241
rect 12371 -2305 12387 -2241
rect 12451 -2305 12467 -2241
rect 12531 -2305 12547 -2241
rect 12611 -2305 12627 -2241
rect 12691 -2305 12698 -2241
rect 11504 -2322 12698 -2305
rect 11504 -2386 11507 -2322
rect 11571 -2386 11587 -2322
rect 11651 -2386 11667 -2322
rect 11731 -2386 11747 -2322
rect 11811 -2386 11827 -2322
rect 11891 -2386 11907 -2322
rect 11971 -2386 11987 -2322
rect 12051 -2386 12067 -2322
rect 12131 -2386 12147 -2322
rect 12211 -2386 12227 -2322
rect 12291 -2386 12307 -2322
rect 12371 -2386 12387 -2322
rect 12451 -2386 12467 -2322
rect 12531 -2386 12547 -2322
rect 12611 -2386 12627 -2322
rect 12691 -2386 12698 -2322
rect 11504 -2403 12698 -2386
rect 11504 -2467 11507 -2403
rect 11571 -2467 11587 -2403
rect 11651 -2467 11667 -2403
rect 11731 -2467 11747 -2403
rect 11811 -2467 11827 -2403
rect 11891 -2467 11907 -2403
rect 11971 -2467 11987 -2403
rect 12051 -2467 12067 -2403
rect 12131 -2467 12147 -2403
rect 12211 -2467 12227 -2403
rect 12291 -2467 12307 -2403
rect 12371 -2467 12387 -2403
rect 12451 -2467 12467 -2403
rect 12531 -2467 12547 -2403
rect 12611 -2467 12627 -2403
rect 12691 -2467 12698 -2403
rect 11504 -2484 12698 -2467
rect 11504 -2548 11507 -2484
rect 11571 -2548 11587 -2484
rect 11651 -2548 11667 -2484
rect 11731 -2548 11747 -2484
rect 11811 -2548 11827 -2484
rect 11891 -2548 11907 -2484
rect 11971 -2548 11987 -2484
rect 12051 -2548 12067 -2484
rect 12131 -2548 12147 -2484
rect 12211 -2548 12227 -2484
rect 12291 -2548 12307 -2484
rect 12371 -2548 12387 -2484
rect 12451 -2548 12467 -2484
rect 12531 -2548 12547 -2484
rect 12611 -2548 12627 -2484
rect 12691 -2548 12698 -2484
rect 11504 -2565 12698 -2548
rect 11504 -2629 11507 -2565
rect 11571 -2629 11587 -2565
rect 11651 -2629 11667 -2565
rect 11731 -2629 11747 -2565
rect 11811 -2629 11827 -2565
rect 11891 -2629 11907 -2565
rect 11971 -2629 11987 -2565
rect 12051 -2629 12067 -2565
rect 12131 -2629 12147 -2565
rect 12211 -2629 12227 -2565
rect 12291 -2629 12307 -2565
rect 12371 -2629 12387 -2565
rect 12451 -2629 12467 -2565
rect 12531 -2629 12547 -2565
rect 12611 -2629 12627 -2565
rect 12691 -2629 12698 -2565
rect 11504 -2646 12698 -2629
rect 11504 -2710 11507 -2646
rect 11571 -2710 11587 -2646
rect 11651 -2710 11667 -2646
rect 11731 -2710 11747 -2646
rect 11811 -2710 11827 -2646
rect 11891 -2710 11907 -2646
rect 11971 -2710 11987 -2646
rect 12051 -2710 12067 -2646
rect 12131 -2710 12147 -2646
rect 12211 -2710 12227 -2646
rect 12291 -2710 12307 -2646
rect 12371 -2710 12387 -2646
rect 12451 -2710 12467 -2646
rect 12531 -2710 12547 -2646
rect 12611 -2710 12627 -2646
rect 12691 -2710 12698 -2646
rect 11504 -2727 12698 -2710
rect 11504 -2791 11507 -2727
rect 11571 -2791 11587 -2727
rect 11651 -2791 11667 -2727
rect 11731 -2791 11747 -2727
rect 11811 -2791 11827 -2727
rect 11891 -2791 11907 -2727
rect 11971 -2791 11987 -2727
rect 12051 -2791 12067 -2727
rect 12131 -2791 12147 -2727
rect 12211 -2791 12227 -2727
rect 12291 -2791 12307 -2727
rect 12371 -2791 12387 -2727
rect 12451 -2791 12467 -2727
rect 12531 -2791 12547 -2727
rect 12611 -2791 12627 -2727
rect 12691 -2791 12698 -2727
rect 11504 -2808 12698 -2791
rect 11504 -2872 11507 -2808
rect 11571 -2872 11587 -2808
rect 11651 -2872 11667 -2808
rect 11731 -2872 11747 -2808
rect 11811 -2872 11827 -2808
rect 11891 -2872 11907 -2808
rect 11971 -2872 11987 -2808
rect 12051 -2872 12067 -2808
rect 12131 -2872 12147 -2808
rect 12211 -2872 12227 -2808
rect 12291 -2872 12307 -2808
rect 12371 -2872 12387 -2808
rect 12451 -2872 12467 -2808
rect 12531 -2872 12547 -2808
rect 12611 -2872 12627 -2808
rect 12691 -2872 12698 -2808
rect 11504 -2889 12698 -2872
rect 11504 -2953 11507 -2889
rect 11571 -2953 11587 -2889
rect 11651 -2953 11667 -2889
rect 11731 -2953 11747 -2889
rect 11811 -2953 11827 -2889
rect 11891 -2953 11907 -2889
rect 11971 -2953 11987 -2889
rect 12051 -2953 12067 -2889
rect 12131 -2953 12147 -2889
rect 12211 -2953 12227 -2889
rect 12291 -2953 12307 -2889
rect 12371 -2953 12387 -2889
rect 12451 -2953 12467 -2889
rect 12531 -2953 12547 -2889
rect 12611 -2953 12627 -2889
rect 12691 -2953 12698 -2889
rect 11504 -2970 12698 -2953
rect 11504 -3034 11507 -2970
rect 11571 -3034 11587 -2970
rect 11651 -3034 11667 -2970
rect 11731 -3034 11747 -2970
rect 11811 -3034 11827 -2970
rect 11891 -3034 11907 -2970
rect 11971 -3034 11987 -2970
rect 12051 -3034 12067 -2970
rect 12131 -3034 12147 -2970
rect 12211 -3034 12227 -2970
rect 12291 -3034 12307 -2970
rect 12371 -3034 12387 -2970
rect 12451 -3034 12467 -2970
rect 12531 -3034 12547 -2970
rect 12611 -3034 12627 -2970
rect 12691 -3034 12698 -2970
rect 11504 -3051 12698 -3034
rect 11504 -3115 11507 -3051
rect 11571 -3115 11587 -3051
rect 11651 -3115 11667 -3051
rect 11731 -3115 11747 -3051
rect 11811 -3115 11827 -3051
rect 11891 -3115 11907 -3051
rect 11971 -3115 11987 -3051
rect 12051 -3115 12067 -3051
rect 12131 -3115 12147 -3051
rect 12211 -3115 12227 -3051
rect 12291 -3115 12307 -3051
rect 12371 -3115 12387 -3051
rect 12451 -3115 12467 -3051
rect 12531 -3115 12547 -3051
rect 12611 -3115 12627 -3051
rect 12691 -3115 12698 -3051
rect 11504 -3132 12698 -3115
rect 11504 -3196 11507 -3132
rect 11571 -3196 11587 -3132
rect 11651 -3196 11667 -3132
rect 11731 -3196 11747 -3132
rect 11811 -3196 11827 -3132
rect 11891 -3196 11907 -3132
rect 11971 -3196 11987 -3132
rect 12051 -3196 12067 -3132
rect 12131 -3196 12147 -3132
rect 12211 -3196 12227 -3132
rect 12291 -3196 12307 -3132
rect 12371 -3196 12387 -3132
rect 12451 -3196 12467 -3132
rect 12531 -3196 12547 -3132
rect 12611 -3196 12627 -3132
rect 12691 -3196 12698 -3132
rect 11504 -3213 12698 -3196
rect 11504 -3277 11507 -3213
rect 11571 -3277 11587 -3213
rect 11651 -3277 11667 -3213
rect 11731 -3277 11747 -3213
rect 11811 -3277 11827 -3213
rect 11891 -3277 11907 -3213
rect 11971 -3277 11987 -3213
rect 12051 -3277 12067 -3213
rect 12131 -3277 12147 -3213
rect 12211 -3277 12227 -3213
rect 12291 -3277 12307 -3213
rect 12371 -3277 12387 -3213
rect 12451 -3277 12467 -3213
rect 12531 -3277 12547 -3213
rect 12611 -3277 12627 -3213
rect 12691 -3277 12698 -3213
rect 11504 -3294 12698 -3277
rect 11504 -3358 11507 -3294
rect 11571 -3358 11587 -3294
rect 11651 -3358 11667 -3294
rect 11731 -3358 11747 -3294
rect 11811 -3358 11827 -3294
rect 11891 -3358 11907 -3294
rect 11971 -3358 11987 -3294
rect 12051 -3358 12067 -3294
rect 12131 -3358 12147 -3294
rect 12211 -3358 12227 -3294
rect 12291 -3358 12307 -3294
rect 12371 -3358 12387 -3294
rect 12451 -3358 12467 -3294
rect 12531 -3358 12547 -3294
rect 12611 -3358 12627 -3294
rect 12691 -3358 12698 -3294
rect 11504 -3375 12698 -3358
rect 11504 -3439 11507 -3375
rect 11571 -3439 11587 -3375
rect 11651 -3439 11667 -3375
rect 11731 -3439 11747 -3375
rect 11811 -3439 11827 -3375
rect 11891 -3439 11907 -3375
rect 11971 -3439 11987 -3375
rect 12051 -3439 12067 -3375
rect 12131 -3439 12147 -3375
rect 12211 -3439 12227 -3375
rect 12291 -3439 12307 -3375
rect 12371 -3439 12387 -3375
rect 12451 -3439 12467 -3375
rect 12531 -3439 12547 -3375
rect 12611 -3439 12627 -3375
rect 12691 -3439 12698 -3375
rect 11504 -3456 12698 -3439
rect 11504 -3520 11507 -3456
rect 11571 -3520 11587 -3456
rect 11651 -3520 11667 -3456
rect 11731 -3520 11747 -3456
rect 11811 -3520 11827 -3456
rect 11891 -3520 11907 -3456
rect 11971 -3520 11987 -3456
rect 12051 -3520 12067 -3456
rect 12131 -3520 12147 -3456
rect 12211 -3520 12227 -3456
rect 12291 -3520 12307 -3456
rect 12371 -3520 12387 -3456
rect 12451 -3520 12467 -3456
rect 12531 -3520 12547 -3456
rect 12611 -3520 12627 -3456
rect 12691 -3520 12698 -3456
rect 11504 -3537 12698 -3520
rect 11504 -3601 11507 -3537
rect 11571 -3601 11587 -3537
rect 11651 -3601 11667 -3537
rect 11731 -3601 11747 -3537
rect 11811 -3601 11827 -3537
rect 11891 -3601 11907 -3537
rect 11971 -3601 11987 -3537
rect 12051 -3601 12067 -3537
rect 12131 -3601 12147 -3537
rect 12211 -3601 12227 -3537
rect 12291 -3601 12307 -3537
rect 12371 -3601 12387 -3537
rect 12451 -3601 12467 -3537
rect 12531 -3601 12547 -3537
rect 12611 -3601 12627 -3537
rect 12691 -3601 12698 -3537
rect 11504 -3618 12698 -3601
rect 11504 -3682 11507 -3618
rect 11571 -3682 11587 -3618
rect 11651 -3682 11667 -3618
rect 11731 -3682 11747 -3618
rect 11811 -3682 11827 -3618
rect 11891 -3682 11907 -3618
rect 11971 -3682 11987 -3618
rect 12051 -3682 12067 -3618
rect 12131 -3682 12147 -3618
rect 12211 -3682 12227 -3618
rect 12291 -3682 12307 -3618
rect 12371 -3682 12387 -3618
rect 12451 -3682 12467 -3618
rect 12531 -3682 12547 -3618
rect 12611 -3682 12627 -3618
rect 12691 -3682 12698 -3618
rect 11504 -3699 12698 -3682
rect 11504 -3763 11507 -3699
rect 11571 -3763 11587 -3699
rect 11651 -3763 11667 -3699
rect 11731 -3763 11747 -3699
rect 11811 -3763 11827 -3699
rect 11891 -3763 11907 -3699
rect 11971 -3763 11987 -3699
rect 12051 -3763 12067 -3699
rect 12131 -3763 12147 -3699
rect 12211 -3763 12227 -3699
rect 12291 -3763 12307 -3699
rect 12371 -3763 12387 -3699
rect 12451 -3763 12467 -3699
rect 12531 -3763 12547 -3699
rect 12611 -3763 12627 -3699
rect 12691 -3763 12698 -3699
rect 11504 -3780 12698 -3763
rect 11504 -3844 11507 -3780
rect 11571 -3844 11587 -3780
rect 11651 -3844 11667 -3780
rect 11731 -3844 11747 -3780
rect 11811 -3844 11827 -3780
rect 11891 -3844 11907 -3780
rect 11971 -3844 11987 -3780
rect 12051 -3844 12067 -3780
rect 12131 -3844 12147 -3780
rect 12211 -3844 12227 -3780
rect 12291 -3844 12307 -3780
rect 12371 -3844 12387 -3780
rect 12451 -3844 12467 -3780
rect 12531 -3844 12547 -3780
rect 12611 -3844 12627 -3780
rect 12691 -3844 12698 -3780
rect 11504 -3861 12698 -3844
rect 11504 -3925 11507 -3861
rect 11571 -3925 11587 -3861
rect 11651 -3925 11667 -3861
rect 11731 -3925 11747 -3861
rect 11811 -3925 11827 -3861
rect 11891 -3925 11907 -3861
rect 11971 -3925 11987 -3861
rect 12051 -3925 12067 -3861
rect 12131 -3925 12147 -3861
rect 12211 -3925 12227 -3861
rect 12291 -3925 12307 -3861
rect 12371 -3925 12387 -3861
rect 12451 -3925 12467 -3861
rect 12531 -3925 12547 -3861
rect 12611 -3925 12627 -3861
rect 12691 -3925 12698 -3861
rect 11504 -3931 12698 -3925
<< via3 >>
rect 5403 -269 5467 -205
rect 5485 -269 5549 -205
rect 5567 -269 5631 -205
rect 5649 -269 5713 -205
rect 5731 -269 5795 -205
rect 5813 -269 5877 -205
rect 5895 -269 5959 -205
rect 5976 -269 6040 -205
rect 6057 -269 6121 -205
rect 6138 -269 6202 -205
rect 6219 -269 6283 -205
rect 6300 -269 6364 -205
rect 6381 -269 6445 -205
rect 6462 -269 6526 -205
rect 5403 -349 5467 -285
rect 5485 -349 5549 -285
rect 5567 -349 5631 -285
rect 5649 -349 5713 -285
rect 5731 -349 5795 -285
rect 5813 -349 5877 -285
rect 5895 -349 5959 -285
rect 5976 -349 6040 -285
rect 6057 -349 6121 -285
rect 6138 -349 6202 -285
rect 6219 -349 6283 -285
rect 6300 -349 6364 -285
rect 6381 -349 6445 -285
rect 6462 -349 6526 -285
rect 5403 -429 5467 -365
rect 5485 -429 5549 -365
rect 5567 -429 5631 -365
rect 5649 -429 5713 -365
rect 5731 -429 5795 -365
rect 5813 -429 5877 -365
rect 5895 -429 5959 -365
rect 5976 -429 6040 -365
rect 6057 -429 6121 -365
rect 6138 -429 6202 -365
rect 6219 -429 6283 -365
rect 6300 -429 6364 -365
rect 6381 -429 6445 -365
rect 6462 -429 6526 -365
rect 5403 -509 5467 -445
rect 5485 -509 5549 -445
rect 5567 -509 5631 -445
rect 5649 -509 5713 -445
rect 5731 -509 5795 -445
rect 5813 -509 5877 -445
rect 5895 -509 5959 -445
rect 5976 -509 6040 -445
rect 6057 -509 6121 -445
rect 6138 -509 6202 -445
rect 6219 -509 6283 -445
rect 6300 -509 6364 -445
rect 6381 -509 6445 -445
rect 6462 -509 6526 -445
rect 5403 -589 5467 -525
rect 5485 -589 5549 -525
rect 5567 -589 5631 -525
rect 5649 -589 5713 -525
rect 5731 -589 5795 -525
rect 5813 -589 5877 -525
rect 5895 -589 5959 -525
rect 5976 -589 6040 -525
rect 6057 -589 6121 -525
rect 6138 -589 6202 -525
rect 6219 -589 6283 -525
rect 6300 -589 6364 -525
rect 6381 -589 6445 -525
rect 6462 -589 6526 -525
rect 5403 -669 5467 -605
rect 5485 -669 5549 -605
rect 5567 -669 5631 -605
rect 5649 -669 5713 -605
rect 5731 -669 5795 -605
rect 5813 -669 5877 -605
rect 5895 -669 5959 -605
rect 5976 -669 6040 -605
rect 6057 -669 6121 -605
rect 6138 -669 6202 -605
rect 6219 -669 6283 -605
rect 6300 -669 6364 -605
rect 6381 -669 6445 -605
rect 6462 -669 6526 -605
rect 5403 -749 5467 -685
rect 5485 -749 5549 -685
rect 5567 -749 5631 -685
rect 5649 -749 5713 -685
rect 5731 -749 5795 -685
rect 5813 -749 5877 -685
rect 5895 -749 5959 -685
rect 5976 -749 6040 -685
rect 6057 -749 6121 -685
rect 6138 -749 6202 -685
rect 6219 -749 6283 -685
rect 6300 -749 6364 -685
rect 6381 -749 6445 -685
rect 6462 -749 6526 -685
rect 5403 -829 5467 -765
rect 5485 -829 5549 -765
rect 5567 -829 5631 -765
rect 5649 -829 5713 -765
rect 5731 -829 5795 -765
rect 5813 -829 5877 -765
rect 5895 -829 5959 -765
rect 5976 -829 6040 -765
rect 6057 -829 6121 -765
rect 6138 -829 6202 -765
rect 6219 -829 6283 -765
rect 6300 -829 6364 -765
rect 6381 -829 6445 -765
rect 6462 -829 6526 -765
rect 5403 -909 5467 -845
rect 5485 -909 5549 -845
rect 5567 -909 5631 -845
rect 5649 -909 5713 -845
rect 5731 -909 5795 -845
rect 5813 -909 5877 -845
rect 5895 -909 5959 -845
rect 5976 -909 6040 -845
rect 6057 -909 6121 -845
rect 6138 -909 6202 -845
rect 6219 -909 6283 -845
rect 6300 -909 6364 -845
rect 6381 -909 6445 -845
rect 6462 -909 6526 -845
rect 5403 -989 5467 -925
rect 5485 -989 5549 -925
rect 5567 -989 5631 -925
rect 5649 -989 5713 -925
rect 5731 -989 5795 -925
rect 5813 -989 5877 -925
rect 5895 -989 5959 -925
rect 5976 -989 6040 -925
rect 6057 -989 6121 -925
rect 6138 -989 6202 -925
rect 6219 -989 6283 -925
rect 6300 -989 6364 -925
rect 6381 -989 6445 -925
rect 6462 -989 6526 -925
rect 7014 -269 7078 -205
rect 7096 -269 7160 -205
rect 7178 -269 7242 -205
rect 7260 -269 7324 -205
rect 7342 -269 7406 -205
rect 7424 -269 7488 -205
rect 7506 -269 7570 -205
rect 7587 -269 7651 -205
rect 7668 -269 7732 -205
rect 7749 -269 7813 -205
rect 7830 -269 7894 -205
rect 7911 -269 7975 -205
rect 7992 -269 8056 -205
rect 8073 -269 8137 -205
rect 7014 -349 7078 -285
rect 7096 -349 7160 -285
rect 7178 -349 7242 -285
rect 7260 -349 7324 -285
rect 7342 -349 7406 -285
rect 7424 -349 7488 -285
rect 7506 -349 7570 -285
rect 7587 -349 7651 -285
rect 7668 -349 7732 -285
rect 7749 -349 7813 -285
rect 7830 -349 7894 -285
rect 7911 -349 7975 -285
rect 7992 -349 8056 -285
rect 8073 -349 8137 -285
rect 9194 -324 9258 -260
rect 9304 -324 9368 -260
rect 9414 -324 9478 -260
rect 9528 -268 9592 -204
rect 9609 -268 9673 -204
rect 9690 -268 9754 -204
rect 9770 -268 9834 -204
rect 9850 -268 9914 -204
rect 9930 -268 9994 -204
rect 10010 -268 10074 -204
rect 10090 -268 10154 -204
rect 10170 -268 10234 -204
rect 10250 -268 10314 -204
rect 10330 -268 10394 -204
rect 10410 -268 10474 -204
rect 10490 -268 10554 -204
rect 7014 -429 7078 -365
rect 7096 -429 7160 -365
rect 7178 -429 7242 -365
rect 7260 -429 7324 -365
rect 7342 -429 7406 -365
rect 7424 -429 7488 -365
rect 7506 -429 7570 -365
rect 7587 -429 7651 -365
rect 7668 -429 7732 -365
rect 7749 -429 7813 -365
rect 7830 -429 7894 -365
rect 7911 -429 7975 -365
rect 7992 -429 8056 -365
rect 8073 -429 8137 -365
rect 7014 -509 7078 -445
rect 7096 -509 7160 -445
rect 7178 -509 7242 -445
rect 7260 -509 7324 -445
rect 7342 -509 7406 -445
rect 7424 -509 7488 -445
rect 7506 -509 7570 -445
rect 7587 -509 7651 -445
rect 7668 -509 7732 -445
rect 7749 -509 7813 -445
rect 7830 -509 7894 -445
rect 7911 -509 7975 -445
rect 7992 -509 8056 -445
rect 8073 -509 8137 -445
rect 7014 -589 7078 -525
rect 7096 -589 7160 -525
rect 7178 -589 7242 -525
rect 7260 -589 7324 -525
rect 7342 -589 7406 -525
rect 7424 -589 7488 -525
rect 7506 -589 7570 -525
rect 7587 -589 7651 -525
rect 7668 -589 7732 -525
rect 7749 -589 7813 -525
rect 7830 -589 7894 -525
rect 7911 -589 7975 -525
rect 7992 -589 8056 -525
rect 8073 -589 8137 -525
rect 7014 -669 7078 -605
rect 7096 -669 7160 -605
rect 7178 -669 7242 -605
rect 7260 -669 7324 -605
rect 7342 -669 7406 -605
rect 7424 -669 7488 -605
rect 7506 -669 7570 -605
rect 7587 -669 7651 -605
rect 7668 -669 7732 -605
rect 7749 -669 7813 -605
rect 7830 -669 7894 -605
rect 7911 -669 7975 -605
rect 7992 -669 8056 -605
rect 8073 -669 8137 -605
rect 9528 -362 9592 -298
rect 9609 -362 9673 -298
rect 9690 -362 9754 -298
rect 9770 -362 9834 -298
rect 9850 -362 9914 -298
rect 9930 -362 9994 -298
rect 10010 -362 10074 -298
rect 10090 -362 10154 -298
rect 10170 -362 10234 -298
rect 10250 -362 10314 -298
rect 10330 -362 10394 -298
rect 10410 -362 10474 -298
rect 10490 -362 10554 -298
rect 9528 -456 9592 -392
rect 9609 -456 9673 -392
rect 9690 -456 9754 -392
rect 9770 -456 9834 -392
rect 9850 -456 9914 -392
rect 9930 -456 9994 -392
rect 10010 -456 10074 -392
rect 10090 -456 10154 -392
rect 10170 -456 10234 -392
rect 10250 -456 10314 -392
rect 10330 -456 10394 -392
rect 10410 -456 10474 -392
rect 10490 -456 10554 -392
rect 10585 -398 10649 -334
rect 10695 -398 10759 -334
rect 10805 -398 10869 -334
rect 10585 -480 10649 -416
rect 10695 -480 10759 -416
rect 10805 -480 10869 -416
rect 9528 -550 9592 -486
rect 9609 -550 9673 -486
rect 9690 -550 9754 -486
rect 9770 -550 9834 -486
rect 9850 -550 9914 -486
rect 9930 -550 9994 -486
rect 10010 -550 10074 -486
rect 10090 -550 10154 -486
rect 10170 -550 10234 -486
rect 10250 -550 10314 -486
rect 10330 -550 10394 -486
rect 10410 -550 10474 -486
rect 10490 -550 10554 -486
rect 10585 -562 10649 -498
rect 10695 -562 10759 -498
rect 10805 -562 10869 -498
rect 11507 -442 12691 -218
rect 11507 -523 11571 -459
rect 11587 -523 11651 -459
rect 11667 -523 11731 -459
rect 11747 -523 11811 -459
rect 11827 -523 11891 -459
rect 11907 -523 11971 -459
rect 11987 -523 12051 -459
rect 12067 -523 12131 -459
rect 12147 -523 12211 -459
rect 12227 -523 12291 -459
rect 12307 -523 12371 -459
rect 12387 -523 12451 -459
rect 12467 -523 12531 -459
rect 12547 -523 12611 -459
rect 12627 -523 12691 -459
rect 9528 -644 9592 -580
rect 9609 -644 9673 -580
rect 9690 -644 9754 -580
rect 9770 -644 9834 -580
rect 9850 -644 9914 -580
rect 9930 -644 9994 -580
rect 10010 -644 10074 -580
rect 10090 -644 10154 -580
rect 10170 -644 10234 -580
rect 10250 -644 10314 -580
rect 10330 -644 10394 -580
rect 10410 -644 10474 -580
rect 10490 -644 10554 -580
rect 10585 -644 10649 -580
rect 10695 -644 10759 -580
rect 10805 -644 10869 -580
rect 11507 -604 11571 -540
rect 11587 -604 11651 -540
rect 11667 -604 11731 -540
rect 11747 -604 11811 -540
rect 11827 -604 11891 -540
rect 11907 -604 11971 -540
rect 11987 -604 12051 -540
rect 12067 -604 12131 -540
rect 12147 -604 12211 -540
rect 12227 -604 12291 -540
rect 12307 -604 12371 -540
rect 12387 -604 12451 -540
rect 12467 -604 12531 -540
rect 12547 -604 12611 -540
rect 12627 -604 12691 -540
rect 7014 -749 7078 -685
rect 7096 -749 7160 -685
rect 7178 -749 7242 -685
rect 7260 -749 7324 -685
rect 7342 -749 7406 -685
rect 7424 -749 7488 -685
rect 7506 -749 7570 -685
rect 7587 -749 7651 -685
rect 7668 -749 7732 -685
rect 7749 -749 7813 -685
rect 7830 -749 7894 -685
rect 7911 -749 7975 -685
rect 7992 -749 8056 -685
rect 8073 -749 8137 -685
rect 7014 -829 7078 -765
rect 7096 -829 7160 -765
rect 7178 -829 7242 -765
rect 7260 -829 7324 -765
rect 7342 -829 7406 -765
rect 7424 -829 7488 -765
rect 7506 -829 7570 -765
rect 7587 -829 7651 -765
rect 7668 -829 7732 -765
rect 7749 -829 7813 -765
rect 7830 -829 7894 -765
rect 7911 -829 7975 -765
rect 7992 -829 8056 -765
rect 8073 -829 8137 -765
rect 7014 -909 7078 -845
rect 7096 -909 7160 -845
rect 7178 -909 7242 -845
rect 7260 -909 7324 -845
rect 7342 -909 7406 -845
rect 7424 -909 7488 -845
rect 7506 -909 7570 -845
rect 7587 -909 7651 -845
rect 7668 -909 7732 -845
rect 7749 -909 7813 -845
rect 7830 -909 7894 -845
rect 7911 -909 7975 -845
rect 7992 -909 8056 -845
rect 8073 -909 8137 -845
rect 9771 -743 9835 -679
rect 9905 -743 9969 -679
rect 9771 -880 9835 -816
rect 9905 -880 9969 -816
rect 7014 -989 7078 -925
rect 7096 -989 7160 -925
rect 7178 -989 7242 -925
rect 7260 -989 7324 -925
rect 7342 -989 7406 -925
rect 7424 -989 7488 -925
rect 7506 -989 7570 -925
rect 7587 -989 7651 -925
rect 7668 -989 7732 -925
rect 7749 -989 7813 -925
rect 7830 -989 7894 -925
rect 7911 -989 7975 -925
rect 7992 -989 8056 -925
rect 8073 -989 8137 -925
rect 10016 -903 11200 -679
rect 10016 -984 10080 -920
rect 10096 -984 10160 -920
rect 10176 -984 10240 -920
rect 10256 -984 10320 -920
rect 10336 -984 10400 -920
rect 10416 -984 10480 -920
rect 10496 -984 10560 -920
rect 10576 -984 10640 -920
rect 10656 -984 10720 -920
rect 10736 -984 10800 -920
rect 10816 -984 10880 -920
rect 10896 -984 10960 -920
rect 10976 -984 11040 -920
rect 11056 -984 11120 -920
rect 11136 -984 11200 -920
rect 10016 -1065 10080 -1001
rect 10096 -1065 10160 -1001
rect 10176 -1065 10240 -1001
rect 10256 -1065 10320 -1001
rect 10336 -1065 10400 -1001
rect 10416 -1065 10480 -1001
rect 10496 -1065 10560 -1001
rect 10576 -1065 10640 -1001
rect 10656 -1065 10720 -1001
rect 10736 -1065 10800 -1001
rect 10816 -1065 10880 -1001
rect 10896 -1065 10960 -1001
rect 10976 -1065 11040 -1001
rect 11056 -1065 11120 -1001
rect 11136 -1065 11200 -1001
rect 10016 -1146 10080 -1082
rect 10096 -1146 10160 -1082
rect 10176 -1146 10240 -1082
rect 10256 -1146 10320 -1082
rect 10336 -1146 10400 -1082
rect 10416 -1146 10480 -1082
rect 10496 -1146 10560 -1082
rect 10576 -1146 10640 -1082
rect 10656 -1146 10720 -1082
rect 10736 -1146 10800 -1082
rect 10816 -1146 10880 -1082
rect 10896 -1146 10960 -1082
rect 10976 -1146 11040 -1082
rect 11056 -1146 11120 -1082
rect 11136 -1146 11200 -1082
rect 10016 -1227 10080 -1163
rect 10096 -1227 10160 -1163
rect 10176 -1227 10240 -1163
rect 10256 -1227 10320 -1163
rect 10336 -1227 10400 -1163
rect 10416 -1227 10480 -1163
rect 10496 -1227 10560 -1163
rect 10576 -1227 10640 -1163
rect 10656 -1227 10720 -1163
rect 10736 -1227 10800 -1163
rect 10816 -1227 10880 -1163
rect 10896 -1227 10960 -1163
rect 10976 -1227 11040 -1163
rect 11056 -1227 11120 -1163
rect 11136 -1227 11200 -1163
rect 10016 -1308 10080 -1244
rect 10096 -1308 10160 -1244
rect 10176 -1308 10240 -1244
rect 10256 -1308 10320 -1244
rect 10336 -1308 10400 -1244
rect 10416 -1308 10480 -1244
rect 10496 -1308 10560 -1244
rect 10576 -1308 10640 -1244
rect 10656 -1308 10720 -1244
rect 10736 -1308 10800 -1244
rect 10816 -1308 10880 -1244
rect 10896 -1308 10960 -1244
rect 10976 -1308 11040 -1244
rect 11056 -1308 11120 -1244
rect 11136 -1308 11200 -1244
rect 10016 -1389 10080 -1325
rect 10096 -1389 10160 -1325
rect 10176 -1389 10240 -1325
rect 10256 -1389 10320 -1325
rect 10336 -1389 10400 -1325
rect 10416 -1389 10480 -1325
rect 10496 -1389 10560 -1325
rect 10576 -1389 10640 -1325
rect 10656 -1389 10720 -1325
rect 10736 -1389 10800 -1325
rect 10816 -1389 10880 -1325
rect 10896 -1389 10960 -1325
rect 10976 -1389 11040 -1325
rect 11056 -1389 11120 -1325
rect 11136 -1389 11200 -1325
rect 10016 -1470 10080 -1406
rect 10096 -1470 10160 -1406
rect 10176 -1470 10240 -1406
rect 10256 -1470 10320 -1406
rect 10336 -1470 10400 -1406
rect 10416 -1470 10480 -1406
rect 10496 -1470 10560 -1406
rect 10576 -1470 10640 -1406
rect 10656 -1470 10720 -1406
rect 10736 -1470 10800 -1406
rect 10816 -1470 10880 -1406
rect 10896 -1470 10960 -1406
rect 10976 -1470 11040 -1406
rect 11056 -1470 11120 -1406
rect 11136 -1470 11200 -1406
rect 10016 -1551 10080 -1487
rect 10096 -1551 10160 -1487
rect 10176 -1551 10240 -1487
rect 10256 -1551 10320 -1487
rect 10336 -1551 10400 -1487
rect 10416 -1551 10480 -1487
rect 10496 -1551 10560 -1487
rect 10576 -1551 10640 -1487
rect 10656 -1551 10720 -1487
rect 10736 -1551 10800 -1487
rect 10816 -1551 10880 -1487
rect 10896 -1551 10960 -1487
rect 10976 -1551 11040 -1487
rect 11056 -1551 11120 -1487
rect 11136 -1551 11200 -1487
rect 10016 -1632 10080 -1568
rect 10096 -1632 10160 -1568
rect 10176 -1632 10240 -1568
rect 10256 -1632 10320 -1568
rect 10336 -1632 10400 -1568
rect 10416 -1632 10480 -1568
rect 10496 -1632 10560 -1568
rect 10576 -1632 10640 -1568
rect 10656 -1632 10720 -1568
rect 10736 -1632 10800 -1568
rect 10816 -1632 10880 -1568
rect 10896 -1632 10960 -1568
rect 10976 -1632 11040 -1568
rect 11056 -1632 11120 -1568
rect 11136 -1632 11200 -1568
rect 10016 -1713 10080 -1649
rect 10096 -1713 10160 -1649
rect 10176 -1713 10240 -1649
rect 10256 -1713 10320 -1649
rect 10336 -1713 10400 -1649
rect 10416 -1713 10480 -1649
rect 10496 -1713 10560 -1649
rect 10576 -1713 10640 -1649
rect 10656 -1713 10720 -1649
rect 10736 -1713 10800 -1649
rect 10816 -1713 10880 -1649
rect 10896 -1713 10960 -1649
rect 10976 -1713 11040 -1649
rect 11056 -1713 11120 -1649
rect 11136 -1713 11200 -1649
rect 10016 -1794 10080 -1730
rect 10096 -1794 10160 -1730
rect 10176 -1794 10240 -1730
rect 10256 -1794 10320 -1730
rect 10336 -1794 10400 -1730
rect 10416 -1794 10480 -1730
rect 10496 -1794 10560 -1730
rect 10576 -1794 10640 -1730
rect 10656 -1794 10720 -1730
rect 10736 -1794 10800 -1730
rect 10816 -1794 10880 -1730
rect 10896 -1794 10960 -1730
rect 10976 -1794 11040 -1730
rect 11056 -1794 11120 -1730
rect 11136 -1794 11200 -1730
rect 10016 -1875 10080 -1811
rect 10096 -1875 10160 -1811
rect 10176 -1875 10240 -1811
rect 10256 -1875 10320 -1811
rect 10336 -1875 10400 -1811
rect 10416 -1875 10480 -1811
rect 10496 -1875 10560 -1811
rect 10576 -1875 10640 -1811
rect 10656 -1875 10720 -1811
rect 10736 -1875 10800 -1811
rect 10816 -1875 10880 -1811
rect 10896 -1875 10960 -1811
rect 10976 -1875 11040 -1811
rect 11056 -1875 11120 -1811
rect 11136 -1875 11200 -1811
rect 10016 -1956 10080 -1892
rect 10096 -1956 10160 -1892
rect 10176 -1956 10240 -1892
rect 10256 -1956 10320 -1892
rect 10336 -1956 10400 -1892
rect 10416 -1956 10480 -1892
rect 10496 -1956 10560 -1892
rect 10576 -1956 10640 -1892
rect 10656 -1956 10720 -1892
rect 10736 -1956 10800 -1892
rect 10816 -1956 10880 -1892
rect 10896 -1956 10960 -1892
rect 10976 -1956 11040 -1892
rect 11056 -1956 11120 -1892
rect 11136 -1956 11200 -1892
rect 10016 -2037 10080 -1973
rect 10096 -2037 10160 -1973
rect 10176 -2037 10240 -1973
rect 10256 -2037 10320 -1973
rect 10336 -2037 10400 -1973
rect 10416 -2037 10480 -1973
rect 10496 -2037 10560 -1973
rect 10576 -2037 10640 -1973
rect 10656 -2037 10720 -1973
rect 10736 -2037 10800 -1973
rect 10816 -2037 10880 -1973
rect 10896 -2037 10960 -1973
rect 10976 -2037 11040 -1973
rect 11056 -2037 11120 -1973
rect 11136 -2037 11200 -1973
rect 10016 -2118 10080 -2054
rect 10096 -2118 10160 -2054
rect 10176 -2118 10240 -2054
rect 10256 -2118 10320 -2054
rect 10336 -2118 10400 -2054
rect 10416 -2118 10480 -2054
rect 10496 -2118 10560 -2054
rect 10576 -2118 10640 -2054
rect 10656 -2118 10720 -2054
rect 10736 -2118 10800 -2054
rect 10816 -2118 10880 -2054
rect 10896 -2118 10960 -2054
rect 10976 -2118 11040 -2054
rect 11056 -2118 11120 -2054
rect 11136 -2118 11200 -2054
rect 10016 -2199 10080 -2135
rect 10096 -2199 10160 -2135
rect 10176 -2199 10240 -2135
rect 10256 -2199 10320 -2135
rect 10336 -2199 10400 -2135
rect 10416 -2199 10480 -2135
rect 10496 -2199 10560 -2135
rect 10576 -2199 10640 -2135
rect 10656 -2199 10720 -2135
rect 10736 -2199 10800 -2135
rect 10816 -2199 10880 -2135
rect 10896 -2199 10960 -2135
rect 10976 -2199 11040 -2135
rect 11056 -2199 11120 -2135
rect 11136 -2199 11200 -2135
rect 10016 -2280 10080 -2216
rect 10096 -2280 10160 -2216
rect 10176 -2280 10240 -2216
rect 10256 -2280 10320 -2216
rect 10336 -2280 10400 -2216
rect 10416 -2280 10480 -2216
rect 10496 -2280 10560 -2216
rect 10576 -2280 10640 -2216
rect 10656 -2280 10720 -2216
rect 10736 -2280 10800 -2216
rect 10816 -2280 10880 -2216
rect 10896 -2280 10960 -2216
rect 10976 -2280 11040 -2216
rect 11056 -2280 11120 -2216
rect 11136 -2280 11200 -2216
rect 10016 -2361 10080 -2297
rect 10096 -2361 10160 -2297
rect 10176 -2361 10240 -2297
rect 10256 -2361 10320 -2297
rect 10336 -2361 10400 -2297
rect 10416 -2361 10480 -2297
rect 10496 -2361 10560 -2297
rect 10576 -2361 10640 -2297
rect 10656 -2361 10720 -2297
rect 10736 -2361 10800 -2297
rect 10816 -2361 10880 -2297
rect 10896 -2361 10960 -2297
rect 10976 -2361 11040 -2297
rect 11056 -2361 11120 -2297
rect 11136 -2361 11200 -2297
rect 10016 -2442 10080 -2378
rect 10096 -2442 10160 -2378
rect 10176 -2442 10240 -2378
rect 10256 -2442 10320 -2378
rect 10336 -2442 10400 -2378
rect 10416 -2442 10480 -2378
rect 10496 -2442 10560 -2378
rect 10576 -2442 10640 -2378
rect 10656 -2442 10720 -2378
rect 10736 -2442 10800 -2378
rect 10816 -2442 10880 -2378
rect 10896 -2442 10960 -2378
rect 10976 -2442 11040 -2378
rect 11056 -2442 11120 -2378
rect 11136 -2442 11200 -2378
rect 10016 -2523 10080 -2459
rect 10096 -2523 10160 -2459
rect 10176 -2523 10240 -2459
rect 10256 -2523 10320 -2459
rect 10336 -2523 10400 -2459
rect 10416 -2523 10480 -2459
rect 10496 -2523 10560 -2459
rect 10576 -2523 10640 -2459
rect 10656 -2523 10720 -2459
rect 10736 -2523 10800 -2459
rect 10816 -2523 10880 -2459
rect 10896 -2523 10960 -2459
rect 10976 -2523 11040 -2459
rect 11056 -2523 11120 -2459
rect 11136 -2523 11200 -2459
rect 10016 -2604 10080 -2540
rect 10096 -2604 10160 -2540
rect 10176 -2604 10240 -2540
rect 10256 -2604 10320 -2540
rect 10336 -2604 10400 -2540
rect 10416 -2604 10480 -2540
rect 10496 -2604 10560 -2540
rect 10576 -2604 10640 -2540
rect 10656 -2604 10720 -2540
rect 10736 -2604 10800 -2540
rect 10816 -2604 10880 -2540
rect 10896 -2604 10960 -2540
rect 10976 -2604 11040 -2540
rect 11056 -2604 11120 -2540
rect 11136 -2604 11200 -2540
rect 10016 -2685 10080 -2621
rect 10096 -2685 10160 -2621
rect 10176 -2685 10240 -2621
rect 10256 -2685 10320 -2621
rect 10336 -2685 10400 -2621
rect 10416 -2685 10480 -2621
rect 10496 -2685 10560 -2621
rect 10576 -2685 10640 -2621
rect 10656 -2685 10720 -2621
rect 10736 -2685 10800 -2621
rect 10816 -2685 10880 -2621
rect 10896 -2685 10960 -2621
rect 10976 -2685 11040 -2621
rect 11056 -2685 11120 -2621
rect 11136 -2685 11200 -2621
rect 10016 -2766 10080 -2702
rect 10096 -2766 10160 -2702
rect 10176 -2766 10240 -2702
rect 10256 -2766 10320 -2702
rect 10336 -2766 10400 -2702
rect 10416 -2766 10480 -2702
rect 10496 -2766 10560 -2702
rect 10576 -2766 10640 -2702
rect 10656 -2766 10720 -2702
rect 10736 -2766 10800 -2702
rect 10816 -2766 10880 -2702
rect 10896 -2766 10960 -2702
rect 10976 -2766 11040 -2702
rect 11056 -2766 11120 -2702
rect 11136 -2766 11200 -2702
rect 10016 -2847 10080 -2783
rect 10096 -2847 10160 -2783
rect 10176 -2847 10240 -2783
rect 10256 -2847 10320 -2783
rect 10336 -2847 10400 -2783
rect 10416 -2847 10480 -2783
rect 10496 -2847 10560 -2783
rect 10576 -2847 10640 -2783
rect 10656 -2847 10720 -2783
rect 10736 -2847 10800 -2783
rect 10816 -2847 10880 -2783
rect 10896 -2847 10960 -2783
rect 10976 -2847 11040 -2783
rect 11056 -2847 11120 -2783
rect 11136 -2847 11200 -2783
rect 10016 -2928 10080 -2864
rect 10096 -2928 10160 -2864
rect 10176 -2928 10240 -2864
rect 10256 -2928 10320 -2864
rect 10336 -2928 10400 -2864
rect 10416 -2928 10480 -2864
rect 10496 -2928 10560 -2864
rect 10576 -2928 10640 -2864
rect 10656 -2928 10720 -2864
rect 10736 -2928 10800 -2864
rect 10816 -2928 10880 -2864
rect 10896 -2928 10960 -2864
rect 10976 -2928 11040 -2864
rect 11056 -2928 11120 -2864
rect 11136 -2928 11200 -2864
rect 10016 -3009 10080 -2945
rect 10096 -3009 10160 -2945
rect 10176 -3009 10240 -2945
rect 10256 -3009 10320 -2945
rect 10336 -3009 10400 -2945
rect 10416 -3009 10480 -2945
rect 10496 -3009 10560 -2945
rect 10576 -3009 10640 -2945
rect 10656 -3009 10720 -2945
rect 10736 -3009 10800 -2945
rect 10816 -3009 10880 -2945
rect 10896 -3009 10960 -2945
rect 10976 -3009 11040 -2945
rect 11056 -3009 11120 -2945
rect 11136 -3009 11200 -2945
rect 10016 -3090 10080 -3026
rect 10096 -3090 10160 -3026
rect 10176 -3090 10240 -3026
rect 10256 -3090 10320 -3026
rect 10336 -3090 10400 -3026
rect 10416 -3090 10480 -3026
rect 10496 -3090 10560 -3026
rect 10576 -3090 10640 -3026
rect 10656 -3090 10720 -3026
rect 10736 -3090 10800 -3026
rect 10816 -3090 10880 -3026
rect 10896 -3090 10960 -3026
rect 10976 -3090 11040 -3026
rect 11056 -3090 11120 -3026
rect 11136 -3090 11200 -3026
rect 10016 -3171 10080 -3107
rect 10096 -3171 10160 -3107
rect 10176 -3171 10240 -3107
rect 10256 -3171 10320 -3107
rect 10336 -3171 10400 -3107
rect 10416 -3171 10480 -3107
rect 10496 -3171 10560 -3107
rect 10576 -3171 10640 -3107
rect 10656 -3171 10720 -3107
rect 10736 -3171 10800 -3107
rect 10816 -3171 10880 -3107
rect 10896 -3171 10960 -3107
rect 10976 -3171 11040 -3107
rect 11056 -3171 11120 -3107
rect 11136 -3171 11200 -3107
rect 10016 -3252 10080 -3188
rect 10096 -3252 10160 -3188
rect 10176 -3252 10240 -3188
rect 10256 -3252 10320 -3188
rect 10336 -3252 10400 -3188
rect 10416 -3252 10480 -3188
rect 10496 -3252 10560 -3188
rect 10576 -3252 10640 -3188
rect 10656 -3252 10720 -3188
rect 10736 -3252 10800 -3188
rect 10816 -3252 10880 -3188
rect 10896 -3252 10960 -3188
rect 10976 -3252 11040 -3188
rect 11056 -3252 11120 -3188
rect 11136 -3252 11200 -3188
rect 10016 -3333 10080 -3269
rect 10096 -3333 10160 -3269
rect 10176 -3333 10240 -3269
rect 10256 -3333 10320 -3269
rect 10336 -3333 10400 -3269
rect 10416 -3333 10480 -3269
rect 10496 -3333 10560 -3269
rect 10576 -3333 10640 -3269
rect 10656 -3333 10720 -3269
rect 10736 -3333 10800 -3269
rect 10816 -3333 10880 -3269
rect 10896 -3333 10960 -3269
rect 10976 -3333 11040 -3269
rect 11056 -3333 11120 -3269
rect 11136 -3333 11200 -3269
rect 10016 -3414 10080 -3350
rect 10096 -3414 10160 -3350
rect 10176 -3414 10240 -3350
rect 10256 -3414 10320 -3350
rect 10336 -3414 10400 -3350
rect 10416 -3414 10480 -3350
rect 10496 -3414 10560 -3350
rect 10576 -3414 10640 -3350
rect 10656 -3414 10720 -3350
rect 10736 -3414 10800 -3350
rect 10816 -3414 10880 -3350
rect 10896 -3414 10960 -3350
rect 10976 -3414 11040 -3350
rect 11056 -3414 11120 -3350
rect 11136 -3414 11200 -3350
rect 11507 -685 11571 -621
rect 11587 -685 11651 -621
rect 11667 -685 11731 -621
rect 11747 -685 11811 -621
rect 11827 -685 11891 -621
rect 11907 -685 11971 -621
rect 11987 -685 12051 -621
rect 12067 -685 12131 -621
rect 12147 -685 12211 -621
rect 12227 -685 12291 -621
rect 12307 -685 12371 -621
rect 12387 -685 12451 -621
rect 12467 -685 12531 -621
rect 12547 -685 12611 -621
rect 12627 -685 12691 -621
rect 11507 -766 11571 -702
rect 11587 -766 11651 -702
rect 11667 -766 11731 -702
rect 11747 -766 11811 -702
rect 11827 -766 11891 -702
rect 11907 -766 11971 -702
rect 11987 -766 12051 -702
rect 12067 -766 12131 -702
rect 12147 -766 12211 -702
rect 12227 -766 12291 -702
rect 12307 -766 12371 -702
rect 12387 -766 12451 -702
rect 12467 -766 12531 -702
rect 12547 -766 12611 -702
rect 12627 -766 12691 -702
rect 11507 -847 11571 -783
rect 11587 -847 11651 -783
rect 11667 -847 11731 -783
rect 11747 -847 11811 -783
rect 11827 -847 11891 -783
rect 11907 -847 11971 -783
rect 11987 -847 12051 -783
rect 12067 -847 12131 -783
rect 12147 -847 12211 -783
rect 12227 -847 12291 -783
rect 12307 -847 12371 -783
rect 12387 -847 12451 -783
rect 12467 -847 12531 -783
rect 12547 -847 12611 -783
rect 12627 -847 12691 -783
rect 11507 -928 11571 -864
rect 11587 -928 11651 -864
rect 11667 -928 11731 -864
rect 11747 -928 11811 -864
rect 11827 -928 11891 -864
rect 11907 -928 11971 -864
rect 11987 -928 12051 -864
rect 12067 -928 12131 -864
rect 12147 -928 12211 -864
rect 12227 -928 12291 -864
rect 12307 -928 12371 -864
rect 12387 -928 12451 -864
rect 12467 -928 12531 -864
rect 12547 -928 12611 -864
rect 12627 -928 12691 -864
rect 11507 -1009 11571 -945
rect 11587 -1009 11651 -945
rect 11667 -1009 11731 -945
rect 11747 -1009 11811 -945
rect 11827 -1009 11891 -945
rect 11907 -1009 11971 -945
rect 11987 -1009 12051 -945
rect 12067 -1009 12131 -945
rect 12147 -1009 12211 -945
rect 12227 -1009 12291 -945
rect 12307 -1009 12371 -945
rect 12387 -1009 12451 -945
rect 12467 -1009 12531 -945
rect 12547 -1009 12611 -945
rect 12627 -1009 12691 -945
rect 11507 -1090 11571 -1026
rect 11587 -1090 11651 -1026
rect 11667 -1090 11731 -1026
rect 11747 -1090 11811 -1026
rect 11827 -1090 11891 -1026
rect 11907 -1090 11971 -1026
rect 11987 -1090 12051 -1026
rect 12067 -1090 12131 -1026
rect 12147 -1090 12211 -1026
rect 12227 -1090 12291 -1026
rect 12307 -1090 12371 -1026
rect 12387 -1090 12451 -1026
rect 12467 -1090 12531 -1026
rect 12547 -1090 12611 -1026
rect 12627 -1090 12691 -1026
rect 11507 -1171 11571 -1107
rect 11587 -1171 11651 -1107
rect 11667 -1171 11731 -1107
rect 11747 -1171 11811 -1107
rect 11827 -1171 11891 -1107
rect 11907 -1171 11971 -1107
rect 11987 -1171 12051 -1107
rect 12067 -1171 12131 -1107
rect 12147 -1171 12211 -1107
rect 12227 -1171 12291 -1107
rect 12307 -1171 12371 -1107
rect 12387 -1171 12451 -1107
rect 12467 -1171 12531 -1107
rect 12547 -1171 12611 -1107
rect 12627 -1171 12691 -1107
rect 11507 -1252 11571 -1188
rect 11587 -1252 11651 -1188
rect 11667 -1252 11731 -1188
rect 11747 -1252 11811 -1188
rect 11827 -1252 11891 -1188
rect 11907 -1252 11971 -1188
rect 11987 -1252 12051 -1188
rect 12067 -1252 12131 -1188
rect 12147 -1252 12211 -1188
rect 12227 -1252 12291 -1188
rect 12307 -1252 12371 -1188
rect 12387 -1252 12451 -1188
rect 12467 -1252 12531 -1188
rect 12547 -1252 12611 -1188
rect 12627 -1252 12691 -1188
rect 11507 -1333 11571 -1269
rect 11587 -1333 11651 -1269
rect 11667 -1333 11731 -1269
rect 11747 -1333 11811 -1269
rect 11827 -1333 11891 -1269
rect 11907 -1333 11971 -1269
rect 11987 -1333 12051 -1269
rect 12067 -1333 12131 -1269
rect 12147 -1333 12211 -1269
rect 12227 -1333 12291 -1269
rect 12307 -1333 12371 -1269
rect 12387 -1333 12451 -1269
rect 12467 -1333 12531 -1269
rect 12547 -1333 12611 -1269
rect 12627 -1333 12691 -1269
rect 11507 -1414 11571 -1350
rect 11587 -1414 11651 -1350
rect 11667 -1414 11731 -1350
rect 11747 -1414 11811 -1350
rect 11827 -1414 11891 -1350
rect 11907 -1414 11971 -1350
rect 11987 -1414 12051 -1350
rect 12067 -1414 12131 -1350
rect 12147 -1414 12211 -1350
rect 12227 -1414 12291 -1350
rect 12307 -1414 12371 -1350
rect 12387 -1414 12451 -1350
rect 12467 -1414 12531 -1350
rect 12547 -1414 12611 -1350
rect 12627 -1414 12691 -1350
rect 11507 -1495 11571 -1431
rect 11587 -1495 11651 -1431
rect 11667 -1495 11731 -1431
rect 11747 -1495 11811 -1431
rect 11827 -1495 11891 -1431
rect 11907 -1495 11971 -1431
rect 11987 -1495 12051 -1431
rect 12067 -1495 12131 -1431
rect 12147 -1495 12211 -1431
rect 12227 -1495 12291 -1431
rect 12307 -1495 12371 -1431
rect 12387 -1495 12451 -1431
rect 12467 -1495 12531 -1431
rect 12547 -1495 12611 -1431
rect 12627 -1495 12691 -1431
rect 11507 -1576 11571 -1512
rect 11587 -1576 11651 -1512
rect 11667 -1576 11731 -1512
rect 11747 -1576 11811 -1512
rect 11827 -1576 11891 -1512
rect 11907 -1576 11971 -1512
rect 11987 -1576 12051 -1512
rect 12067 -1576 12131 -1512
rect 12147 -1576 12211 -1512
rect 12227 -1576 12291 -1512
rect 12307 -1576 12371 -1512
rect 12387 -1576 12451 -1512
rect 12467 -1576 12531 -1512
rect 12547 -1576 12611 -1512
rect 12627 -1576 12691 -1512
rect 11507 -1657 11571 -1593
rect 11587 -1657 11651 -1593
rect 11667 -1657 11731 -1593
rect 11747 -1657 11811 -1593
rect 11827 -1657 11891 -1593
rect 11907 -1657 11971 -1593
rect 11987 -1657 12051 -1593
rect 12067 -1657 12131 -1593
rect 12147 -1657 12211 -1593
rect 12227 -1657 12291 -1593
rect 12307 -1657 12371 -1593
rect 12387 -1657 12451 -1593
rect 12467 -1657 12531 -1593
rect 12547 -1657 12611 -1593
rect 12627 -1657 12691 -1593
rect 11507 -1738 11571 -1674
rect 11587 -1738 11651 -1674
rect 11667 -1738 11731 -1674
rect 11747 -1738 11811 -1674
rect 11827 -1738 11891 -1674
rect 11907 -1738 11971 -1674
rect 11987 -1738 12051 -1674
rect 12067 -1738 12131 -1674
rect 12147 -1738 12211 -1674
rect 12227 -1738 12291 -1674
rect 12307 -1738 12371 -1674
rect 12387 -1738 12451 -1674
rect 12467 -1738 12531 -1674
rect 12547 -1738 12611 -1674
rect 12627 -1738 12691 -1674
rect 11507 -1819 11571 -1755
rect 11587 -1819 11651 -1755
rect 11667 -1819 11731 -1755
rect 11747 -1819 11811 -1755
rect 11827 -1819 11891 -1755
rect 11907 -1819 11971 -1755
rect 11987 -1819 12051 -1755
rect 12067 -1819 12131 -1755
rect 12147 -1819 12211 -1755
rect 12227 -1819 12291 -1755
rect 12307 -1819 12371 -1755
rect 12387 -1819 12451 -1755
rect 12467 -1819 12531 -1755
rect 12547 -1819 12611 -1755
rect 12627 -1819 12691 -1755
rect 11507 -1900 11571 -1836
rect 11587 -1900 11651 -1836
rect 11667 -1900 11731 -1836
rect 11747 -1900 11811 -1836
rect 11827 -1900 11891 -1836
rect 11907 -1900 11971 -1836
rect 11987 -1900 12051 -1836
rect 12067 -1900 12131 -1836
rect 12147 -1900 12211 -1836
rect 12227 -1900 12291 -1836
rect 12307 -1900 12371 -1836
rect 12387 -1900 12451 -1836
rect 12467 -1900 12531 -1836
rect 12547 -1900 12611 -1836
rect 12627 -1900 12691 -1836
rect 11507 -1981 11571 -1917
rect 11587 -1981 11651 -1917
rect 11667 -1981 11731 -1917
rect 11747 -1981 11811 -1917
rect 11827 -1981 11891 -1917
rect 11907 -1981 11971 -1917
rect 11987 -1981 12051 -1917
rect 12067 -1981 12131 -1917
rect 12147 -1981 12211 -1917
rect 12227 -1981 12291 -1917
rect 12307 -1981 12371 -1917
rect 12387 -1981 12451 -1917
rect 12467 -1981 12531 -1917
rect 12547 -1981 12611 -1917
rect 12627 -1981 12691 -1917
rect 11507 -2062 11571 -1998
rect 11587 -2062 11651 -1998
rect 11667 -2062 11731 -1998
rect 11747 -2062 11811 -1998
rect 11827 -2062 11891 -1998
rect 11907 -2062 11971 -1998
rect 11987 -2062 12051 -1998
rect 12067 -2062 12131 -1998
rect 12147 -2062 12211 -1998
rect 12227 -2062 12291 -1998
rect 12307 -2062 12371 -1998
rect 12387 -2062 12451 -1998
rect 12467 -2062 12531 -1998
rect 12547 -2062 12611 -1998
rect 12627 -2062 12691 -1998
rect 11507 -2143 11571 -2079
rect 11587 -2143 11651 -2079
rect 11667 -2143 11731 -2079
rect 11747 -2143 11811 -2079
rect 11827 -2143 11891 -2079
rect 11907 -2143 11971 -2079
rect 11987 -2143 12051 -2079
rect 12067 -2143 12131 -2079
rect 12147 -2143 12211 -2079
rect 12227 -2143 12291 -2079
rect 12307 -2143 12371 -2079
rect 12387 -2143 12451 -2079
rect 12467 -2143 12531 -2079
rect 12547 -2143 12611 -2079
rect 12627 -2143 12691 -2079
rect 11507 -2224 11571 -2160
rect 11587 -2224 11651 -2160
rect 11667 -2224 11731 -2160
rect 11747 -2224 11811 -2160
rect 11827 -2224 11891 -2160
rect 11907 -2224 11971 -2160
rect 11987 -2224 12051 -2160
rect 12067 -2224 12131 -2160
rect 12147 -2224 12211 -2160
rect 12227 -2224 12291 -2160
rect 12307 -2224 12371 -2160
rect 12387 -2224 12451 -2160
rect 12467 -2224 12531 -2160
rect 12547 -2224 12611 -2160
rect 12627 -2224 12691 -2160
rect 11507 -2305 11571 -2241
rect 11587 -2305 11651 -2241
rect 11667 -2305 11731 -2241
rect 11747 -2305 11811 -2241
rect 11827 -2305 11891 -2241
rect 11907 -2305 11971 -2241
rect 11987 -2305 12051 -2241
rect 12067 -2305 12131 -2241
rect 12147 -2305 12211 -2241
rect 12227 -2305 12291 -2241
rect 12307 -2305 12371 -2241
rect 12387 -2305 12451 -2241
rect 12467 -2305 12531 -2241
rect 12547 -2305 12611 -2241
rect 12627 -2305 12691 -2241
rect 11507 -2386 11571 -2322
rect 11587 -2386 11651 -2322
rect 11667 -2386 11731 -2322
rect 11747 -2386 11811 -2322
rect 11827 -2386 11891 -2322
rect 11907 -2386 11971 -2322
rect 11987 -2386 12051 -2322
rect 12067 -2386 12131 -2322
rect 12147 -2386 12211 -2322
rect 12227 -2386 12291 -2322
rect 12307 -2386 12371 -2322
rect 12387 -2386 12451 -2322
rect 12467 -2386 12531 -2322
rect 12547 -2386 12611 -2322
rect 12627 -2386 12691 -2322
rect 11507 -2467 11571 -2403
rect 11587 -2467 11651 -2403
rect 11667 -2467 11731 -2403
rect 11747 -2467 11811 -2403
rect 11827 -2467 11891 -2403
rect 11907 -2467 11971 -2403
rect 11987 -2467 12051 -2403
rect 12067 -2467 12131 -2403
rect 12147 -2467 12211 -2403
rect 12227 -2467 12291 -2403
rect 12307 -2467 12371 -2403
rect 12387 -2467 12451 -2403
rect 12467 -2467 12531 -2403
rect 12547 -2467 12611 -2403
rect 12627 -2467 12691 -2403
rect 11507 -2548 11571 -2484
rect 11587 -2548 11651 -2484
rect 11667 -2548 11731 -2484
rect 11747 -2548 11811 -2484
rect 11827 -2548 11891 -2484
rect 11907 -2548 11971 -2484
rect 11987 -2548 12051 -2484
rect 12067 -2548 12131 -2484
rect 12147 -2548 12211 -2484
rect 12227 -2548 12291 -2484
rect 12307 -2548 12371 -2484
rect 12387 -2548 12451 -2484
rect 12467 -2548 12531 -2484
rect 12547 -2548 12611 -2484
rect 12627 -2548 12691 -2484
rect 11507 -2629 11571 -2565
rect 11587 -2629 11651 -2565
rect 11667 -2629 11731 -2565
rect 11747 -2629 11811 -2565
rect 11827 -2629 11891 -2565
rect 11907 -2629 11971 -2565
rect 11987 -2629 12051 -2565
rect 12067 -2629 12131 -2565
rect 12147 -2629 12211 -2565
rect 12227 -2629 12291 -2565
rect 12307 -2629 12371 -2565
rect 12387 -2629 12451 -2565
rect 12467 -2629 12531 -2565
rect 12547 -2629 12611 -2565
rect 12627 -2629 12691 -2565
rect 11507 -2710 11571 -2646
rect 11587 -2710 11651 -2646
rect 11667 -2710 11731 -2646
rect 11747 -2710 11811 -2646
rect 11827 -2710 11891 -2646
rect 11907 -2710 11971 -2646
rect 11987 -2710 12051 -2646
rect 12067 -2710 12131 -2646
rect 12147 -2710 12211 -2646
rect 12227 -2710 12291 -2646
rect 12307 -2710 12371 -2646
rect 12387 -2710 12451 -2646
rect 12467 -2710 12531 -2646
rect 12547 -2710 12611 -2646
rect 12627 -2710 12691 -2646
rect 11507 -2791 11571 -2727
rect 11587 -2791 11651 -2727
rect 11667 -2791 11731 -2727
rect 11747 -2791 11811 -2727
rect 11827 -2791 11891 -2727
rect 11907 -2791 11971 -2727
rect 11987 -2791 12051 -2727
rect 12067 -2791 12131 -2727
rect 12147 -2791 12211 -2727
rect 12227 -2791 12291 -2727
rect 12307 -2791 12371 -2727
rect 12387 -2791 12451 -2727
rect 12467 -2791 12531 -2727
rect 12547 -2791 12611 -2727
rect 12627 -2791 12691 -2727
rect 11507 -2872 11571 -2808
rect 11587 -2872 11651 -2808
rect 11667 -2872 11731 -2808
rect 11747 -2872 11811 -2808
rect 11827 -2872 11891 -2808
rect 11907 -2872 11971 -2808
rect 11987 -2872 12051 -2808
rect 12067 -2872 12131 -2808
rect 12147 -2872 12211 -2808
rect 12227 -2872 12291 -2808
rect 12307 -2872 12371 -2808
rect 12387 -2872 12451 -2808
rect 12467 -2872 12531 -2808
rect 12547 -2872 12611 -2808
rect 12627 -2872 12691 -2808
rect 11507 -2953 11571 -2889
rect 11587 -2953 11651 -2889
rect 11667 -2953 11731 -2889
rect 11747 -2953 11811 -2889
rect 11827 -2953 11891 -2889
rect 11907 -2953 11971 -2889
rect 11987 -2953 12051 -2889
rect 12067 -2953 12131 -2889
rect 12147 -2953 12211 -2889
rect 12227 -2953 12291 -2889
rect 12307 -2953 12371 -2889
rect 12387 -2953 12451 -2889
rect 12467 -2953 12531 -2889
rect 12547 -2953 12611 -2889
rect 12627 -2953 12691 -2889
rect 11507 -3034 11571 -2970
rect 11587 -3034 11651 -2970
rect 11667 -3034 11731 -2970
rect 11747 -3034 11811 -2970
rect 11827 -3034 11891 -2970
rect 11907 -3034 11971 -2970
rect 11987 -3034 12051 -2970
rect 12067 -3034 12131 -2970
rect 12147 -3034 12211 -2970
rect 12227 -3034 12291 -2970
rect 12307 -3034 12371 -2970
rect 12387 -3034 12451 -2970
rect 12467 -3034 12531 -2970
rect 12547 -3034 12611 -2970
rect 12627 -3034 12691 -2970
rect 11507 -3115 11571 -3051
rect 11587 -3115 11651 -3051
rect 11667 -3115 11731 -3051
rect 11747 -3115 11811 -3051
rect 11827 -3115 11891 -3051
rect 11907 -3115 11971 -3051
rect 11987 -3115 12051 -3051
rect 12067 -3115 12131 -3051
rect 12147 -3115 12211 -3051
rect 12227 -3115 12291 -3051
rect 12307 -3115 12371 -3051
rect 12387 -3115 12451 -3051
rect 12467 -3115 12531 -3051
rect 12547 -3115 12611 -3051
rect 12627 -3115 12691 -3051
rect 11507 -3196 11571 -3132
rect 11587 -3196 11651 -3132
rect 11667 -3196 11731 -3132
rect 11747 -3196 11811 -3132
rect 11827 -3196 11891 -3132
rect 11907 -3196 11971 -3132
rect 11987 -3196 12051 -3132
rect 12067 -3196 12131 -3132
rect 12147 -3196 12211 -3132
rect 12227 -3196 12291 -3132
rect 12307 -3196 12371 -3132
rect 12387 -3196 12451 -3132
rect 12467 -3196 12531 -3132
rect 12547 -3196 12611 -3132
rect 12627 -3196 12691 -3132
rect 11507 -3277 11571 -3213
rect 11587 -3277 11651 -3213
rect 11667 -3277 11731 -3213
rect 11747 -3277 11811 -3213
rect 11827 -3277 11891 -3213
rect 11907 -3277 11971 -3213
rect 11987 -3277 12051 -3213
rect 12067 -3277 12131 -3213
rect 12147 -3277 12211 -3213
rect 12227 -3277 12291 -3213
rect 12307 -3277 12371 -3213
rect 12387 -3277 12451 -3213
rect 12467 -3277 12531 -3213
rect 12547 -3277 12611 -3213
rect 12627 -3277 12691 -3213
rect 11507 -3358 11571 -3294
rect 11587 -3358 11651 -3294
rect 11667 -3358 11731 -3294
rect 11747 -3358 11811 -3294
rect 11827 -3358 11891 -3294
rect 11907 -3358 11971 -3294
rect 11987 -3358 12051 -3294
rect 12067 -3358 12131 -3294
rect 12147 -3358 12211 -3294
rect 12227 -3358 12291 -3294
rect 12307 -3358 12371 -3294
rect 12387 -3358 12451 -3294
rect 12467 -3358 12531 -3294
rect 12547 -3358 12611 -3294
rect 12627 -3358 12691 -3294
rect 11507 -3439 11571 -3375
rect 11587 -3439 11651 -3375
rect 11667 -3439 11731 -3375
rect 11747 -3439 11811 -3375
rect 11827 -3439 11891 -3375
rect 11907 -3439 11971 -3375
rect 11987 -3439 12051 -3375
rect 12067 -3439 12131 -3375
rect 12147 -3439 12211 -3375
rect 12227 -3439 12291 -3375
rect 12307 -3439 12371 -3375
rect 12387 -3439 12451 -3375
rect 12467 -3439 12531 -3375
rect 12547 -3439 12611 -3375
rect 12627 -3439 12691 -3375
rect 11507 -3520 11571 -3456
rect 11587 -3520 11651 -3456
rect 11667 -3520 11731 -3456
rect 11747 -3520 11811 -3456
rect 11827 -3520 11891 -3456
rect 11907 -3520 11971 -3456
rect 11987 -3520 12051 -3456
rect 12067 -3520 12131 -3456
rect 12147 -3520 12211 -3456
rect 12227 -3520 12291 -3456
rect 12307 -3520 12371 -3456
rect 12387 -3520 12451 -3456
rect 12467 -3520 12531 -3456
rect 12547 -3520 12611 -3456
rect 12627 -3520 12691 -3456
rect 11507 -3601 11571 -3537
rect 11587 -3601 11651 -3537
rect 11667 -3601 11731 -3537
rect 11747 -3601 11811 -3537
rect 11827 -3601 11891 -3537
rect 11907 -3601 11971 -3537
rect 11987 -3601 12051 -3537
rect 12067 -3601 12131 -3537
rect 12147 -3601 12211 -3537
rect 12227 -3601 12291 -3537
rect 12307 -3601 12371 -3537
rect 12387 -3601 12451 -3537
rect 12467 -3601 12531 -3537
rect 12547 -3601 12611 -3537
rect 12627 -3601 12691 -3537
rect 11507 -3682 11571 -3618
rect 11587 -3682 11651 -3618
rect 11667 -3682 11731 -3618
rect 11747 -3682 11811 -3618
rect 11827 -3682 11891 -3618
rect 11907 -3682 11971 -3618
rect 11987 -3682 12051 -3618
rect 12067 -3682 12131 -3618
rect 12147 -3682 12211 -3618
rect 12227 -3682 12291 -3618
rect 12307 -3682 12371 -3618
rect 12387 -3682 12451 -3618
rect 12467 -3682 12531 -3618
rect 12547 -3682 12611 -3618
rect 12627 -3682 12691 -3618
rect 11507 -3763 11571 -3699
rect 11587 -3763 11651 -3699
rect 11667 -3763 11731 -3699
rect 11747 -3763 11811 -3699
rect 11827 -3763 11891 -3699
rect 11907 -3763 11971 -3699
rect 11987 -3763 12051 -3699
rect 12067 -3763 12131 -3699
rect 12147 -3763 12211 -3699
rect 12227 -3763 12291 -3699
rect 12307 -3763 12371 -3699
rect 12387 -3763 12451 -3699
rect 12467 -3763 12531 -3699
rect 12547 -3763 12611 -3699
rect 12627 -3763 12691 -3699
rect 11507 -3844 11571 -3780
rect 11587 -3844 11651 -3780
rect 11667 -3844 11731 -3780
rect 11747 -3844 11811 -3780
rect 11827 -3844 11891 -3780
rect 11907 -3844 11971 -3780
rect 11987 -3844 12051 -3780
rect 12067 -3844 12131 -3780
rect 12147 -3844 12211 -3780
rect 12227 -3844 12291 -3780
rect 12307 -3844 12371 -3780
rect 12387 -3844 12451 -3780
rect 12467 -3844 12531 -3780
rect 12547 -3844 12611 -3780
rect 12627 -3844 12691 -3780
rect 11507 -3925 11571 -3861
rect 11587 -3925 11651 -3861
rect 11667 -3925 11731 -3861
rect 11747 -3925 11811 -3861
rect 11827 -3925 11891 -3861
rect 11907 -3925 11971 -3861
rect 11987 -3925 12051 -3861
rect 12067 -3925 12131 -3861
rect 12147 -3925 12211 -3861
rect 12227 -3925 12291 -3861
rect 12307 -3925 12371 -3861
rect 12387 -3925 12451 -3861
rect 12467 -3925 12531 -3861
rect 12547 -3925 12611 -3861
rect 12627 -3925 12691 -3861
<< metal4 >>
rect 5402 -205 8138 -202
rect 5402 -269 5403 -205
rect 5467 -269 5485 -205
rect 5549 -269 5567 -205
rect 5631 -269 5649 -205
rect 5713 -269 5731 -205
rect 5795 -269 5813 -205
rect 5877 -269 5895 -205
rect 5959 -269 5976 -205
rect 6040 -269 6057 -205
rect 6121 -269 6138 -205
rect 6202 -269 6219 -205
rect 6283 -269 6300 -205
rect 6364 -269 6381 -205
rect 6445 -269 6462 -205
rect 6526 -269 7014 -205
rect 7078 -269 7096 -205
rect 7160 -269 7178 -205
rect 7242 -269 7260 -205
rect 7324 -269 7342 -205
rect 7406 -269 7424 -205
rect 7488 -269 7506 -205
rect 7570 -269 7587 -205
rect 7651 -269 7668 -205
rect 7732 -269 7749 -205
rect 7813 -269 7830 -205
rect 7894 -269 7911 -205
rect 7975 -269 7992 -205
rect 8056 -269 8073 -205
rect 8137 -269 8138 -205
rect 5402 -285 8138 -269
rect 5402 -349 5403 -285
rect 5467 -349 5485 -285
rect 5549 -349 5567 -285
rect 5631 -349 5649 -285
rect 5713 -349 5731 -285
rect 5795 -349 5813 -285
rect 5877 -349 5895 -285
rect 5959 -349 5976 -285
rect 6040 -349 6057 -285
rect 6121 -349 6138 -285
rect 6202 -349 6219 -285
rect 6283 -349 6300 -285
rect 6364 -349 6381 -285
rect 6445 -349 6462 -285
rect 6526 -349 7014 -285
rect 7078 -349 7096 -285
rect 7160 -349 7178 -285
rect 7242 -349 7260 -285
rect 7324 -349 7342 -285
rect 7406 -349 7424 -285
rect 7488 -349 7506 -285
rect 7570 -349 7587 -285
rect 7651 -349 7668 -285
rect 7732 -349 7749 -285
rect 7813 -349 7830 -285
rect 7894 -349 7911 -285
rect 7975 -349 7992 -285
rect 8056 -349 8073 -285
rect 8137 -349 8138 -285
rect 9193 -260 9479 -203
rect 9193 -324 9194 -260
rect 9258 -324 9304 -260
rect 9368 -324 9414 -260
rect 9478 -324 9479 -260
rect 9193 -325 9479 -324
rect 9527 -204 10555 -202
rect 9527 -268 9528 -204
rect 9592 -268 9609 -204
rect 9673 -268 9690 -204
rect 9754 -268 9770 -204
rect 9834 -268 9850 -204
rect 9914 -268 9930 -204
rect 9994 -268 10010 -204
rect 10074 -268 10090 -204
rect 10154 -268 10170 -204
rect 10234 -268 10250 -204
rect 10314 -268 10330 -204
rect 10394 -268 10410 -204
rect 10474 -268 10490 -204
rect 10554 -268 10555 -204
rect 9527 -298 10555 -268
rect 5402 -359 8138 -349
rect 5402 -365 6527 -359
rect 5402 -429 5403 -365
rect 5467 -429 5485 -365
rect 5549 -429 5567 -365
rect 5631 -429 5649 -365
rect 5713 -429 5731 -365
rect 5795 -429 5813 -365
rect 5877 -429 5895 -365
rect 5959 -429 5976 -365
rect 6040 -429 6057 -365
rect 6121 -429 6138 -365
rect 6202 -429 6219 -365
rect 6283 -429 6300 -365
rect 6364 -429 6381 -365
rect 6445 -429 6462 -365
rect 6526 -429 6527 -365
rect 5402 -445 6527 -429
rect 5402 -509 5403 -445
rect 5467 -509 5485 -445
rect 5549 -509 5567 -445
rect 5631 -509 5649 -445
rect 5713 -509 5731 -445
rect 5795 -509 5813 -445
rect 5877 -509 5895 -445
rect 5959 -509 5976 -445
rect 6040 -509 6057 -445
rect 6121 -509 6138 -445
rect 6202 -509 6219 -445
rect 6283 -509 6300 -445
rect 6364 -509 6381 -445
rect 6445 -509 6462 -445
rect 6526 -509 6527 -445
rect 5402 -525 6527 -509
rect 5402 -589 5403 -525
rect 5467 -589 5485 -525
rect 5549 -589 5567 -525
rect 5631 -589 5649 -525
rect 5713 -589 5731 -525
rect 5795 -589 5813 -525
rect 5877 -589 5895 -525
rect 5959 -589 5976 -525
rect 6040 -589 6057 -525
rect 6121 -589 6138 -525
rect 6202 -589 6219 -525
rect 6283 -589 6300 -525
rect 6364 -589 6381 -525
rect 6445 -589 6462 -525
rect 6526 -589 6527 -525
rect 5402 -605 6527 -589
rect 5402 -669 5403 -605
rect 5467 -669 5485 -605
rect 5549 -669 5567 -605
rect 5631 -669 5649 -605
rect 5713 -669 5731 -605
rect 5795 -669 5813 -605
rect 5877 -669 5895 -605
rect 5959 -669 5976 -605
rect 6040 -669 6057 -605
rect 6121 -669 6138 -605
rect 6202 -669 6219 -605
rect 6283 -669 6300 -605
rect 6364 -669 6381 -605
rect 6445 -669 6462 -605
rect 6526 -669 6527 -605
rect 5402 -685 6527 -669
rect 5402 -749 5403 -685
rect 5467 -749 5485 -685
rect 5549 -749 5567 -685
rect 5631 -749 5649 -685
rect 5713 -749 5731 -685
rect 5795 -749 5813 -685
rect 5877 -749 5895 -685
rect 5959 -749 5976 -685
rect 6040 -749 6057 -685
rect 6121 -749 6138 -685
rect 6202 -749 6219 -685
rect 6283 -749 6300 -685
rect 6364 -749 6381 -685
rect 6445 -749 6462 -685
rect 6526 -749 6527 -685
rect 5402 -765 6527 -749
rect 5402 -829 5403 -765
rect 5467 -829 5485 -765
rect 5549 -829 5567 -765
rect 5631 -829 5649 -765
rect 5713 -829 5731 -765
rect 5795 -829 5813 -765
rect 5877 -829 5895 -765
rect 5959 -829 5976 -765
rect 6040 -829 6057 -765
rect 6121 -829 6138 -765
rect 6202 -829 6219 -765
rect 6283 -829 6300 -765
rect 6364 -829 6381 -765
rect 6445 -829 6462 -765
rect 6526 -829 6527 -765
rect 5402 -845 6527 -829
rect 5402 -909 5403 -845
rect 5467 -909 5485 -845
rect 5549 -909 5567 -845
rect 5631 -909 5649 -845
rect 5713 -909 5731 -845
rect 5795 -909 5813 -845
rect 5877 -909 5895 -845
rect 5959 -909 5976 -845
rect 6040 -909 6057 -845
rect 6121 -909 6138 -845
rect 6202 -909 6219 -845
rect 6283 -909 6300 -845
rect 6364 -909 6381 -845
rect 6445 -909 6462 -845
rect 6526 -909 6527 -845
rect 5402 -925 6527 -909
rect 5402 -989 5403 -925
rect 5467 -989 5485 -925
rect 5549 -989 5567 -925
rect 5631 -989 5649 -925
rect 5713 -989 5731 -925
rect 5795 -989 5813 -925
rect 5877 -989 5895 -925
rect 5959 -989 5976 -925
rect 6040 -989 6057 -925
rect 6121 -989 6138 -925
rect 6202 -989 6219 -925
rect 6283 -989 6300 -925
rect 6364 -989 6381 -925
rect 6445 -989 6462 -925
rect 6526 -989 6527 -925
rect 5402 -992 6527 -989
rect 7013 -365 8138 -359
rect 7013 -429 7014 -365
rect 7078 -429 7096 -365
rect 7160 -429 7178 -365
rect 7242 -429 7260 -365
rect 7324 -429 7342 -365
rect 7406 -429 7424 -365
rect 7488 -429 7506 -365
rect 7570 -429 7587 -365
rect 7651 -429 7668 -365
rect 7732 -429 7749 -365
rect 7813 -429 7830 -365
rect 7894 -429 7911 -365
rect 7975 -429 7992 -365
rect 8056 -429 8073 -365
rect 8137 -429 8138 -365
rect 7013 -445 8138 -429
rect 7013 -509 7014 -445
rect 7078 -509 7096 -445
rect 7160 -509 7178 -445
rect 7242 -509 7260 -445
rect 7324 -509 7342 -445
rect 7406 -509 7424 -445
rect 7488 -509 7506 -445
rect 7570 -509 7587 -445
rect 7651 -509 7668 -445
rect 7732 -509 7749 -445
rect 7813 -509 7830 -445
rect 7894 -509 7911 -445
rect 7975 -509 7992 -445
rect 8056 -509 8073 -445
rect 8137 -509 8138 -445
rect 7013 -525 8138 -509
rect 7013 -589 7014 -525
rect 7078 -589 7096 -525
rect 7160 -589 7178 -525
rect 7242 -589 7260 -525
rect 7324 -589 7342 -525
rect 7406 -589 7424 -525
rect 7488 -589 7506 -525
rect 7570 -589 7587 -525
rect 7651 -589 7668 -525
rect 7732 -589 7749 -525
rect 7813 -589 7830 -525
rect 7894 -589 7911 -525
rect 7975 -589 7992 -525
rect 8056 -589 8073 -525
rect 8137 -589 8138 -525
rect 7013 -605 8138 -589
rect 7013 -669 7014 -605
rect 7078 -669 7096 -605
rect 7160 -669 7178 -605
rect 7242 -669 7260 -605
rect 7324 -669 7342 -605
rect 7406 -669 7424 -605
rect 7488 -669 7506 -605
rect 7570 -669 7587 -605
rect 7651 -669 7668 -605
rect 7732 -669 7749 -605
rect 7813 -669 7830 -605
rect 7894 -669 7911 -605
rect 7975 -669 7992 -605
rect 8056 -669 8073 -605
rect 8137 -669 8138 -605
rect 9527 -362 9528 -298
rect 9592 -362 9609 -298
rect 9673 -362 9690 -298
rect 9754 -362 9770 -298
rect 9834 -362 9850 -298
rect 9914 -362 9930 -298
rect 9994 -362 10010 -298
rect 10074 -362 10090 -298
rect 10154 -362 10170 -298
rect 10234 -362 10250 -298
rect 10314 -362 10330 -298
rect 10394 -362 10410 -298
rect 10474 -362 10490 -298
rect 10554 -362 10555 -298
rect 11504 -218 12694 -217
rect 9527 -392 10555 -362
rect 9527 -456 9528 -392
rect 9592 -456 9609 -392
rect 9673 -456 9690 -392
rect 9754 -456 9770 -392
rect 9834 -456 9850 -392
rect 9914 -456 9930 -392
rect 9994 -456 10010 -392
rect 10074 -456 10090 -392
rect 10154 -456 10170 -392
rect 10234 -456 10250 -392
rect 10314 -456 10330 -392
rect 10394 -456 10410 -392
rect 10474 -456 10490 -392
rect 10554 -456 10555 -392
rect 9527 -486 10555 -456
rect 9527 -550 9528 -486
rect 9592 -550 9609 -486
rect 9673 -550 9690 -486
rect 9754 -550 9770 -486
rect 9834 -550 9850 -486
rect 9914 -550 9930 -486
rect 9994 -550 10010 -486
rect 10074 -550 10090 -486
rect 10154 -550 10170 -486
rect 10234 -550 10250 -486
rect 10314 -550 10330 -486
rect 10394 -550 10410 -486
rect 10474 -550 10490 -486
rect 10554 -550 10555 -486
rect 9527 -580 10555 -550
rect 9527 -644 9528 -580
rect 9592 -644 9609 -580
rect 9673 -644 9690 -580
rect 9754 -644 9770 -580
rect 9834 -644 9850 -580
rect 9914 -644 9930 -580
rect 9994 -644 10010 -580
rect 10074 -644 10090 -580
rect 10154 -644 10170 -580
rect 10234 -644 10250 -580
rect 10314 -644 10330 -580
rect 10394 -644 10410 -580
rect 10474 -644 10490 -580
rect 10554 -644 10555 -580
rect 9527 -646 10555 -644
rect 10584 -334 10870 -333
rect 10584 -398 10585 -334
rect 10649 -398 10695 -334
rect 10759 -398 10805 -334
rect 10869 -398 10870 -334
rect 10584 -416 10870 -398
rect 10584 -480 10585 -416
rect 10649 -480 10695 -416
rect 10759 -480 10805 -416
rect 10869 -480 10870 -416
rect 10584 -498 10870 -480
rect 10584 -562 10585 -498
rect 10649 -562 10695 -498
rect 10759 -562 10805 -498
rect 10869 -562 10870 -498
rect 10584 -580 10870 -562
rect 10584 -644 10585 -580
rect 10649 -644 10695 -580
rect 10759 -644 10805 -580
rect 10869 -644 10870 -580
rect 10584 -645 10870 -644
rect 11504 -442 11507 -218
rect 12691 -442 12694 -218
rect 11504 -459 12694 -442
rect 11504 -523 11507 -459
rect 11571 -523 11587 -459
rect 11651 -523 11667 -459
rect 11731 -523 11747 -459
rect 11811 -523 11827 -459
rect 11891 -523 11907 -459
rect 11971 -523 11987 -459
rect 12051 -523 12067 -459
rect 12131 -523 12147 -459
rect 12211 -523 12227 -459
rect 12291 -523 12307 -459
rect 12371 -523 12387 -459
rect 12451 -523 12467 -459
rect 12531 -523 12547 -459
rect 12611 -523 12627 -459
rect 12691 -523 12694 -459
rect 11504 -540 12694 -523
rect 11504 -604 11507 -540
rect 11571 -604 11587 -540
rect 11651 -604 11667 -540
rect 11731 -604 11747 -540
rect 11811 -604 11827 -540
rect 11891 -604 11907 -540
rect 11971 -604 11987 -540
rect 12051 -604 12067 -540
rect 12131 -604 12147 -540
rect 12211 -604 12227 -540
rect 12291 -604 12307 -540
rect 12371 -604 12387 -540
rect 12451 -604 12467 -540
rect 12531 -604 12547 -540
rect 12611 -604 12627 -540
rect 12691 -604 12694 -540
rect 11504 -621 12694 -604
rect 7013 -685 8138 -669
rect 7013 -749 7014 -685
rect 7078 -749 7096 -685
rect 7160 -749 7178 -685
rect 7242 -749 7260 -685
rect 7324 -749 7342 -685
rect 7406 -749 7424 -685
rect 7488 -749 7506 -685
rect 7570 -749 7587 -685
rect 7651 -749 7668 -685
rect 7732 -749 7749 -685
rect 7813 -749 7830 -685
rect 7894 -749 7911 -685
rect 7975 -749 7992 -685
rect 8056 -749 8073 -685
rect 8137 -749 8138 -685
rect 7013 -765 8138 -749
rect 7013 -829 7014 -765
rect 7078 -829 7096 -765
rect 7160 -829 7178 -765
rect 7242 -829 7260 -765
rect 7324 -829 7342 -765
rect 7406 -829 7424 -765
rect 7488 -829 7506 -765
rect 7570 -829 7587 -765
rect 7651 -829 7668 -765
rect 7732 -829 7749 -765
rect 7813 -829 7830 -765
rect 7894 -829 7911 -765
rect 7975 -829 7992 -765
rect 8056 -829 8073 -765
rect 8137 -829 8138 -765
rect 7013 -845 8138 -829
rect 7013 -909 7014 -845
rect 7078 -909 7096 -845
rect 7160 -909 7178 -845
rect 7242 -909 7260 -845
rect 7324 -909 7342 -845
rect 7406 -909 7424 -845
rect 7488 -909 7506 -845
rect 7570 -909 7587 -845
rect 7651 -909 7668 -845
rect 7732 -909 7749 -845
rect 7813 -909 7830 -845
rect 7894 -909 7911 -845
rect 7975 -909 7992 -845
rect 8056 -909 8073 -845
rect 8137 -909 8138 -845
rect 9770 -679 9970 -678
rect 9770 -743 9771 -679
rect 9835 -743 9905 -679
rect 9969 -743 9970 -679
rect 9770 -816 9970 -743
rect 9770 -880 9771 -816
rect 9835 -880 9905 -816
rect 9969 -880 9970 -816
rect 9770 -881 9970 -880
rect 10013 -679 11203 -678
rect 7013 -925 8138 -909
rect 7013 -989 7014 -925
rect 7078 -989 7096 -925
rect 7160 -989 7178 -925
rect 7242 -989 7260 -925
rect 7324 -989 7342 -925
rect 7406 -989 7424 -925
rect 7488 -989 7506 -925
rect 7570 -989 7587 -925
rect 7651 -989 7668 -925
rect 7732 -989 7749 -925
rect 7813 -989 7830 -925
rect 7894 -989 7911 -925
rect 7975 -989 7992 -925
rect 8056 -989 8073 -925
rect 8137 -989 8138 -925
rect 7013 -992 8138 -989
rect 10013 -903 10016 -679
rect 11200 -903 11203 -679
rect 10013 -920 11203 -903
rect 10013 -984 10016 -920
rect 10080 -984 10096 -920
rect 10160 -984 10176 -920
rect 10240 -984 10256 -920
rect 10320 -984 10336 -920
rect 10400 -984 10416 -920
rect 10480 -984 10496 -920
rect 10560 -984 10576 -920
rect 10640 -984 10656 -920
rect 10720 -984 10736 -920
rect 10800 -984 10816 -920
rect 10880 -984 10896 -920
rect 10960 -984 10976 -920
rect 11040 -984 11056 -920
rect 11120 -984 11136 -920
rect 11200 -984 11203 -920
rect 10013 -1001 11203 -984
rect 10013 -1065 10016 -1001
rect 10080 -1065 10096 -1001
rect 10160 -1065 10176 -1001
rect 10240 -1065 10256 -1001
rect 10320 -1065 10336 -1001
rect 10400 -1065 10416 -1001
rect 10480 -1065 10496 -1001
rect 10560 -1065 10576 -1001
rect 10640 -1065 10656 -1001
rect 10720 -1065 10736 -1001
rect 10800 -1065 10816 -1001
rect 10880 -1065 10896 -1001
rect 10960 -1065 10976 -1001
rect 11040 -1065 11056 -1001
rect 11120 -1065 11136 -1001
rect 11200 -1065 11203 -1001
rect 10013 -1082 11203 -1065
rect 10013 -1146 10016 -1082
rect 10080 -1146 10096 -1082
rect 10160 -1146 10176 -1082
rect 10240 -1146 10256 -1082
rect 10320 -1146 10336 -1082
rect 10400 -1146 10416 -1082
rect 10480 -1146 10496 -1082
rect 10560 -1146 10576 -1082
rect 10640 -1146 10656 -1082
rect 10720 -1146 10736 -1082
rect 10800 -1146 10816 -1082
rect 10880 -1146 10896 -1082
rect 10960 -1146 10976 -1082
rect 11040 -1146 11056 -1082
rect 11120 -1146 11136 -1082
rect 11200 -1146 11203 -1082
rect 10013 -1163 11203 -1146
rect 10013 -1227 10016 -1163
rect 10080 -1227 10096 -1163
rect 10160 -1227 10176 -1163
rect 10240 -1227 10256 -1163
rect 10320 -1227 10336 -1163
rect 10400 -1227 10416 -1163
rect 10480 -1227 10496 -1163
rect 10560 -1227 10576 -1163
rect 10640 -1227 10656 -1163
rect 10720 -1227 10736 -1163
rect 10800 -1227 10816 -1163
rect 10880 -1227 10896 -1163
rect 10960 -1227 10976 -1163
rect 11040 -1227 11056 -1163
rect 11120 -1227 11136 -1163
rect 11200 -1227 11203 -1163
rect 10013 -1244 11203 -1227
rect 10013 -1308 10016 -1244
rect 10080 -1308 10096 -1244
rect 10160 -1308 10176 -1244
rect 10240 -1308 10256 -1244
rect 10320 -1308 10336 -1244
rect 10400 -1308 10416 -1244
rect 10480 -1308 10496 -1244
rect 10560 -1308 10576 -1244
rect 10640 -1308 10656 -1244
rect 10720 -1308 10736 -1244
rect 10800 -1308 10816 -1244
rect 10880 -1308 10896 -1244
rect 10960 -1308 10976 -1244
rect 11040 -1308 11056 -1244
rect 11120 -1308 11136 -1244
rect 11200 -1308 11203 -1244
rect 10013 -1325 11203 -1308
rect 10013 -1389 10016 -1325
rect 10080 -1389 10096 -1325
rect 10160 -1389 10176 -1325
rect 10240 -1389 10256 -1325
rect 10320 -1389 10336 -1325
rect 10400 -1389 10416 -1325
rect 10480 -1389 10496 -1325
rect 10560 -1389 10576 -1325
rect 10640 -1389 10656 -1325
rect 10720 -1389 10736 -1325
rect 10800 -1389 10816 -1325
rect 10880 -1389 10896 -1325
rect 10960 -1389 10976 -1325
rect 11040 -1389 11056 -1325
rect 11120 -1389 11136 -1325
rect 11200 -1389 11203 -1325
rect 10013 -1406 11203 -1389
rect 10013 -1470 10016 -1406
rect 10080 -1470 10096 -1406
rect 10160 -1470 10176 -1406
rect 10240 -1470 10256 -1406
rect 10320 -1470 10336 -1406
rect 10400 -1470 10416 -1406
rect 10480 -1470 10496 -1406
rect 10560 -1470 10576 -1406
rect 10640 -1470 10656 -1406
rect 10720 -1470 10736 -1406
rect 10800 -1470 10816 -1406
rect 10880 -1470 10896 -1406
rect 10960 -1470 10976 -1406
rect 11040 -1470 11056 -1406
rect 11120 -1470 11136 -1406
rect 11200 -1470 11203 -1406
rect 10013 -1487 11203 -1470
rect 10013 -1551 10016 -1487
rect 10080 -1551 10096 -1487
rect 10160 -1551 10176 -1487
rect 10240 -1551 10256 -1487
rect 10320 -1551 10336 -1487
rect 10400 -1551 10416 -1487
rect 10480 -1551 10496 -1487
rect 10560 -1551 10576 -1487
rect 10640 -1551 10656 -1487
rect 10720 -1551 10736 -1487
rect 10800 -1551 10816 -1487
rect 10880 -1551 10896 -1487
rect 10960 -1551 10976 -1487
rect 11040 -1551 11056 -1487
rect 11120 -1551 11136 -1487
rect 11200 -1551 11203 -1487
rect 10013 -1568 11203 -1551
rect 10013 -1632 10016 -1568
rect 10080 -1632 10096 -1568
rect 10160 -1632 10176 -1568
rect 10240 -1632 10256 -1568
rect 10320 -1632 10336 -1568
rect 10400 -1632 10416 -1568
rect 10480 -1632 10496 -1568
rect 10560 -1632 10576 -1568
rect 10640 -1632 10656 -1568
rect 10720 -1632 10736 -1568
rect 10800 -1632 10816 -1568
rect 10880 -1632 10896 -1568
rect 10960 -1632 10976 -1568
rect 11040 -1632 11056 -1568
rect 11120 -1632 11136 -1568
rect 11200 -1632 11203 -1568
rect 10013 -1649 11203 -1632
rect 10013 -1713 10016 -1649
rect 10080 -1713 10096 -1649
rect 10160 -1713 10176 -1649
rect 10240 -1713 10256 -1649
rect 10320 -1713 10336 -1649
rect 10400 -1713 10416 -1649
rect 10480 -1713 10496 -1649
rect 10560 -1713 10576 -1649
rect 10640 -1713 10656 -1649
rect 10720 -1713 10736 -1649
rect 10800 -1713 10816 -1649
rect 10880 -1713 10896 -1649
rect 10960 -1713 10976 -1649
rect 11040 -1713 11056 -1649
rect 11120 -1713 11136 -1649
rect 11200 -1713 11203 -1649
rect 10013 -1730 11203 -1713
rect 10013 -1794 10016 -1730
rect 10080 -1794 10096 -1730
rect 10160 -1794 10176 -1730
rect 10240 -1794 10256 -1730
rect 10320 -1794 10336 -1730
rect 10400 -1794 10416 -1730
rect 10480 -1794 10496 -1730
rect 10560 -1794 10576 -1730
rect 10640 -1794 10656 -1730
rect 10720 -1794 10736 -1730
rect 10800 -1794 10816 -1730
rect 10880 -1794 10896 -1730
rect 10960 -1794 10976 -1730
rect 11040 -1794 11056 -1730
rect 11120 -1794 11136 -1730
rect 11200 -1794 11203 -1730
rect 10013 -1811 11203 -1794
rect 10013 -1875 10016 -1811
rect 10080 -1875 10096 -1811
rect 10160 -1875 10176 -1811
rect 10240 -1875 10256 -1811
rect 10320 -1875 10336 -1811
rect 10400 -1875 10416 -1811
rect 10480 -1875 10496 -1811
rect 10560 -1875 10576 -1811
rect 10640 -1875 10656 -1811
rect 10720 -1875 10736 -1811
rect 10800 -1875 10816 -1811
rect 10880 -1875 10896 -1811
rect 10960 -1875 10976 -1811
rect 11040 -1875 11056 -1811
rect 11120 -1875 11136 -1811
rect 11200 -1875 11203 -1811
rect 10013 -1892 11203 -1875
rect 10013 -1956 10016 -1892
rect 10080 -1956 10096 -1892
rect 10160 -1956 10176 -1892
rect 10240 -1956 10256 -1892
rect 10320 -1956 10336 -1892
rect 10400 -1956 10416 -1892
rect 10480 -1956 10496 -1892
rect 10560 -1956 10576 -1892
rect 10640 -1956 10656 -1892
rect 10720 -1956 10736 -1892
rect 10800 -1956 10816 -1892
rect 10880 -1956 10896 -1892
rect 10960 -1956 10976 -1892
rect 11040 -1956 11056 -1892
rect 11120 -1956 11136 -1892
rect 11200 -1956 11203 -1892
rect 10013 -1973 11203 -1956
rect 10013 -2037 10016 -1973
rect 10080 -2037 10096 -1973
rect 10160 -2037 10176 -1973
rect 10240 -2037 10256 -1973
rect 10320 -2037 10336 -1973
rect 10400 -2037 10416 -1973
rect 10480 -2037 10496 -1973
rect 10560 -2037 10576 -1973
rect 10640 -2037 10656 -1973
rect 10720 -2037 10736 -1973
rect 10800 -2037 10816 -1973
rect 10880 -2037 10896 -1973
rect 10960 -2037 10976 -1973
rect 11040 -2037 11056 -1973
rect 11120 -2037 11136 -1973
rect 11200 -2037 11203 -1973
rect 10013 -2054 11203 -2037
rect 10013 -2118 10016 -2054
rect 10080 -2118 10096 -2054
rect 10160 -2118 10176 -2054
rect 10240 -2118 10256 -2054
rect 10320 -2118 10336 -2054
rect 10400 -2118 10416 -2054
rect 10480 -2118 10496 -2054
rect 10560 -2118 10576 -2054
rect 10640 -2118 10656 -2054
rect 10720 -2118 10736 -2054
rect 10800 -2118 10816 -2054
rect 10880 -2118 10896 -2054
rect 10960 -2118 10976 -2054
rect 11040 -2118 11056 -2054
rect 11120 -2118 11136 -2054
rect 11200 -2118 11203 -2054
rect 10013 -2135 11203 -2118
rect 10013 -2199 10016 -2135
rect 10080 -2199 10096 -2135
rect 10160 -2199 10176 -2135
rect 10240 -2199 10256 -2135
rect 10320 -2199 10336 -2135
rect 10400 -2199 10416 -2135
rect 10480 -2199 10496 -2135
rect 10560 -2199 10576 -2135
rect 10640 -2199 10656 -2135
rect 10720 -2199 10736 -2135
rect 10800 -2199 10816 -2135
rect 10880 -2199 10896 -2135
rect 10960 -2199 10976 -2135
rect 11040 -2199 11056 -2135
rect 11120 -2199 11136 -2135
rect 11200 -2199 11203 -2135
rect 10013 -2216 11203 -2199
rect 10013 -2280 10016 -2216
rect 10080 -2280 10096 -2216
rect 10160 -2280 10176 -2216
rect 10240 -2280 10256 -2216
rect 10320 -2280 10336 -2216
rect 10400 -2280 10416 -2216
rect 10480 -2280 10496 -2216
rect 10560 -2280 10576 -2216
rect 10640 -2280 10656 -2216
rect 10720 -2280 10736 -2216
rect 10800 -2280 10816 -2216
rect 10880 -2280 10896 -2216
rect 10960 -2280 10976 -2216
rect 11040 -2280 11056 -2216
rect 11120 -2280 11136 -2216
rect 11200 -2280 11203 -2216
rect 10013 -2297 11203 -2280
rect 10013 -2361 10016 -2297
rect 10080 -2361 10096 -2297
rect 10160 -2361 10176 -2297
rect 10240 -2361 10256 -2297
rect 10320 -2361 10336 -2297
rect 10400 -2361 10416 -2297
rect 10480 -2361 10496 -2297
rect 10560 -2361 10576 -2297
rect 10640 -2361 10656 -2297
rect 10720 -2361 10736 -2297
rect 10800 -2361 10816 -2297
rect 10880 -2361 10896 -2297
rect 10960 -2361 10976 -2297
rect 11040 -2361 11056 -2297
rect 11120 -2361 11136 -2297
rect 11200 -2361 11203 -2297
rect 10013 -2378 11203 -2361
rect 10013 -2442 10016 -2378
rect 10080 -2442 10096 -2378
rect 10160 -2442 10176 -2378
rect 10240 -2442 10256 -2378
rect 10320 -2442 10336 -2378
rect 10400 -2442 10416 -2378
rect 10480 -2442 10496 -2378
rect 10560 -2442 10576 -2378
rect 10640 -2442 10656 -2378
rect 10720 -2442 10736 -2378
rect 10800 -2442 10816 -2378
rect 10880 -2442 10896 -2378
rect 10960 -2442 10976 -2378
rect 11040 -2442 11056 -2378
rect 11120 -2442 11136 -2378
rect 11200 -2442 11203 -2378
rect 10013 -2459 11203 -2442
rect 10013 -2523 10016 -2459
rect 10080 -2523 10096 -2459
rect 10160 -2523 10176 -2459
rect 10240 -2523 10256 -2459
rect 10320 -2523 10336 -2459
rect 10400 -2523 10416 -2459
rect 10480 -2523 10496 -2459
rect 10560 -2523 10576 -2459
rect 10640 -2523 10656 -2459
rect 10720 -2523 10736 -2459
rect 10800 -2523 10816 -2459
rect 10880 -2523 10896 -2459
rect 10960 -2523 10976 -2459
rect 11040 -2523 11056 -2459
rect 11120 -2523 11136 -2459
rect 11200 -2523 11203 -2459
rect 10013 -2540 11203 -2523
rect 10013 -2604 10016 -2540
rect 10080 -2604 10096 -2540
rect 10160 -2604 10176 -2540
rect 10240 -2604 10256 -2540
rect 10320 -2604 10336 -2540
rect 10400 -2604 10416 -2540
rect 10480 -2604 10496 -2540
rect 10560 -2604 10576 -2540
rect 10640 -2604 10656 -2540
rect 10720 -2604 10736 -2540
rect 10800 -2604 10816 -2540
rect 10880 -2604 10896 -2540
rect 10960 -2604 10976 -2540
rect 11040 -2604 11056 -2540
rect 11120 -2604 11136 -2540
rect 11200 -2604 11203 -2540
rect 10013 -2621 11203 -2604
rect 10013 -2685 10016 -2621
rect 10080 -2685 10096 -2621
rect 10160 -2685 10176 -2621
rect 10240 -2685 10256 -2621
rect 10320 -2685 10336 -2621
rect 10400 -2685 10416 -2621
rect 10480 -2685 10496 -2621
rect 10560 -2685 10576 -2621
rect 10640 -2685 10656 -2621
rect 10720 -2685 10736 -2621
rect 10800 -2685 10816 -2621
rect 10880 -2685 10896 -2621
rect 10960 -2685 10976 -2621
rect 11040 -2685 11056 -2621
rect 11120 -2685 11136 -2621
rect 11200 -2685 11203 -2621
rect 10013 -2702 11203 -2685
rect 10013 -2766 10016 -2702
rect 10080 -2766 10096 -2702
rect 10160 -2766 10176 -2702
rect 10240 -2766 10256 -2702
rect 10320 -2766 10336 -2702
rect 10400 -2766 10416 -2702
rect 10480 -2766 10496 -2702
rect 10560 -2766 10576 -2702
rect 10640 -2766 10656 -2702
rect 10720 -2766 10736 -2702
rect 10800 -2766 10816 -2702
rect 10880 -2766 10896 -2702
rect 10960 -2766 10976 -2702
rect 11040 -2766 11056 -2702
rect 11120 -2766 11136 -2702
rect 11200 -2766 11203 -2702
rect 10013 -2783 11203 -2766
rect 10013 -2847 10016 -2783
rect 10080 -2847 10096 -2783
rect 10160 -2847 10176 -2783
rect 10240 -2847 10256 -2783
rect 10320 -2847 10336 -2783
rect 10400 -2847 10416 -2783
rect 10480 -2847 10496 -2783
rect 10560 -2847 10576 -2783
rect 10640 -2847 10656 -2783
rect 10720 -2847 10736 -2783
rect 10800 -2847 10816 -2783
rect 10880 -2847 10896 -2783
rect 10960 -2847 10976 -2783
rect 11040 -2847 11056 -2783
rect 11120 -2847 11136 -2783
rect 11200 -2847 11203 -2783
rect 10013 -2864 11203 -2847
rect 10013 -2928 10016 -2864
rect 10080 -2928 10096 -2864
rect 10160 -2928 10176 -2864
rect 10240 -2928 10256 -2864
rect 10320 -2928 10336 -2864
rect 10400 -2928 10416 -2864
rect 10480 -2928 10496 -2864
rect 10560 -2928 10576 -2864
rect 10640 -2928 10656 -2864
rect 10720 -2928 10736 -2864
rect 10800 -2928 10816 -2864
rect 10880 -2928 10896 -2864
rect 10960 -2928 10976 -2864
rect 11040 -2928 11056 -2864
rect 11120 -2928 11136 -2864
rect 11200 -2928 11203 -2864
rect 10013 -2945 11203 -2928
rect 10013 -3009 10016 -2945
rect 10080 -3009 10096 -2945
rect 10160 -3009 10176 -2945
rect 10240 -3009 10256 -2945
rect 10320 -3009 10336 -2945
rect 10400 -3009 10416 -2945
rect 10480 -3009 10496 -2945
rect 10560 -3009 10576 -2945
rect 10640 -3009 10656 -2945
rect 10720 -3009 10736 -2945
rect 10800 -3009 10816 -2945
rect 10880 -3009 10896 -2945
rect 10960 -3009 10976 -2945
rect 11040 -3009 11056 -2945
rect 11120 -3009 11136 -2945
rect 11200 -3009 11203 -2945
rect 10013 -3026 11203 -3009
rect 10013 -3090 10016 -3026
rect 10080 -3090 10096 -3026
rect 10160 -3090 10176 -3026
rect 10240 -3090 10256 -3026
rect 10320 -3090 10336 -3026
rect 10400 -3090 10416 -3026
rect 10480 -3090 10496 -3026
rect 10560 -3090 10576 -3026
rect 10640 -3090 10656 -3026
rect 10720 -3090 10736 -3026
rect 10800 -3090 10816 -3026
rect 10880 -3090 10896 -3026
rect 10960 -3090 10976 -3026
rect 11040 -3090 11056 -3026
rect 11120 -3090 11136 -3026
rect 11200 -3090 11203 -3026
rect 10013 -3107 11203 -3090
rect 10013 -3171 10016 -3107
rect 10080 -3171 10096 -3107
rect 10160 -3171 10176 -3107
rect 10240 -3171 10256 -3107
rect 10320 -3171 10336 -3107
rect 10400 -3171 10416 -3107
rect 10480 -3171 10496 -3107
rect 10560 -3171 10576 -3107
rect 10640 -3171 10656 -3107
rect 10720 -3171 10736 -3107
rect 10800 -3171 10816 -3107
rect 10880 -3171 10896 -3107
rect 10960 -3171 10976 -3107
rect 11040 -3171 11056 -3107
rect 11120 -3171 11136 -3107
rect 11200 -3171 11203 -3107
rect 10013 -3188 11203 -3171
rect 10013 -3252 10016 -3188
rect 10080 -3252 10096 -3188
rect 10160 -3252 10176 -3188
rect 10240 -3252 10256 -3188
rect 10320 -3252 10336 -3188
rect 10400 -3252 10416 -3188
rect 10480 -3252 10496 -3188
rect 10560 -3252 10576 -3188
rect 10640 -3252 10656 -3188
rect 10720 -3252 10736 -3188
rect 10800 -3252 10816 -3188
rect 10880 -3252 10896 -3188
rect 10960 -3252 10976 -3188
rect 11040 -3252 11056 -3188
rect 11120 -3252 11136 -3188
rect 11200 -3252 11203 -3188
rect 10013 -3269 11203 -3252
rect 10013 -3333 10016 -3269
rect 10080 -3333 10096 -3269
rect 10160 -3333 10176 -3269
rect 10240 -3333 10256 -3269
rect 10320 -3333 10336 -3269
rect 10400 -3333 10416 -3269
rect 10480 -3333 10496 -3269
rect 10560 -3333 10576 -3269
rect 10640 -3333 10656 -3269
rect 10720 -3333 10736 -3269
rect 10800 -3333 10816 -3269
rect 10880 -3333 10896 -3269
rect 10960 -3333 10976 -3269
rect 11040 -3333 11056 -3269
rect 11120 -3333 11136 -3269
rect 11200 -3333 11203 -3269
rect 10013 -3350 11203 -3333
rect 10013 -3414 10016 -3350
rect 10080 -3414 10096 -3350
rect 10160 -3414 10176 -3350
rect 10240 -3414 10256 -3350
rect 10320 -3414 10336 -3350
rect 10400 -3414 10416 -3350
rect 10480 -3414 10496 -3350
rect 10560 -3414 10576 -3350
rect 10640 -3414 10656 -3350
rect 10720 -3414 10736 -3350
rect 10800 -3414 10816 -3350
rect 10880 -3414 10896 -3350
rect 10960 -3414 10976 -3350
rect 11040 -3414 11056 -3350
rect 11120 -3414 11136 -3350
rect 11200 -3414 11203 -3350
rect 10013 -3415 11203 -3414
rect 11504 -685 11507 -621
rect 11571 -685 11587 -621
rect 11651 -685 11667 -621
rect 11731 -685 11747 -621
rect 11811 -685 11827 -621
rect 11891 -685 11907 -621
rect 11971 -685 11987 -621
rect 12051 -685 12067 -621
rect 12131 -685 12147 -621
rect 12211 -685 12227 -621
rect 12291 -685 12307 -621
rect 12371 -685 12387 -621
rect 12451 -685 12467 -621
rect 12531 -685 12547 -621
rect 12611 -685 12627 -621
rect 12691 -685 12694 -621
rect 11504 -702 12694 -685
rect 11504 -766 11507 -702
rect 11571 -766 11587 -702
rect 11651 -766 11667 -702
rect 11731 -766 11747 -702
rect 11811 -766 11827 -702
rect 11891 -766 11907 -702
rect 11971 -766 11987 -702
rect 12051 -766 12067 -702
rect 12131 -766 12147 -702
rect 12211 -766 12227 -702
rect 12291 -766 12307 -702
rect 12371 -766 12387 -702
rect 12451 -766 12467 -702
rect 12531 -766 12547 -702
rect 12611 -766 12627 -702
rect 12691 -766 12694 -702
rect 11504 -783 12694 -766
rect 11504 -847 11507 -783
rect 11571 -847 11587 -783
rect 11651 -847 11667 -783
rect 11731 -847 11747 -783
rect 11811 -847 11827 -783
rect 11891 -847 11907 -783
rect 11971 -847 11987 -783
rect 12051 -847 12067 -783
rect 12131 -847 12147 -783
rect 12211 -847 12227 -783
rect 12291 -847 12307 -783
rect 12371 -847 12387 -783
rect 12451 -847 12467 -783
rect 12531 -847 12547 -783
rect 12611 -847 12627 -783
rect 12691 -847 12694 -783
rect 11504 -864 12694 -847
rect 11504 -928 11507 -864
rect 11571 -928 11587 -864
rect 11651 -928 11667 -864
rect 11731 -928 11747 -864
rect 11811 -928 11827 -864
rect 11891 -928 11907 -864
rect 11971 -928 11987 -864
rect 12051 -928 12067 -864
rect 12131 -928 12147 -864
rect 12211 -928 12227 -864
rect 12291 -928 12307 -864
rect 12371 -928 12387 -864
rect 12451 -928 12467 -864
rect 12531 -928 12547 -864
rect 12611 -928 12627 -864
rect 12691 -928 12694 -864
rect 11504 -945 12694 -928
rect 11504 -1009 11507 -945
rect 11571 -1009 11587 -945
rect 11651 -1009 11667 -945
rect 11731 -1009 11747 -945
rect 11811 -1009 11827 -945
rect 11891 -1009 11907 -945
rect 11971 -1009 11987 -945
rect 12051 -1009 12067 -945
rect 12131 -1009 12147 -945
rect 12211 -1009 12227 -945
rect 12291 -1009 12307 -945
rect 12371 -1009 12387 -945
rect 12451 -1009 12467 -945
rect 12531 -1009 12547 -945
rect 12611 -1009 12627 -945
rect 12691 -1009 12694 -945
rect 11504 -1026 12694 -1009
rect 11504 -1090 11507 -1026
rect 11571 -1090 11587 -1026
rect 11651 -1090 11667 -1026
rect 11731 -1090 11747 -1026
rect 11811 -1090 11827 -1026
rect 11891 -1090 11907 -1026
rect 11971 -1090 11987 -1026
rect 12051 -1090 12067 -1026
rect 12131 -1090 12147 -1026
rect 12211 -1090 12227 -1026
rect 12291 -1090 12307 -1026
rect 12371 -1090 12387 -1026
rect 12451 -1090 12467 -1026
rect 12531 -1090 12547 -1026
rect 12611 -1090 12627 -1026
rect 12691 -1090 12694 -1026
rect 11504 -1107 12694 -1090
rect 11504 -1171 11507 -1107
rect 11571 -1171 11587 -1107
rect 11651 -1171 11667 -1107
rect 11731 -1171 11747 -1107
rect 11811 -1171 11827 -1107
rect 11891 -1171 11907 -1107
rect 11971 -1171 11987 -1107
rect 12051 -1171 12067 -1107
rect 12131 -1171 12147 -1107
rect 12211 -1171 12227 -1107
rect 12291 -1171 12307 -1107
rect 12371 -1171 12387 -1107
rect 12451 -1171 12467 -1107
rect 12531 -1171 12547 -1107
rect 12611 -1171 12627 -1107
rect 12691 -1171 12694 -1107
rect 11504 -1188 12694 -1171
rect 11504 -1252 11507 -1188
rect 11571 -1252 11587 -1188
rect 11651 -1252 11667 -1188
rect 11731 -1252 11747 -1188
rect 11811 -1252 11827 -1188
rect 11891 -1252 11907 -1188
rect 11971 -1252 11987 -1188
rect 12051 -1252 12067 -1188
rect 12131 -1252 12147 -1188
rect 12211 -1252 12227 -1188
rect 12291 -1252 12307 -1188
rect 12371 -1252 12387 -1188
rect 12451 -1252 12467 -1188
rect 12531 -1252 12547 -1188
rect 12611 -1252 12627 -1188
rect 12691 -1252 12694 -1188
rect 11504 -1269 12694 -1252
rect 11504 -1333 11507 -1269
rect 11571 -1333 11587 -1269
rect 11651 -1333 11667 -1269
rect 11731 -1333 11747 -1269
rect 11811 -1333 11827 -1269
rect 11891 -1333 11907 -1269
rect 11971 -1333 11987 -1269
rect 12051 -1333 12067 -1269
rect 12131 -1333 12147 -1269
rect 12211 -1333 12227 -1269
rect 12291 -1333 12307 -1269
rect 12371 -1333 12387 -1269
rect 12451 -1333 12467 -1269
rect 12531 -1333 12547 -1269
rect 12611 -1333 12627 -1269
rect 12691 -1333 12694 -1269
rect 11504 -1350 12694 -1333
rect 11504 -1414 11507 -1350
rect 11571 -1414 11587 -1350
rect 11651 -1414 11667 -1350
rect 11731 -1414 11747 -1350
rect 11811 -1414 11827 -1350
rect 11891 -1414 11907 -1350
rect 11971 -1414 11987 -1350
rect 12051 -1414 12067 -1350
rect 12131 -1414 12147 -1350
rect 12211 -1414 12227 -1350
rect 12291 -1414 12307 -1350
rect 12371 -1414 12387 -1350
rect 12451 -1414 12467 -1350
rect 12531 -1414 12547 -1350
rect 12611 -1414 12627 -1350
rect 12691 -1414 12694 -1350
rect 11504 -1431 12694 -1414
rect 11504 -1495 11507 -1431
rect 11571 -1495 11587 -1431
rect 11651 -1495 11667 -1431
rect 11731 -1495 11747 -1431
rect 11811 -1495 11827 -1431
rect 11891 -1495 11907 -1431
rect 11971 -1495 11987 -1431
rect 12051 -1495 12067 -1431
rect 12131 -1495 12147 -1431
rect 12211 -1495 12227 -1431
rect 12291 -1495 12307 -1431
rect 12371 -1495 12387 -1431
rect 12451 -1495 12467 -1431
rect 12531 -1495 12547 -1431
rect 12611 -1495 12627 -1431
rect 12691 -1495 12694 -1431
rect 11504 -1512 12694 -1495
rect 11504 -1576 11507 -1512
rect 11571 -1576 11587 -1512
rect 11651 -1576 11667 -1512
rect 11731 -1576 11747 -1512
rect 11811 -1576 11827 -1512
rect 11891 -1576 11907 -1512
rect 11971 -1576 11987 -1512
rect 12051 -1576 12067 -1512
rect 12131 -1576 12147 -1512
rect 12211 -1576 12227 -1512
rect 12291 -1576 12307 -1512
rect 12371 -1576 12387 -1512
rect 12451 -1576 12467 -1512
rect 12531 -1576 12547 -1512
rect 12611 -1576 12627 -1512
rect 12691 -1576 12694 -1512
rect 11504 -1593 12694 -1576
rect 11504 -1657 11507 -1593
rect 11571 -1657 11587 -1593
rect 11651 -1657 11667 -1593
rect 11731 -1657 11747 -1593
rect 11811 -1657 11827 -1593
rect 11891 -1657 11907 -1593
rect 11971 -1657 11987 -1593
rect 12051 -1657 12067 -1593
rect 12131 -1657 12147 -1593
rect 12211 -1657 12227 -1593
rect 12291 -1657 12307 -1593
rect 12371 -1657 12387 -1593
rect 12451 -1657 12467 -1593
rect 12531 -1657 12547 -1593
rect 12611 -1657 12627 -1593
rect 12691 -1657 12694 -1593
rect 11504 -1674 12694 -1657
rect 11504 -1738 11507 -1674
rect 11571 -1738 11587 -1674
rect 11651 -1738 11667 -1674
rect 11731 -1738 11747 -1674
rect 11811 -1738 11827 -1674
rect 11891 -1738 11907 -1674
rect 11971 -1738 11987 -1674
rect 12051 -1738 12067 -1674
rect 12131 -1738 12147 -1674
rect 12211 -1738 12227 -1674
rect 12291 -1738 12307 -1674
rect 12371 -1738 12387 -1674
rect 12451 -1738 12467 -1674
rect 12531 -1738 12547 -1674
rect 12611 -1738 12627 -1674
rect 12691 -1738 12694 -1674
rect 11504 -1755 12694 -1738
rect 11504 -1819 11507 -1755
rect 11571 -1819 11587 -1755
rect 11651 -1819 11667 -1755
rect 11731 -1819 11747 -1755
rect 11811 -1819 11827 -1755
rect 11891 -1819 11907 -1755
rect 11971 -1819 11987 -1755
rect 12051 -1819 12067 -1755
rect 12131 -1819 12147 -1755
rect 12211 -1819 12227 -1755
rect 12291 -1819 12307 -1755
rect 12371 -1819 12387 -1755
rect 12451 -1819 12467 -1755
rect 12531 -1819 12547 -1755
rect 12611 -1819 12627 -1755
rect 12691 -1819 12694 -1755
rect 11504 -1836 12694 -1819
rect 11504 -1900 11507 -1836
rect 11571 -1900 11587 -1836
rect 11651 -1900 11667 -1836
rect 11731 -1900 11747 -1836
rect 11811 -1900 11827 -1836
rect 11891 -1900 11907 -1836
rect 11971 -1900 11987 -1836
rect 12051 -1900 12067 -1836
rect 12131 -1900 12147 -1836
rect 12211 -1900 12227 -1836
rect 12291 -1900 12307 -1836
rect 12371 -1900 12387 -1836
rect 12451 -1900 12467 -1836
rect 12531 -1900 12547 -1836
rect 12611 -1900 12627 -1836
rect 12691 -1900 12694 -1836
rect 11504 -1917 12694 -1900
rect 11504 -1981 11507 -1917
rect 11571 -1981 11587 -1917
rect 11651 -1981 11667 -1917
rect 11731 -1981 11747 -1917
rect 11811 -1981 11827 -1917
rect 11891 -1981 11907 -1917
rect 11971 -1981 11987 -1917
rect 12051 -1981 12067 -1917
rect 12131 -1981 12147 -1917
rect 12211 -1981 12227 -1917
rect 12291 -1981 12307 -1917
rect 12371 -1981 12387 -1917
rect 12451 -1981 12467 -1917
rect 12531 -1981 12547 -1917
rect 12611 -1981 12627 -1917
rect 12691 -1981 12694 -1917
rect 11504 -1998 12694 -1981
rect 11504 -2062 11507 -1998
rect 11571 -2062 11587 -1998
rect 11651 -2062 11667 -1998
rect 11731 -2062 11747 -1998
rect 11811 -2062 11827 -1998
rect 11891 -2062 11907 -1998
rect 11971 -2062 11987 -1998
rect 12051 -2062 12067 -1998
rect 12131 -2062 12147 -1998
rect 12211 -2062 12227 -1998
rect 12291 -2062 12307 -1998
rect 12371 -2062 12387 -1998
rect 12451 -2062 12467 -1998
rect 12531 -2062 12547 -1998
rect 12611 -2062 12627 -1998
rect 12691 -2062 12694 -1998
rect 11504 -2079 12694 -2062
rect 11504 -2143 11507 -2079
rect 11571 -2143 11587 -2079
rect 11651 -2143 11667 -2079
rect 11731 -2143 11747 -2079
rect 11811 -2143 11827 -2079
rect 11891 -2143 11907 -2079
rect 11971 -2143 11987 -2079
rect 12051 -2143 12067 -2079
rect 12131 -2143 12147 -2079
rect 12211 -2143 12227 -2079
rect 12291 -2143 12307 -2079
rect 12371 -2143 12387 -2079
rect 12451 -2143 12467 -2079
rect 12531 -2143 12547 -2079
rect 12611 -2143 12627 -2079
rect 12691 -2143 12694 -2079
rect 11504 -2160 12694 -2143
rect 11504 -2224 11507 -2160
rect 11571 -2224 11587 -2160
rect 11651 -2224 11667 -2160
rect 11731 -2224 11747 -2160
rect 11811 -2224 11827 -2160
rect 11891 -2224 11907 -2160
rect 11971 -2224 11987 -2160
rect 12051 -2224 12067 -2160
rect 12131 -2224 12147 -2160
rect 12211 -2224 12227 -2160
rect 12291 -2224 12307 -2160
rect 12371 -2224 12387 -2160
rect 12451 -2224 12467 -2160
rect 12531 -2224 12547 -2160
rect 12611 -2224 12627 -2160
rect 12691 -2224 12694 -2160
rect 11504 -2241 12694 -2224
rect 11504 -2305 11507 -2241
rect 11571 -2305 11587 -2241
rect 11651 -2305 11667 -2241
rect 11731 -2305 11747 -2241
rect 11811 -2305 11827 -2241
rect 11891 -2305 11907 -2241
rect 11971 -2305 11987 -2241
rect 12051 -2305 12067 -2241
rect 12131 -2305 12147 -2241
rect 12211 -2305 12227 -2241
rect 12291 -2305 12307 -2241
rect 12371 -2305 12387 -2241
rect 12451 -2305 12467 -2241
rect 12531 -2305 12547 -2241
rect 12611 -2305 12627 -2241
rect 12691 -2305 12694 -2241
rect 11504 -2322 12694 -2305
rect 11504 -2386 11507 -2322
rect 11571 -2386 11587 -2322
rect 11651 -2386 11667 -2322
rect 11731 -2386 11747 -2322
rect 11811 -2386 11827 -2322
rect 11891 -2386 11907 -2322
rect 11971 -2386 11987 -2322
rect 12051 -2386 12067 -2322
rect 12131 -2386 12147 -2322
rect 12211 -2386 12227 -2322
rect 12291 -2386 12307 -2322
rect 12371 -2386 12387 -2322
rect 12451 -2386 12467 -2322
rect 12531 -2386 12547 -2322
rect 12611 -2386 12627 -2322
rect 12691 -2386 12694 -2322
rect 11504 -2403 12694 -2386
rect 11504 -2467 11507 -2403
rect 11571 -2467 11587 -2403
rect 11651 -2467 11667 -2403
rect 11731 -2467 11747 -2403
rect 11811 -2467 11827 -2403
rect 11891 -2467 11907 -2403
rect 11971 -2467 11987 -2403
rect 12051 -2467 12067 -2403
rect 12131 -2467 12147 -2403
rect 12211 -2467 12227 -2403
rect 12291 -2467 12307 -2403
rect 12371 -2467 12387 -2403
rect 12451 -2467 12467 -2403
rect 12531 -2467 12547 -2403
rect 12611 -2467 12627 -2403
rect 12691 -2467 12694 -2403
rect 11504 -2484 12694 -2467
rect 11504 -2548 11507 -2484
rect 11571 -2548 11587 -2484
rect 11651 -2548 11667 -2484
rect 11731 -2548 11747 -2484
rect 11811 -2548 11827 -2484
rect 11891 -2548 11907 -2484
rect 11971 -2548 11987 -2484
rect 12051 -2548 12067 -2484
rect 12131 -2548 12147 -2484
rect 12211 -2548 12227 -2484
rect 12291 -2548 12307 -2484
rect 12371 -2548 12387 -2484
rect 12451 -2548 12467 -2484
rect 12531 -2548 12547 -2484
rect 12611 -2548 12627 -2484
rect 12691 -2548 12694 -2484
rect 11504 -2565 12694 -2548
rect 11504 -2629 11507 -2565
rect 11571 -2629 11587 -2565
rect 11651 -2629 11667 -2565
rect 11731 -2629 11747 -2565
rect 11811 -2629 11827 -2565
rect 11891 -2629 11907 -2565
rect 11971 -2629 11987 -2565
rect 12051 -2629 12067 -2565
rect 12131 -2629 12147 -2565
rect 12211 -2629 12227 -2565
rect 12291 -2629 12307 -2565
rect 12371 -2629 12387 -2565
rect 12451 -2629 12467 -2565
rect 12531 -2629 12547 -2565
rect 12611 -2629 12627 -2565
rect 12691 -2629 12694 -2565
rect 11504 -2646 12694 -2629
rect 11504 -2710 11507 -2646
rect 11571 -2710 11587 -2646
rect 11651 -2710 11667 -2646
rect 11731 -2710 11747 -2646
rect 11811 -2710 11827 -2646
rect 11891 -2710 11907 -2646
rect 11971 -2710 11987 -2646
rect 12051 -2710 12067 -2646
rect 12131 -2710 12147 -2646
rect 12211 -2710 12227 -2646
rect 12291 -2710 12307 -2646
rect 12371 -2710 12387 -2646
rect 12451 -2710 12467 -2646
rect 12531 -2710 12547 -2646
rect 12611 -2710 12627 -2646
rect 12691 -2710 12694 -2646
rect 11504 -2727 12694 -2710
rect 11504 -2791 11507 -2727
rect 11571 -2791 11587 -2727
rect 11651 -2791 11667 -2727
rect 11731 -2791 11747 -2727
rect 11811 -2791 11827 -2727
rect 11891 -2791 11907 -2727
rect 11971 -2791 11987 -2727
rect 12051 -2791 12067 -2727
rect 12131 -2791 12147 -2727
rect 12211 -2791 12227 -2727
rect 12291 -2791 12307 -2727
rect 12371 -2791 12387 -2727
rect 12451 -2791 12467 -2727
rect 12531 -2791 12547 -2727
rect 12611 -2791 12627 -2727
rect 12691 -2791 12694 -2727
rect 11504 -2808 12694 -2791
rect 11504 -2872 11507 -2808
rect 11571 -2872 11587 -2808
rect 11651 -2872 11667 -2808
rect 11731 -2872 11747 -2808
rect 11811 -2872 11827 -2808
rect 11891 -2872 11907 -2808
rect 11971 -2872 11987 -2808
rect 12051 -2872 12067 -2808
rect 12131 -2872 12147 -2808
rect 12211 -2872 12227 -2808
rect 12291 -2872 12307 -2808
rect 12371 -2872 12387 -2808
rect 12451 -2872 12467 -2808
rect 12531 -2872 12547 -2808
rect 12611 -2872 12627 -2808
rect 12691 -2872 12694 -2808
rect 11504 -2889 12694 -2872
rect 11504 -2953 11507 -2889
rect 11571 -2953 11587 -2889
rect 11651 -2953 11667 -2889
rect 11731 -2953 11747 -2889
rect 11811 -2953 11827 -2889
rect 11891 -2953 11907 -2889
rect 11971 -2953 11987 -2889
rect 12051 -2953 12067 -2889
rect 12131 -2953 12147 -2889
rect 12211 -2953 12227 -2889
rect 12291 -2953 12307 -2889
rect 12371 -2953 12387 -2889
rect 12451 -2953 12467 -2889
rect 12531 -2953 12547 -2889
rect 12611 -2953 12627 -2889
rect 12691 -2953 12694 -2889
rect 11504 -2970 12694 -2953
rect 11504 -3034 11507 -2970
rect 11571 -3034 11587 -2970
rect 11651 -3034 11667 -2970
rect 11731 -3034 11747 -2970
rect 11811 -3034 11827 -2970
rect 11891 -3034 11907 -2970
rect 11971 -3034 11987 -2970
rect 12051 -3034 12067 -2970
rect 12131 -3034 12147 -2970
rect 12211 -3034 12227 -2970
rect 12291 -3034 12307 -2970
rect 12371 -3034 12387 -2970
rect 12451 -3034 12467 -2970
rect 12531 -3034 12547 -2970
rect 12611 -3034 12627 -2970
rect 12691 -3034 12694 -2970
rect 11504 -3051 12694 -3034
rect 11504 -3115 11507 -3051
rect 11571 -3115 11587 -3051
rect 11651 -3115 11667 -3051
rect 11731 -3115 11747 -3051
rect 11811 -3115 11827 -3051
rect 11891 -3115 11907 -3051
rect 11971 -3115 11987 -3051
rect 12051 -3115 12067 -3051
rect 12131 -3115 12147 -3051
rect 12211 -3115 12227 -3051
rect 12291 -3115 12307 -3051
rect 12371 -3115 12387 -3051
rect 12451 -3115 12467 -3051
rect 12531 -3115 12547 -3051
rect 12611 -3115 12627 -3051
rect 12691 -3115 12694 -3051
rect 11504 -3132 12694 -3115
rect 11504 -3196 11507 -3132
rect 11571 -3196 11587 -3132
rect 11651 -3196 11667 -3132
rect 11731 -3196 11747 -3132
rect 11811 -3196 11827 -3132
rect 11891 -3196 11907 -3132
rect 11971 -3196 11987 -3132
rect 12051 -3196 12067 -3132
rect 12131 -3196 12147 -3132
rect 12211 -3196 12227 -3132
rect 12291 -3196 12307 -3132
rect 12371 -3196 12387 -3132
rect 12451 -3196 12467 -3132
rect 12531 -3196 12547 -3132
rect 12611 -3196 12627 -3132
rect 12691 -3196 12694 -3132
rect 11504 -3213 12694 -3196
rect 11504 -3277 11507 -3213
rect 11571 -3277 11587 -3213
rect 11651 -3277 11667 -3213
rect 11731 -3277 11747 -3213
rect 11811 -3277 11827 -3213
rect 11891 -3277 11907 -3213
rect 11971 -3277 11987 -3213
rect 12051 -3277 12067 -3213
rect 12131 -3277 12147 -3213
rect 12211 -3277 12227 -3213
rect 12291 -3277 12307 -3213
rect 12371 -3277 12387 -3213
rect 12451 -3277 12467 -3213
rect 12531 -3277 12547 -3213
rect 12611 -3277 12627 -3213
rect 12691 -3277 12694 -3213
rect 11504 -3294 12694 -3277
rect 11504 -3358 11507 -3294
rect 11571 -3358 11587 -3294
rect 11651 -3358 11667 -3294
rect 11731 -3358 11747 -3294
rect 11811 -3358 11827 -3294
rect 11891 -3358 11907 -3294
rect 11971 -3358 11987 -3294
rect 12051 -3358 12067 -3294
rect 12131 -3358 12147 -3294
rect 12211 -3358 12227 -3294
rect 12291 -3358 12307 -3294
rect 12371 -3358 12387 -3294
rect 12451 -3358 12467 -3294
rect 12531 -3358 12547 -3294
rect 12611 -3358 12627 -3294
rect 12691 -3358 12694 -3294
rect 11504 -3375 12694 -3358
rect 11504 -3439 11507 -3375
rect 11571 -3439 11587 -3375
rect 11651 -3439 11667 -3375
rect 11731 -3439 11747 -3375
rect 11811 -3439 11827 -3375
rect 11891 -3439 11907 -3375
rect 11971 -3439 11987 -3375
rect 12051 -3439 12067 -3375
rect 12131 -3439 12147 -3375
rect 12211 -3439 12227 -3375
rect 12291 -3439 12307 -3375
rect 12371 -3439 12387 -3375
rect 12451 -3439 12467 -3375
rect 12531 -3439 12547 -3375
rect 12611 -3439 12627 -3375
rect 12691 -3439 12694 -3375
rect 11504 -3456 12694 -3439
rect 11504 -3520 11507 -3456
rect 11571 -3520 11587 -3456
rect 11651 -3520 11667 -3456
rect 11731 -3520 11747 -3456
rect 11811 -3520 11827 -3456
rect 11891 -3520 11907 -3456
rect 11971 -3520 11987 -3456
rect 12051 -3520 12067 -3456
rect 12131 -3520 12147 -3456
rect 12211 -3520 12227 -3456
rect 12291 -3520 12307 -3456
rect 12371 -3520 12387 -3456
rect 12451 -3520 12467 -3456
rect 12531 -3520 12547 -3456
rect 12611 -3520 12627 -3456
rect 12691 -3520 12694 -3456
rect 11504 -3537 12694 -3520
rect 11504 -3601 11507 -3537
rect 11571 -3601 11587 -3537
rect 11651 -3601 11667 -3537
rect 11731 -3601 11747 -3537
rect 11811 -3601 11827 -3537
rect 11891 -3601 11907 -3537
rect 11971 -3601 11987 -3537
rect 12051 -3601 12067 -3537
rect 12131 -3601 12147 -3537
rect 12211 -3601 12227 -3537
rect 12291 -3601 12307 -3537
rect 12371 -3601 12387 -3537
rect 12451 -3601 12467 -3537
rect 12531 -3601 12547 -3537
rect 12611 -3601 12627 -3537
rect 12691 -3601 12694 -3537
rect 11504 -3618 12694 -3601
rect 11504 -3682 11507 -3618
rect 11571 -3682 11587 -3618
rect 11651 -3682 11667 -3618
rect 11731 -3682 11747 -3618
rect 11811 -3682 11827 -3618
rect 11891 -3682 11907 -3618
rect 11971 -3682 11987 -3618
rect 12051 -3682 12067 -3618
rect 12131 -3682 12147 -3618
rect 12211 -3682 12227 -3618
rect 12291 -3682 12307 -3618
rect 12371 -3682 12387 -3618
rect 12451 -3682 12467 -3618
rect 12531 -3682 12547 -3618
rect 12611 -3682 12627 -3618
rect 12691 -3682 12694 -3618
rect 11504 -3699 12694 -3682
rect 11504 -3763 11507 -3699
rect 11571 -3763 11587 -3699
rect 11651 -3763 11667 -3699
rect 11731 -3763 11747 -3699
rect 11811 -3763 11827 -3699
rect 11891 -3763 11907 -3699
rect 11971 -3763 11987 -3699
rect 12051 -3763 12067 -3699
rect 12131 -3763 12147 -3699
rect 12211 -3763 12227 -3699
rect 12291 -3763 12307 -3699
rect 12371 -3763 12387 -3699
rect 12451 -3763 12467 -3699
rect 12531 -3763 12547 -3699
rect 12611 -3763 12627 -3699
rect 12691 -3763 12694 -3699
rect 11504 -3780 12694 -3763
rect 11504 -3844 11507 -3780
rect 11571 -3844 11587 -3780
rect 11651 -3844 11667 -3780
rect 11731 -3844 11747 -3780
rect 11811 -3844 11827 -3780
rect 11891 -3844 11907 -3780
rect 11971 -3844 11987 -3780
rect 12051 -3844 12067 -3780
rect 12131 -3844 12147 -3780
rect 12211 -3844 12227 -3780
rect 12291 -3844 12307 -3780
rect 12371 -3844 12387 -3780
rect 12451 -3844 12467 -3780
rect 12531 -3844 12547 -3780
rect 12611 -3844 12627 -3780
rect 12691 -3844 12694 -3780
rect 11504 -3861 12694 -3844
rect 11504 -3925 11507 -3861
rect 11571 -3925 11587 -3861
rect 11651 -3925 11667 -3861
rect 11731 -3925 11747 -3861
rect 11811 -3925 11827 -3861
rect 11891 -3925 11907 -3861
rect 11971 -3925 11987 -3861
rect 12051 -3925 12067 -3861
rect 12131 -3925 12147 -3861
rect 12211 -3925 12227 -3861
rect 12291 -3925 12307 -3861
rect 12371 -3925 12387 -3861
rect 12451 -3925 12467 -3861
rect 12531 -3925 12547 -3861
rect 12611 -3925 12627 -3861
rect 12691 -3925 12694 -3861
rect 11504 -3926 12694 -3925
use sky130_fd_io__gpio_odrvr_subv2  sky130_fd_io__gpio_odrvr_subv2_0
timestamp 1666199351
transform 1 0 0 0 1 0
box -973 -13613 15198 16619
<< labels >>
flabel locali s 310 1322 402 1368 3 FreeSans 520 0 0 0 VGND
port 1 nsew
flabel metal2 s 4692 12367 7591 13421 3 FreeSans 520 0 0 0 VGND_IO
port 2 nsew
flabel metal2 s 11116 4023 12657 5116 3 FreeSans 520 0 0 0 PAD
port 3 nsew
flabel metal2 s 11116 10856 12657 11949 3 FreeSans 520 0 0 0 PAD
port 3 nsew
flabel metal2 s 14708 -6 14748 186 3 FreeSans 520 90 0 0 PD_H[0]
port 4 nsew
flabel metal2 s 14788 -6 14828 186 3 FreeSans 520 90 0 0 PD_H[1]
port 5 nsew
flabel metal2 s 14868 -6 14908 186 3 FreeSans 520 90 0 0 PD_H[2]
port 6 nsew
flabel metal2 s 14948 -6 14988 186 3 FreeSans 520 90 0 0 PD_H[3]
port 7 nsew
flabel metal2 s 15028 -6 15068 186 3 FreeSans 520 90 0 0 TIE_LO_ESD
port 8 nsew
flabel metal2 s 13327 2545 14496 3616 3 FreeSans 520 0 0 0 VCC_IO
port 9 nsew
flabel metal1 s 13310 7954 13365 8287 3 FreeSans 520 0 0 0 PAD
port 3 nsew
flabel metal1 s 761 681 794 713 3 FreeSans 520 0 0 0 PU_H_N[0]
port 10 nsew
flabel metal1 s 6540 685 6596 718 3 FreeSans 520 0 0 0 PU_H_N[1]
port 11 nsew
flabel metal1 s 14167 280 14252 332 3 FreeSans 520 0 0 0 PU_H_N[2]
port 12 nsew
flabel metal1 s 13921 168 14073 220 3 FreeSans 520 0 0 0 PU_H_N[3]
port 13 nsew
flabel metal1 s 14164 88 14240 140 3 FreeSans 520 0 0 0 TIE_HI_ESD
port 14 nsew
flabel metal1 s 11799 737 11831 795 3 FreeSans 520 0 0 0 VCC_IO
port 9 nsew
flabel metal1 s 451 932 1620 1077 3 FreeSans 520 0 0 0 VCC_IO
port 9 nsew
flabel metal1 s 4107 173 5276 318 3 FreeSans 520 0 0 0 VCC_IO
port 9 nsew
flabel metal1 s 2496 8314 2549 8360 3 FreeSans 520 0 0 0 VGND_IO
port 2 nsew
flabel metal1 s 49 -1067 83 -1013 3 FreeSans 520 270 0 0 FORCE_HI_H_N
port 15 nsew
flabel metal1 s 377 -1075 415 -1020 3 FreeSans 520 270 0 0 FORCE_LO_H
port 16 nsew
flabel metal1 s 258 -1075 313 -1023 3 FreeSans 520 270 0 0 FORCE_LOVOL_H
port 17 nsew
flabel metal1 s 168 -1074 206 -1007 3 FreeSans 520 270 0 0 VSSIO_AMX
port 18 nsew
<< properties >>
string GDS_END 48517894
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 48364862
<< end >>
