magic
tech sky130B
magscale 1 2
timestamp 1669056001
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 348786 700340 348792 700392
rect 348844 700380 348850 700392
rect 364334 700380 364340 700392
rect 348844 700352 364340 700380
rect 348844 700340 348850 700352
rect 364334 700340 364340 700352
rect 364392 700340 364398 700392
rect 8110 700272 8116 700324
rect 8168 700312 8174 700324
rect 250438 700312 250444 700324
rect 8168 700284 250444 700312
rect 8168 700272 8174 700284
rect 250438 700272 250444 700284
rect 250496 700272 250502 700324
rect 332502 700272 332508 700324
rect 332560 700312 332566 700324
rect 364426 700312 364432 700324
rect 332560 700284 364432 700312
rect 332560 700272 332566 700284
rect 364426 700272 364432 700284
rect 364484 700272 364490 700324
rect 218974 699660 218980 699712
rect 219032 699700 219038 699712
rect 220078 699700 220084 699712
rect 219032 699672 220084 699700
rect 219032 699660 219038 699672
rect 220078 699660 220084 699672
rect 220136 699660 220142 699712
rect 396718 699660 396724 699712
rect 396776 699700 396782 699712
rect 397454 699700 397460 699712
rect 396776 699672 397460 699700
rect 396776 699660 396782 699672
rect 397454 699660 397460 699672
rect 397512 699660 397518 699712
rect 363598 698640 363604 698692
rect 363656 698680 363662 698692
rect 364978 698680 364984 698692
rect 363656 698652 364984 698680
rect 363656 698640 363662 698652
rect 364978 698640 364984 698652
rect 365036 698640 365042 698692
rect 266354 697552 266360 697604
rect 266412 697592 266418 697604
rect 267642 697592 267648 697604
rect 266412 697564 267648 697592
rect 266412 697552 266418 697564
rect 267642 697552 267648 697564
rect 267700 697552 267706 697604
rect 378778 696940 378784 696992
rect 378836 696980 378842 696992
rect 580166 696980 580172 696992
rect 378836 696952 580172 696980
rect 378836 696940 378842 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 369854 683176 369860 683188
rect 3476 683148 369860 683176
rect 3476 683136 3482 683148
rect 369854 683136 369860 683148
rect 369912 683136 369918 683188
rect 3418 671032 3424 671084
rect 3476 671072 3482 671084
rect 7558 671072 7564 671084
rect 3476 671044 7564 671072
rect 3476 671032 3482 671044
rect 7558 671032 7564 671044
rect 7616 671032 7622 671084
rect 359458 670692 359464 670744
rect 359516 670732 359522 670744
rect 580166 670732 580172 670744
rect 359516 670704 580172 670732
rect 359516 670692 359522 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 2774 656956 2780 657008
rect 2832 656996 2838 657008
rect 4798 656996 4804 657008
rect 2832 656968 4804 656996
rect 2832 656956 2838 656968
rect 4798 656956 4804 656968
rect 4856 656956 4862 657008
rect 359550 643084 359556 643136
rect 359608 643124 359614 643136
rect 580166 643124 580172 643136
rect 359608 643096 580172 643124
rect 359608 643084 359614 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 371418 632108 371424 632120
rect 3476 632080 371424 632108
rect 3476 632068 3482 632080
rect 371418 632068 371424 632080
rect 371476 632068 371482 632120
rect 359642 630640 359648 630692
rect 359700 630680 359706 630692
rect 579982 630680 579988 630692
rect 359700 630652 579988 630680
rect 359700 630640 359706 630652
rect 579982 630640 579988 630652
rect 580040 630640 580046 630692
rect 382918 616836 382924 616888
rect 382976 616876 382982 616888
rect 580166 616876 580172 616888
rect 382976 616848 580172 616876
rect 382976 616836 382982 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3510 605820 3516 605872
rect 3568 605860 3574 605872
rect 142798 605860 142804 605872
rect 3568 605832 142804 605860
rect 3568 605820 3574 605832
rect 142798 605820 142804 605832
rect 142856 605820 142862 605872
rect 367738 590656 367744 590708
rect 367796 590696 367802 590708
rect 580166 590696 580172 590708
rect 367796 590668 580172 590696
rect 367796 590656 367802 590668
rect 580166 590656 580172 590668
rect 580224 590656 580230 590708
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 372614 579680 372620 579692
rect 3384 579652 372620 579680
rect 3384 579640 3390 579652
rect 372614 579640 372620 579652
rect 372672 579640 372678 579692
rect 358446 576852 358452 576904
rect 358504 576892 358510 576904
rect 580166 576892 580172 576904
rect 358504 576864 580172 576892
rect 358504 576852 358510 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 3234 565836 3240 565888
rect 3292 565876 3298 565888
rect 195238 565876 195244 565888
rect 3292 565848 195244 565876
rect 3292 565836 3298 565848
rect 195238 565836 195244 565848
rect 195296 565836 195302 565888
rect 376018 563048 376024 563100
rect 376076 563088 376082 563100
rect 580166 563088 580172 563100
rect 376076 563060 580172 563088
rect 376076 563048 376082 563060
rect 580166 563048 580172 563060
rect 580224 563048 580230 563100
rect 3326 553392 3332 553444
rect 3384 553432 3390 553444
rect 10318 553432 10324 553444
rect 3384 553404 10324 553432
rect 3384 553392 3390 553404
rect 10318 553392 10324 553404
rect 10376 553392 10382 553444
rect 377398 536800 377404 536852
rect 377456 536840 377462 536852
rect 579890 536840 579896 536852
rect 377456 536812 579896 536840
rect 377456 536800 377462 536812
rect 579890 536800 579896 536812
rect 579948 536800 579954 536852
rect 2958 527144 2964 527196
rect 3016 527184 3022 527196
rect 373994 527184 374000 527196
rect 3016 527156 374000 527184
rect 3016 527144 3022 527156
rect 373994 527144 374000 527156
rect 374052 527144 374058 527196
rect 392578 524424 392584 524476
rect 392636 524464 392642 524476
rect 580166 524464 580172 524476
rect 392636 524436 580172 524464
rect 392636 524424 392642 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3510 514768 3516 514820
rect 3568 514808 3574 514820
rect 13078 514808 13084 514820
rect 3568 514780 13084 514808
rect 3568 514768 3574 514780
rect 13078 514768 13084 514780
rect 13136 514768 13142 514820
rect 360838 511232 360844 511284
rect 360896 511272 360902 511284
rect 580258 511272 580264 511284
rect 360896 511244 580264 511272
rect 360896 511232 360902 511244
rect 580258 511232 580264 511244
rect 580316 511232 580322 511284
rect 3050 500964 3056 501016
rect 3108 501004 3114 501016
rect 298738 501004 298744 501016
rect 3108 500976 298744 501004
rect 3108 500964 3114 500976
rect 298738 500964 298744 500976
rect 298796 500964 298802 501016
rect 355318 484372 355324 484424
rect 355376 484412 355382 484424
rect 580166 484412 580172 484424
rect 355376 484384 580172 484412
rect 355376 484372 355382 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 3050 474716 3056 474768
rect 3108 474756 3114 474768
rect 374086 474756 374092 474768
rect 3108 474728 374092 474756
rect 3108 474716 3114 474728
rect 374086 474716 374092 474728
rect 374144 474716 374150 474768
rect 363690 473968 363696 474020
rect 363748 474008 363754 474020
rect 412634 474008 412640 474020
rect 363748 473980 412640 474008
rect 363748 473968 363754 473980
rect 412634 473968 412640 473980
rect 412692 473968 412698 474020
rect 356698 472608 356704 472660
rect 356756 472648 356762 472660
rect 392578 472648 392584 472660
rect 356756 472620 392584 472648
rect 356756 472608 356762 472620
rect 392578 472608 392584 472620
rect 392636 472608 392642 472660
rect 367830 470568 367836 470620
rect 367888 470608 367894 470620
rect 580074 470608 580080 470620
rect 367888 470580 580080 470608
rect 367888 470568 367894 470580
rect 580074 470568 580080 470580
rect 580132 470568 580138 470620
rect 360930 469820 360936 469872
rect 360988 469860 360994 469872
rect 527174 469860 527180 469872
rect 360988 469832 527180 469860
rect 360988 469820 360994 469832
rect 527174 469820 527180 469832
rect 527232 469820 527238 469872
rect 358078 468460 358084 468512
rect 358136 468500 358142 468512
rect 367738 468500 367744 468512
rect 358136 468472 367744 468500
rect 358136 468460 358142 468472
rect 367738 468460 367744 468472
rect 367796 468460 367802 468512
rect 40034 467100 40040 467152
rect 40092 467140 40098 467152
rect 368566 467140 368572 467152
rect 40092 467112 368572 467140
rect 40092 467100 40098 467112
rect 368566 467100 368572 467112
rect 368624 467100 368630 467152
rect 104894 465672 104900 465724
rect 104952 465712 104958 465724
rect 276014 465712 276020 465724
rect 104952 465684 276020 465712
rect 104952 465672 104958 465684
rect 276014 465672 276020 465684
rect 276072 465672 276078 465724
rect 362310 465672 362316 465724
rect 362368 465712 362374 465724
rect 477494 465712 477500 465724
rect 362368 465684 477500 465712
rect 362368 465672 362374 465684
rect 477494 465672 477500 465684
rect 477552 465672 477558 465724
rect 276014 465060 276020 465112
rect 276072 465100 276078 465112
rect 277302 465100 277308 465112
rect 276072 465072 277308 465100
rect 276072 465060 276078 465072
rect 277302 465060 277308 465072
rect 277360 465100 277366 465112
rect 368658 465100 368664 465112
rect 277360 465072 368664 465100
rect 277360 465060 277366 465072
rect 368658 465060 368664 465072
rect 368716 465060 368722 465112
rect 169754 464312 169760 464364
rect 169812 464352 169818 464364
rect 273254 464352 273260 464364
rect 169812 464324 273260 464352
rect 169812 464312 169818 464324
rect 273254 464312 273260 464324
rect 273312 464312 273318 464364
rect 362218 464312 362224 464364
rect 362276 464352 362282 464364
rect 542354 464352 542360 464364
rect 362276 464324 542360 464352
rect 362276 464312 362282 464324
rect 542354 464312 542360 464324
rect 542412 464312 542418 464364
rect 273254 463700 273260 463752
rect 273312 463740 273318 463752
rect 274542 463740 274548 463752
rect 273312 463712 274548 463740
rect 273312 463700 273318 463712
rect 274542 463700 274548 463712
rect 274600 463740 274606 463752
rect 367094 463740 367100 463752
rect 274600 463712 367100 463740
rect 274600 463700 274606 463712
rect 367094 463700 367100 463712
rect 367152 463700 367158 463752
rect 356238 462952 356244 463004
rect 356296 462992 356302 463004
rect 377398 462992 377404 463004
rect 356296 462964 377404 462992
rect 356296 462952 356302 462964
rect 377398 462952 377404 462964
rect 377456 462952 377462 463004
rect 3510 462544 3516 462596
rect 3568 462584 3574 462596
rect 8938 462584 8944 462596
rect 3568 462556 8944 462584
rect 3568 462544 3574 462556
rect 8938 462544 8944 462556
rect 8996 462544 9002 462596
rect 234614 461592 234620 461644
rect 234672 461632 234678 461644
rect 275278 461632 275284 461644
rect 234672 461604 275284 461632
rect 234672 461592 234678 461604
rect 275278 461592 275284 461604
rect 275336 461592 275342 461644
rect 363046 461592 363052 461644
rect 363104 461632 363110 461644
rect 396718 461632 396724 461644
rect 363104 461604 396724 461632
rect 363104 461592 363110 461604
rect 396718 461592 396724 461604
rect 396776 461592 396782 461644
rect 275278 460912 275284 460964
rect 275336 460952 275342 460964
rect 365806 460952 365812 460964
rect 275336 460924 365812 460952
rect 275336 460912 275342 460924
rect 365806 460912 365812 460924
rect 365864 460912 365870 460964
rect 357250 460232 357256 460284
rect 357308 460272 357314 460284
rect 367830 460272 367836 460284
rect 357308 460244 367836 460272
rect 357308 460232 357314 460244
rect 367830 460232 367836 460244
rect 367888 460232 367894 460284
rect 363230 460164 363236 460216
rect 363288 460204 363294 460216
rect 429194 460204 429200 460216
rect 363288 460176 429200 460204
rect 363288 460164 363294 460176
rect 429194 460164 429200 460176
rect 429252 460164 429258 460216
rect 360654 458804 360660 458856
rect 360712 458844 360718 458856
rect 558914 458844 558920 458856
rect 360712 458816 558920 458844
rect 360712 458804 360718 458816
rect 558914 458804 558920 458816
rect 558972 458804 558978 458856
rect 334710 457104 334716 457156
rect 334768 457144 334774 457156
rect 373534 457144 373540 457156
rect 334768 457116 373540 457144
rect 334768 457104 334774 457116
rect 373534 457104 373540 457116
rect 373592 457104 373598 457156
rect 334894 457036 334900 457088
rect 334952 457076 334958 457088
rect 375742 457076 375748 457088
rect 334952 457048 375748 457076
rect 334952 457036 334958 457048
rect 375742 457036 375748 457048
rect 375800 457036 375806 457088
rect 333514 456968 333520 457020
rect 333572 457008 333578 457020
rect 380158 457008 380164 457020
rect 333572 456980 380164 457008
rect 333572 456968 333578 456980
rect 380158 456968 380164 456980
rect 380216 456968 380222 457020
rect 332042 456900 332048 456952
rect 332100 456940 332106 456952
rect 378226 456940 378232 456952
rect 332100 456912 378232 456940
rect 332100 456900 332106 456912
rect 378226 456900 378232 456912
rect 378284 456900 378290 456952
rect 320818 456832 320824 456884
rect 320876 456872 320882 456884
rect 381262 456872 381268 456884
rect 320876 456844 381268 456872
rect 320876 456832 320882 456844
rect 381262 456832 381268 456844
rect 381320 456832 381326 456884
rect 355962 456764 355968 456816
rect 356020 456804 356026 456816
rect 580166 456804 580172 456816
rect 356020 456776 580172 456804
rect 356020 456764 356026 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 358630 456084 358636 456136
rect 358688 456124 358694 456136
rect 382918 456124 382924 456136
rect 358688 456096 382924 456124
rect 358688 456084 358694 456096
rect 382918 456084 382924 456096
rect 382976 456084 382982 456136
rect 362310 456016 362316 456068
rect 362368 456056 362374 456068
rect 462314 456056 462320 456068
rect 362368 456028 462320 456056
rect 362368 456016 362374 456028
rect 462314 456016 462320 456028
rect 462372 456016 462378 456068
rect 359182 455880 359188 455932
rect 359240 455920 359246 455932
rect 359642 455920 359648 455932
rect 359240 455892 359648 455920
rect 359240 455880 359246 455892
rect 359642 455880 359648 455892
rect 359700 455880 359706 455932
rect 363506 455880 363512 455932
rect 363564 455920 363570 455932
rect 363690 455920 363696 455932
rect 363564 455892 363696 455920
rect 363564 455880 363570 455892
rect 363690 455880 363696 455892
rect 363748 455880 363754 455932
rect 336458 455812 336464 455864
rect 336516 455852 336522 455864
rect 364426 455852 364432 455864
rect 336516 455824 364432 455852
rect 336516 455812 336522 455824
rect 364426 455812 364432 455824
rect 364484 455812 364490 455864
rect 327810 455744 327816 455796
rect 327868 455784 327874 455796
rect 360470 455784 360476 455796
rect 327868 455756 360476 455784
rect 327868 455744 327874 455756
rect 360470 455744 360476 455756
rect 360528 455744 360534 455796
rect 324958 455676 324964 455728
rect 325016 455716 325022 455728
rect 362494 455716 362500 455728
rect 325016 455688 362500 455716
rect 325016 455676 325022 455688
rect 362494 455676 362500 455688
rect 362552 455676 362558 455728
rect 322198 455608 322204 455660
rect 322256 455648 322262 455660
rect 363506 455648 363512 455660
rect 322256 455620 363512 455648
rect 322256 455608 322262 455620
rect 363506 455608 363512 455620
rect 363564 455608 363570 455660
rect 301498 455540 301504 455592
rect 301556 455580 301562 455592
rect 356698 455580 356704 455592
rect 301556 455552 356704 455580
rect 301556 455540 301562 455552
rect 356698 455540 356704 455552
rect 356756 455580 356762 455592
rect 356974 455580 356980 455592
rect 356756 455552 356980 455580
rect 356756 455540 356762 455552
rect 356974 455540 356980 455552
rect 357032 455540 357038 455592
rect 304258 455472 304264 455524
rect 304316 455512 304322 455524
rect 364334 455512 364340 455524
rect 304316 455484 364340 455512
rect 304316 455472 304322 455484
rect 364334 455472 364340 455484
rect 364392 455512 364398 455524
rect 364702 455512 364708 455524
rect 364392 455484 364708 455512
rect 364392 455472 364398 455484
rect 364702 455472 364708 455484
rect 364760 455472 364766 455524
rect 298830 455404 298836 455456
rect 298888 455444 298894 455456
rect 359182 455444 359188 455456
rect 298888 455416 359188 455444
rect 298888 455404 298894 455416
rect 359182 455404 359188 455416
rect 359240 455404 359246 455456
rect 278590 454928 278596 454980
rect 278648 454968 278654 454980
rect 350718 454968 350724 454980
rect 278648 454940 350724 454968
rect 278648 454928 278654 454940
rect 350718 454928 350724 454940
rect 350776 454928 350782 454980
rect 307018 454860 307024 454912
rect 307076 454900 307082 454912
rect 367186 454900 367192 454912
rect 307076 454872 367192 454900
rect 307076 454860 307082 454872
rect 367186 454860 367192 454872
rect 367244 454860 367250 454912
rect 278682 454792 278688 454844
rect 278740 454832 278746 454844
rect 352098 454832 352104 454844
rect 278740 454804 352104 454832
rect 278740 454792 278746 454804
rect 352098 454792 352104 454804
rect 352156 454792 352162 454844
rect 358722 454792 358728 454844
rect 358780 454832 358786 454844
rect 376018 454832 376024 454844
rect 358780 454804 376024 454832
rect 358780 454792 358786 454804
rect 376018 454792 376024 454804
rect 376076 454792 376082 454844
rect 337930 454724 337936 454776
rect 337988 454764 337994 454776
rect 363230 454764 363236 454776
rect 337988 454736 363236 454764
rect 337988 454724 337994 454736
rect 363230 454724 363236 454736
rect 363288 454724 363294 454776
rect 338022 454656 338028 454708
rect 338080 454696 338086 454708
rect 360654 454696 360660 454708
rect 338080 454668 360660 454696
rect 338080 454656 338086 454668
rect 360654 454656 360660 454668
rect 360712 454656 360718 454708
rect 361574 454656 361580 454708
rect 361632 454696 361638 454708
rect 494054 454696 494060 454708
rect 361632 454668 494060 454696
rect 361632 454656 361638 454668
rect 494054 454656 494060 454668
rect 494112 454656 494118 454708
rect 334618 454588 334624 454640
rect 334676 454628 334682 454640
rect 363322 454628 363328 454640
rect 334676 454600 363328 454628
rect 334676 454588 334682 454600
rect 363322 454588 363328 454600
rect 363380 454588 363386 454640
rect 289814 454520 289820 454572
rect 289872 454560 289878 454572
rect 349982 454560 349988 454572
rect 289872 454532 349988 454560
rect 289872 454520 289878 454532
rect 349982 454520 349988 454532
rect 350040 454520 350046 454572
rect 317598 454452 317604 454504
rect 317656 454492 317662 454504
rect 377582 454492 377588 454504
rect 317656 454464 377588 454492
rect 317656 454452 317662 454464
rect 377582 454452 377588 454464
rect 377640 454452 377646 454504
rect 322382 454384 322388 454436
rect 322440 454424 322446 454436
rect 382458 454424 382464 454436
rect 322440 454396 382464 454424
rect 322440 454384 322446 454396
rect 382458 454384 382464 454396
rect 382516 454384 382522 454436
rect 316862 454316 316868 454368
rect 316920 454356 316926 454368
rect 376938 454356 376944 454368
rect 316920 454328 376944 454356
rect 316920 454316 316926 454328
rect 376938 454316 376944 454328
rect 376996 454316 377002 454368
rect 319438 454248 319444 454300
rect 319496 454288 319502 454300
rect 379790 454288 379796 454300
rect 319496 454260 379796 454288
rect 319496 454248 319502 454260
rect 379790 454248 379796 454260
rect 379848 454248 379854 454300
rect 340782 454180 340788 454232
rect 340840 454220 340846 454232
rect 357618 454220 357624 454232
rect 340840 454192 357624 454220
rect 340840 454180 340846 454192
rect 357618 454180 357624 454192
rect 357676 454220 357682 454232
rect 358722 454220 358728 454232
rect 357676 454192 358728 454220
rect 357676 454180 357682 454192
rect 358722 454180 358728 454192
rect 358780 454180 358786 454232
rect 341518 454112 341524 454164
rect 341576 454152 341582 454164
rect 360930 454152 360936 454164
rect 341576 454124 360936 454152
rect 341576 454112 341582 454124
rect 360930 454112 360936 454124
rect 360988 454112 360994 454164
rect 340506 454044 340512 454096
rect 340564 454084 340570 454096
rect 361574 454084 361580 454096
rect 340564 454056 361580 454084
rect 340564 454044 340570 454056
rect 361574 454044 361580 454056
rect 361632 454044 361638 454096
rect 359090 453976 359096 454028
rect 359148 454016 359154 454028
rect 359550 454016 359556 454028
rect 359148 453988 359556 454016
rect 359148 453976 359154 453988
rect 359550 453976 359556 453988
rect 359608 453976 359614 454028
rect 337838 453568 337844 453620
rect 337896 453608 337902 453620
rect 358078 453608 358084 453620
rect 337896 453580 358084 453608
rect 337896 453568 337902 453580
rect 358078 453568 358084 453580
rect 358136 453568 358142 453620
rect 294598 453500 294604 453552
rect 294656 453540 294662 453552
rect 355410 453540 355416 453552
rect 294656 453512 355416 453540
rect 294656 453500 294662 453512
rect 355410 453500 355416 453512
rect 355468 453540 355474 453552
rect 355962 453540 355968 453552
rect 355468 453512 355968 453540
rect 355468 453500 355474 453512
rect 355962 453500 355968 453512
rect 356020 453500 356026 453552
rect 335078 453432 335084 453484
rect 335136 453472 335142 453484
rect 359090 453472 359096 453484
rect 335136 453444 359096 453472
rect 335136 453432 335142 453444
rect 359090 453432 359096 453444
rect 359148 453432 359154 453484
rect 360378 453432 360384 453484
rect 360436 453472 360442 453484
rect 378778 453472 378784 453484
rect 360436 453444 378784 453472
rect 360436 453432 360442 453444
rect 378778 453432 378784 453444
rect 378836 453432 378842 453484
rect 299474 453364 299480 453416
rect 299532 453404 299538 453416
rect 309042 453404 309048 453416
rect 299532 453376 309048 453404
rect 299532 453364 299538 453376
rect 309042 453364 309048 453376
rect 309100 453364 309106 453416
rect 357342 453296 357348 453348
rect 357400 453336 357406 453348
rect 580350 453336 580356 453348
rect 357400 453308 580356 453336
rect 357400 453296 357406 453308
rect 580350 453296 580356 453308
rect 580408 453296 580414 453348
rect 327902 453228 327908 453280
rect 327960 453268 327966 453280
rect 356054 453268 356060 453280
rect 327960 453240 356060 453268
rect 327960 453228 327966 453240
rect 356054 453228 356060 453240
rect 356112 453268 356118 453280
rect 357250 453268 357256 453280
rect 356112 453240 357256 453268
rect 356112 453228 356118 453240
rect 357250 453228 357256 453240
rect 357308 453228 357314 453280
rect 325050 453160 325056 453212
rect 325108 453200 325114 453212
rect 371234 453200 371240 453212
rect 325108 453172 371240 453200
rect 325108 453160 325114 453172
rect 371234 453160 371240 453172
rect 371292 453160 371298 453212
rect 315298 453092 315304 453144
rect 315356 453132 315362 453144
rect 369946 453132 369952 453144
rect 315356 453104 369952 453132
rect 315356 453092 315362 453104
rect 369946 453092 369952 453104
rect 370004 453092 370010 453144
rect 323670 453024 323676 453076
rect 323728 453064 323734 453076
rect 382734 453064 382740 453076
rect 323728 453036 382740 453064
rect 323728 453024 323734 453036
rect 382734 453024 382740 453036
rect 382792 453024 382798 453076
rect 322290 452956 322296 453008
rect 322348 452996 322354 453008
rect 381630 452996 381636 453008
rect 322348 452968 381636 452996
rect 322348 452956 322354 452968
rect 381630 452956 381636 452968
rect 381688 452956 381694 453008
rect 316770 452888 316776 452940
rect 316828 452928 316834 452940
rect 376110 452928 376116 452940
rect 316828 452900 376116 452928
rect 316828 452888 316834 452900
rect 376110 452888 376116 452900
rect 376168 452888 376174 452940
rect 318058 452820 318064 452872
rect 318116 452860 318122 452872
rect 377214 452860 377220 452872
rect 318116 452832 377220 452860
rect 318116 452820 318122 452832
rect 377214 452820 377220 452832
rect 377272 452820 377278 452872
rect 323578 452752 323584 452804
rect 323636 452792 323642 452804
rect 383838 452792 383844 452804
rect 323636 452764 383844 452792
rect 323636 452752 323642 452764
rect 383838 452752 383844 452764
rect 383896 452752 383902 452804
rect 316678 452684 316684 452736
rect 316736 452724 316742 452736
rect 376754 452724 376760 452736
rect 316736 452696 376760 452724
rect 316736 452684 316742 452696
rect 376754 452684 376760 452696
rect 376812 452684 376818 452736
rect 340690 452616 340696 452668
rect 340748 452656 340754 452668
rect 356330 452656 356336 452668
rect 340748 452628 356336 452656
rect 340748 452616 340754 452628
rect 356330 452616 356336 452628
rect 356388 452656 356394 452668
rect 357342 452656 357348 452668
rect 356388 452628 357348 452656
rect 356388 452616 356394 452628
rect 357342 452616 357348 452628
rect 357400 452616 357406 452668
rect 281258 452140 281264 452192
rect 281316 452180 281322 452192
rect 347406 452180 347412 452192
rect 281316 452152 347412 452180
rect 281316 452140 281322 452152
rect 347406 452140 347412 452152
rect 347464 452140 347470 452192
rect 294690 452072 294696 452124
rect 294748 452112 294754 452124
rect 353662 452112 353668 452124
rect 294748 452084 353668 452112
rect 294748 452072 294754 452084
rect 353662 452072 353668 452084
rect 353720 452072 353726 452124
rect 340138 452004 340144 452056
rect 340196 452044 340202 452056
rect 384574 452044 384580 452056
rect 340196 452016 384580 452044
rect 340196 452004 340202 452016
rect 384574 452004 384580 452016
rect 384632 452004 384638 452056
rect 279878 451936 279884 451988
rect 279936 451976 279942 451988
rect 354858 451976 354864 451988
rect 279936 451948 354864 451976
rect 279936 451936 279942 451948
rect 354858 451936 354864 451948
rect 354916 451936 354922 451988
rect 291838 451868 291844 451920
rect 291896 451908 291902 451920
rect 350534 451908 350540 451920
rect 291896 451880 350540 451908
rect 291896 451868 291902 451880
rect 350534 451868 350540 451880
rect 350592 451868 350598 451920
rect 371234 451868 371240 451920
rect 371292 451908 371298 451920
rect 385034 451908 385040 451920
rect 371292 451880 385040 451908
rect 371292 451868 371298 451880
rect 385034 451868 385040 451880
rect 385092 451868 385098 451920
rect 341794 451800 341800 451852
rect 341852 451840 341858 451852
rect 379054 451840 379060 451852
rect 341852 451812 379060 451840
rect 341852 451800 341858 451812
rect 379054 451800 379060 451812
rect 379112 451800 379118 451852
rect 337378 451732 337384 451784
rect 337436 451772 337442 451784
rect 351454 451772 351460 451784
rect 337436 451744 351460 451772
rect 337436 451732 337442 451744
rect 351454 451732 351460 451744
rect 351512 451732 351518 451784
rect 338758 451664 338764 451716
rect 338816 451704 338822 451716
rect 352558 451704 352564 451716
rect 338816 451676 352564 451704
rect 338816 451664 338822 451676
rect 352558 451664 352564 451676
rect 352616 451664 352622 451716
rect 334802 451596 334808 451648
rect 334860 451636 334866 451648
rect 370222 451636 370228 451648
rect 334860 451608 370228 451636
rect 334860 451596 334866 451608
rect 370222 451596 370228 451608
rect 370280 451596 370286 451648
rect 340966 451528 340972 451580
rect 341024 451568 341030 451580
rect 382550 451568 382556 451580
rect 341024 451540 382556 451568
rect 341024 451528 341030 451540
rect 382550 451528 382556 451540
rect 382608 451528 382614 451580
rect 341610 451460 341616 451512
rect 341668 451500 341674 451512
rect 341668 451472 350534 451500
rect 341668 451460 341674 451472
rect 342254 451392 342260 451444
rect 342312 451432 342318 451444
rect 350506 451432 350534 451472
rect 365806 451432 365812 451444
rect 342312 451404 348280 451432
rect 350506 451404 365812 451432
rect 342312 451392 342318 451404
rect 348142 451364 348148 451376
rect 340846 451336 348148 451364
rect 340322 451256 340328 451308
rect 340380 451296 340386 451308
rect 340846 451296 340874 451336
rect 348142 451324 348148 451336
rect 348200 451324 348206 451376
rect 348252 451364 348280 451404
rect 365806 451392 365812 451404
rect 365864 451392 365870 451444
rect 352190 451364 352196 451376
rect 348252 451336 352196 451364
rect 352190 451324 352196 451336
rect 352248 451324 352254 451376
rect 362218 451324 362224 451376
rect 362276 451364 362282 451376
rect 369118 451364 369124 451376
rect 362276 451336 369124 451364
rect 362276 451324 362282 451336
rect 369118 451324 369124 451336
rect 369176 451324 369182 451376
rect 340380 451268 340874 451296
rect 340380 451256 340386 451268
rect 341886 451256 341892 451308
rect 341944 451296 341950 451308
rect 349246 451296 349252 451308
rect 341944 451268 349252 451296
rect 341944 451256 341950 451268
rect 349246 451256 349252 451268
rect 349304 451256 349310 451308
rect 358538 451256 358544 451308
rect 358596 451296 358602 451308
rect 363966 451296 363972 451308
rect 358596 451268 363972 451296
rect 358596 451256 358602 451268
rect 363966 451256 363972 451268
rect 364024 451256 364030 451308
rect 369946 451256 369952 451308
rect 370004 451296 370010 451308
rect 375374 451296 375380 451308
rect 370004 451268 375380 451296
rect 370004 451256 370010 451268
rect 375374 451256 375380 451268
rect 375432 451256 375438 451308
rect 297358 450848 297364 450900
rect 297416 450888 297422 450900
rect 356238 450888 356244 450900
rect 297416 450860 356244 450888
rect 297416 450848 297422 450860
rect 356238 450848 356244 450860
rect 356296 450848 356302 450900
rect 266354 450780 266360 450832
rect 266412 450820 266418 450832
rect 271322 450820 271328 450832
rect 266412 450792 271328 450820
rect 266412 450780 266418 450792
rect 271322 450780 271328 450792
rect 271380 450820 271386 450832
rect 365714 450820 365720 450832
rect 271380 450792 365720 450820
rect 271380 450780 271386 450792
rect 365714 450780 365720 450792
rect 365772 450780 365778 450832
rect 302878 450712 302884 450764
rect 302936 450752 302942 450764
rect 362310 450752 362316 450764
rect 302936 450724 362316 450752
rect 302936 450712 302942 450724
rect 362310 450712 362316 450724
rect 362368 450712 362374 450764
rect 294782 450644 294788 450696
rect 294840 450684 294846 450696
rect 353294 450684 353300 450696
rect 294840 450656 353300 450684
rect 294840 450644 294846 450656
rect 353294 450644 353300 450656
rect 353352 450644 353358 450696
rect 355226 450644 355232 450696
rect 355284 450684 355290 450696
rect 356698 450684 356704 450696
rect 355284 450656 356704 450684
rect 355284 450644 355290 450656
rect 356698 450644 356704 450656
rect 356756 450644 356762 450696
rect 320910 450576 320916 450628
rect 320968 450616 320974 450628
rect 380526 450616 380532 450628
rect 320968 450588 380532 450616
rect 320968 450576 320974 450588
rect 380526 450576 380532 450588
rect 380584 450576 380590 450628
rect 136634 450508 136640 450560
rect 136692 450548 136698 450560
rect 136692 450520 296714 450548
rect 136692 450508 136698 450520
rect 296686 450480 296714 450520
rect 356238 450508 356244 450560
rect 356296 450548 356302 450560
rect 356606 450548 356612 450560
rect 356296 450520 356612 450548
rect 356296 450508 356302 450520
rect 356606 450508 356612 450520
rect 356664 450508 356670 450560
rect 356698 450508 356704 450560
rect 356756 450548 356762 450560
rect 580258 450548 580264 450560
rect 356756 450520 580264 450548
rect 356756 450508 356762 450520
rect 580258 450508 580264 450520
rect 580316 450508 580322 450560
rect 307754 450480 307760 450492
rect 296686 450452 307760 450480
rect 307754 450440 307760 450452
rect 307812 450480 307818 450492
rect 367646 450480 367652 450492
rect 307812 450452 367652 450480
rect 307812 450440 307818 450452
rect 367646 450440 367652 450452
rect 367704 450440 367710 450492
rect 295978 450372 295984 450424
rect 296036 450412 296042 450424
rect 355318 450412 355324 450424
rect 296036 450384 355324 450412
rect 296036 450372 296042 450384
rect 355318 450372 355324 450384
rect 355376 450412 355382 450424
rect 355502 450412 355508 450424
rect 355376 450384 355508 450412
rect 355376 450372 355382 450384
rect 355502 450372 355508 450384
rect 355560 450372 355566 450424
rect 321002 450304 321008 450356
rect 321060 450344 321066 450356
rect 380894 450344 380900 450356
rect 321060 450316 380900 450344
rect 321060 450304 321066 450316
rect 380894 450304 380900 450316
rect 380952 450304 380958 450356
rect 318150 450236 318156 450288
rect 318208 450276 318214 450288
rect 378318 450276 378324 450288
rect 318208 450248 378324 450276
rect 318208 450236 318214 450248
rect 378318 450236 378324 450248
rect 378376 450236 378382 450288
rect 319530 450168 319536 450220
rect 319588 450208 319594 450220
rect 379652 450208 379658 450220
rect 319588 450180 379658 450208
rect 319588 450168 319594 450180
rect 379652 450168 379658 450180
rect 379710 450168 379716 450220
rect 313918 450100 313924 450152
rect 313976 450140 313982 450152
rect 374500 450140 374506 450152
rect 313976 450112 374506 450140
rect 313976 450100 313982 450112
rect 374500 450100 374506 450112
rect 374558 450100 374564 450152
rect 339310 450032 339316 450084
rect 339368 450072 339374 450084
rect 366542 450072 366548 450084
rect 339368 450044 366548 450072
rect 339368 450032 339374 450044
rect 366542 450032 366548 450044
rect 366600 450032 366606 450084
rect 342162 449964 342168 450016
rect 342220 450004 342226 450016
rect 351086 450004 351092 450016
rect 342220 449976 351092 450004
rect 342220 449964 342226 449976
rect 351086 449964 351092 449976
rect 351144 449964 351150 450016
rect 353294 449964 353300 450016
rect 353352 450004 353358 450016
rect 354122 450004 354128 450016
rect 353352 449976 354128 450004
rect 353352 449964 353358 449976
rect 354122 449964 354128 449976
rect 354180 450004 354186 450016
rect 388438 450004 388444 450016
rect 354180 449976 388444 450004
rect 354180 449964 354186 449976
rect 388438 449964 388444 449976
rect 388496 449964 388502 450016
rect 332226 449896 332232 449948
rect 332284 449936 332290 449948
rect 354766 449936 354772 449948
rect 332284 449908 354772 449936
rect 332284 449896 332290 449908
rect 354766 449896 354772 449908
rect 354824 449936 354830 449948
rect 389818 449936 389824 449948
rect 354824 449908 389824 449936
rect 354824 449896 354830 449908
rect 389818 449896 389824 449908
rect 389876 449896 389882 449948
rect 342346 449488 342352 449540
rect 342404 449528 342410 449540
rect 349614 449528 349620 449540
rect 342404 449500 349620 449528
rect 342404 449488 342410 449500
rect 349614 449488 349620 449500
rect 349672 449488 349678 449540
rect 358538 449460 358544 449472
rect 335326 449432 358544 449460
rect 304350 449284 304356 449336
rect 304408 449324 304414 449336
rect 335326 449324 335354 449432
rect 358538 449420 358544 449432
rect 358596 449420 358602 449472
rect 365070 449460 365076 449472
rect 358648 449432 365076 449460
rect 341702 449352 341708 449404
rect 341760 449392 341766 449404
rect 344094 449392 344100 449404
rect 341760 449364 344100 449392
rect 341760 449352 341766 449364
rect 344094 449352 344100 449364
rect 344152 449352 344158 449404
rect 348510 449352 348516 449404
rect 348568 449352 348574 449404
rect 358648 449392 358676 449432
rect 365070 449420 365076 449432
rect 365128 449420 365134 449472
rect 369854 449420 369860 449472
rect 369912 449460 369918 449472
rect 370590 449460 370596 449472
rect 369912 449432 370596 449460
rect 369912 449420 369918 449432
rect 370590 449420 370596 449432
rect 370648 449420 370654 449472
rect 354646 449364 358676 449392
rect 304408 449296 335354 449324
rect 304408 449284 304414 449296
rect 342438 449284 342444 449336
rect 342496 449324 342502 449336
rect 348528 449324 348556 449352
rect 342496 449296 348556 449324
rect 342496 449284 342502 449296
rect 305638 449216 305644 449268
rect 305696 449256 305702 449268
rect 309042 449256 309048 449268
rect 305696 449228 309048 449256
rect 305696 449216 305702 449228
rect 309042 449216 309048 449228
rect 309100 449256 309106 449268
rect 354646 449256 354674 449364
rect 362218 449352 362224 449404
rect 362276 449352 362282 449404
rect 362236 449324 362264 449352
rect 309100 449228 354674 449256
rect 358464 449296 362264 449324
rect 309100 449216 309106 449228
rect 88334 449148 88340 449200
rect 88392 449188 88398 449200
rect 309134 449188 309140 449200
rect 88392 449160 309140 449188
rect 88392 449148 88398 449160
rect 309134 449148 309140 449160
rect 309192 449188 309198 449200
rect 358464 449188 358492 449296
rect 309192 449160 358492 449188
rect 309192 449148 309198 449160
rect 3050 448604 3056 448656
rect 3108 448644 3114 448656
rect 281534 448644 281540 448656
rect 3108 448616 281540 448644
rect 3108 448604 3114 448616
rect 281534 448604 281540 448616
rect 281592 448604 281598 448656
rect 282822 448604 282828 448656
rect 282880 448644 282886 448656
rect 342438 448644 342444 448656
rect 282880 448616 342444 448644
rect 282880 448604 282886 448616
rect 342438 448604 342444 448616
rect 342496 448604 342502 448656
rect 281166 448536 281172 448588
rect 281224 448576 281230 448588
rect 342346 448576 342352 448588
rect 281224 448548 342352 448576
rect 281224 448536 281230 448548
rect 342346 448536 342352 448548
rect 342404 448536 342410 448588
rect 322474 445000 322480 445052
rect 322532 445040 322538 445052
rect 340966 445040 340972 445052
rect 322532 445012 340972 445040
rect 322532 445000 322538 445012
rect 340966 445000 340972 445012
rect 341024 445000 341030 445052
rect 311158 443640 311164 443692
rect 311216 443680 311222 443692
rect 340874 443680 340880 443692
rect 311216 443652 340880 443680
rect 311216 443640 311222 443652
rect 340874 443640 340880 443652
rect 340932 443640 340938 443692
rect 289722 438132 289728 438184
rect 289780 438172 289786 438184
rect 340966 438172 340972 438184
rect 289780 438144 340972 438172
rect 289780 438132 289786 438144
rect 340966 438132 340972 438144
rect 341024 438132 341030 438184
rect 319622 436704 319628 436756
rect 319680 436744 319686 436756
rect 340966 436744 340972 436756
rect 319680 436716 340972 436744
rect 319680 436704 319686 436716
rect 340966 436704 340972 436716
rect 341024 436704 341030 436756
rect 389818 431876 389824 431928
rect 389876 431916 389882 431928
rect 580166 431916 580172 431928
rect 389876 431888 580172 431916
rect 389876 431876 389882 431888
rect 580166 431876 580172 431888
rect 580224 431876 580230 431928
rect 284938 428408 284944 428460
rect 284996 428448 285002 428460
rect 340966 428448 340972 428460
rect 284996 428420 340972 428448
rect 284996 428408 285002 428420
rect 340966 428408 340972 428420
rect 341024 428408 341030 428460
rect 288342 424328 288348 424380
rect 288400 424368 288406 424380
rect 340322 424368 340328 424380
rect 288400 424340 340328 424368
rect 288400 424328 288406 424340
rect 340322 424328 340328 424340
rect 340380 424328 340386 424380
rect 3510 422288 3516 422340
rect 3568 422328 3574 422340
rect 315574 422328 315580 422340
rect 3568 422300 315580 422328
rect 3568 422288 3574 422300
rect 315574 422288 315580 422300
rect 315632 422328 315638 422340
rect 316770 422328 316776 422340
rect 315632 422300 316776 422328
rect 315632 422288 315638 422300
rect 316770 422288 316776 422300
rect 316828 422288 316834 422340
rect 8938 421540 8944 421592
rect 8996 421580 9002 421592
rect 314654 421580 314660 421592
rect 8996 421552 314660 421580
rect 8996 421540 9002 421552
rect 314654 421540 314660 421552
rect 314712 421540 314718 421592
rect 314654 420860 314660 420912
rect 314712 420900 314718 420912
rect 315390 420900 315396 420912
rect 314712 420872 315396 420900
rect 314712 420860 314718 420872
rect 315390 420860 315396 420872
rect 315448 420900 315454 420912
rect 334894 420900 334900 420912
rect 315448 420872 334900 420900
rect 315448 420860 315454 420872
rect 334894 420860 334900 420872
rect 334952 420860 334958 420912
rect 3418 420180 3424 420232
rect 3476 420220 3482 420232
rect 311894 420220 311900 420232
rect 3476 420192 311900 420220
rect 3476 420180 3482 420192
rect 311894 420180 311900 420192
rect 311952 420180 311958 420232
rect 7558 419432 7564 419484
rect 7616 419472 7622 419484
rect 311158 419472 311164 419484
rect 7616 419444 311164 419472
rect 7616 419432 7622 419444
rect 311158 419432 311164 419444
rect 311216 419432 311222 419484
rect 311894 419432 311900 419484
rect 311952 419472 311958 419484
rect 312630 419472 312636 419484
rect 311952 419444 312636 419472
rect 311952 419432 311958 419444
rect 312630 419432 312636 419444
rect 312688 419472 312694 419484
rect 337654 419472 337660 419484
rect 312688 419444 337660 419472
rect 312688 419432 312694 419444
rect 337654 419432 337660 419444
rect 337712 419432 337718 419484
rect 310698 418140 310704 418192
rect 310756 418180 310762 418192
rect 311158 418180 311164 418192
rect 310756 418152 311164 418180
rect 310756 418140 310762 418152
rect 311158 418140 311164 418152
rect 311216 418140 311222 418192
rect 10318 418072 10324 418124
rect 10376 418112 10382 418124
rect 313550 418112 313556 418124
rect 10376 418084 313556 418112
rect 10376 418072 10382 418084
rect 313550 418072 313556 418084
rect 313608 418072 313614 418124
rect 313550 417664 313556 417716
rect 313608 417704 313614 417716
rect 314010 417704 314016 417716
rect 313608 417676 314016 417704
rect 313608 417664 313614 417676
rect 314010 417664 314016 417676
rect 314068 417664 314074 417716
rect 142798 416032 142804 416084
rect 142856 416072 142862 416084
rect 312722 416072 312728 416084
rect 142856 416044 312728 416072
rect 142856 416032 142862 416044
rect 312722 416032 312728 416044
rect 312780 416032 312786 416084
rect 4798 414672 4804 414724
rect 4856 414712 4862 414724
rect 310514 414712 310520 414724
rect 4856 414684 310520 414712
rect 4856 414672 4862 414684
rect 310514 414672 310520 414684
rect 310572 414672 310578 414724
rect 310514 413924 310520 413976
rect 310572 413964 310578 413976
rect 337470 413964 337476 413976
rect 310572 413936 337476 413964
rect 310572 413924 310578 413936
rect 337470 413924 337476 413936
rect 337528 413924 337534 413976
rect 71774 411884 71780 411936
rect 71832 411924 71838 411936
rect 308122 411924 308128 411936
rect 71832 411896 308128 411924
rect 71832 411884 71838 411896
rect 308122 411884 308128 411896
rect 308180 411884 308186 411936
rect 308122 411204 308128 411256
rect 308180 411244 308186 411256
rect 309042 411244 309048 411256
rect 308180 411216 309048 411244
rect 308180 411204 308186 411216
rect 309042 411204 309048 411216
rect 309100 411244 309106 411256
rect 340230 411244 340236 411256
rect 309100 411216 340236 411244
rect 309100 411204 309106 411216
rect 340230 411204 340236 411216
rect 340288 411204 340294 411256
rect 282914 409164 282920 409216
rect 282972 409204 282978 409216
rect 304994 409204 305000 409216
rect 282972 409176 305000 409204
rect 282972 409164 282978 409176
rect 304994 409164 305000 409176
rect 305052 409164 305058 409216
rect 293218 409096 293224 409148
rect 293276 409136 293282 409148
rect 338758 409136 338764 409148
rect 293276 409108 338764 409136
rect 293276 409096 293282 409108
rect 338758 409096 338764 409108
rect 338816 409096 338822 409148
rect 23474 407736 23480 407788
rect 23532 407776 23538 407788
rect 310422 407776 310428 407788
rect 23532 407748 310428 407776
rect 23532 407736 23538 407748
rect 310422 407736 310428 407748
rect 310480 407736 310486 407788
rect 325142 407736 325148 407788
rect 325200 407776 325206 407788
rect 340138 407776 340144 407788
rect 325200 407748 340144 407776
rect 325200 407736 325206 407748
rect 340138 407736 340144 407748
rect 340196 407736 340202 407788
rect 3418 407056 3424 407108
rect 3476 407096 3482 407108
rect 316218 407096 316224 407108
rect 3476 407068 316224 407096
rect 3476 407056 3482 407068
rect 316218 407056 316224 407068
rect 316276 407096 316282 407108
rect 316862 407096 316868 407108
rect 316276 407068 316868 407096
rect 316276 407056 316282 407068
rect 316862 407056 316868 407068
rect 316920 407056 316926 407108
rect 309870 406988 309876 407040
rect 309928 407028 309934 407040
rect 310422 407028 310428 407040
rect 309928 407000 310428 407028
rect 309928 406988 309934 407000
rect 310422 406988 310428 407000
rect 310480 407028 310486 407040
rect 334802 407028 334808 407040
rect 310480 407000 334808 407028
rect 310480 406988 310486 407000
rect 334802 406988 334808 407000
rect 334860 406988 334866 407040
rect 292022 406376 292028 406428
rect 292080 406416 292086 406428
rect 337378 406416 337384 406428
rect 292080 406388 337384 406416
rect 292080 406376 292086 406388
rect 337378 406376 337384 406388
rect 337436 406376 337442 406428
rect 304994 405628 305000 405680
rect 305052 405668 305058 405680
rect 305730 405668 305736 405680
rect 305052 405640 305736 405668
rect 305052 405628 305058 405640
rect 305730 405628 305736 405640
rect 305788 405668 305794 405680
rect 340966 405668 340972 405680
rect 305788 405640 340972 405668
rect 305788 405628 305794 405640
rect 340966 405628 340972 405640
rect 341024 405628 341030 405680
rect 388990 405628 388996 405680
rect 389048 405668 389054 405680
rect 580166 405668 580172 405680
rect 389048 405640 580172 405668
rect 389048 405628 389054 405640
rect 580166 405628 580172 405640
rect 580224 405628 580230 405680
rect 195238 404948 195244 405000
rect 195296 404988 195302 405000
rect 314010 404988 314016 405000
rect 195296 404960 314016 404988
rect 195296 404948 195302 404960
rect 314010 404948 314016 404960
rect 314068 404948 314074 405000
rect 281534 404268 281540 404320
rect 281592 404308 281598 404320
rect 281994 404308 282000 404320
rect 281592 404280 282000 404308
rect 281592 404268 281598 404280
rect 281994 404268 282000 404280
rect 282052 404308 282058 404320
rect 315298 404308 315304 404320
rect 282052 404280 315304 404308
rect 282052 404268 282058 404280
rect 315298 404268 315304 404280
rect 315356 404268 315362 404320
rect 314010 404200 314016 404252
rect 314068 404240 314074 404252
rect 334710 404240 334716 404252
rect 314068 404212 334716 404240
rect 314068 404200 314074 404212
rect 334710 404200 334716 404212
rect 334768 404200 334774 404252
rect 13078 403588 13084 403640
rect 13136 403628 13142 403640
rect 220170 403628 220176 403640
rect 13136 403600 220176 403628
rect 13136 403588 13142 403600
rect 220170 403588 220176 403600
rect 220228 403588 220234 403640
rect 255958 403588 255964 403640
rect 256016 403628 256022 403640
rect 281994 403628 282000 403640
rect 256016 403600 282000 403628
rect 256016 403588 256022 403600
rect 281994 403588 282000 403600
rect 282052 403588 282058 403640
rect 220170 402976 220176 403028
rect 220228 403016 220234 403028
rect 315482 403016 315488 403028
rect 220228 402988 315488 403016
rect 220228 402976 220234 402988
rect 315482 402976 315488 402988
rect 315540 402976 315546 403028
rect 298738 402908 298744 402960
rect 298796 402948 298802 402960
rect 313918 402948 313924 402960
rect 298796 402920 313924 402948
rect 298796 402908 298802 402920
rect 313918 402908 313924 402920
rect 313976 402908 313982 402960
rect 315574 402840 315580 402892
rect 315632 402880 315638 402892
rect 316126 402880 316132 402892
rect 315632 402852 316132 402880
rect 315632 402840 315638 402852
rect 316126 402840 316132 402852
rect 316184 402840 316190 402892
rect 313366 402228 313372 402280
rect 313424 402268 313430 402280
rect 313918 402268 313924 402280
rect 313424 402240 313924 402268
rect 313424 402228 313430 402240
rect 313918 402228 313924 402240
rect 313976 402228 313982 402280
rect 341886 400936 341892 400988
rect 341944 400976 341950 400988
rect 341944 400948 347084 400976
rect 341944 400936 341950 400948
rect 347056 400704 347084 400948
rect 343790 400676 344922 400704
rect 347056 400676 353294 400704
rect 341702 400636 341708 400648
rect 335326 400608 341708 400636
rect 333330 400528 333336 400580
rect 333388 400568 333394 400580
rect 335326 400568 335354 400608
rect 341702 400596 341708 400608
rect 341760 400596 341766 400648
rect 343790 400636 343818 400676
rect 341996 400608 343818 400636
rect 333388 400540 335354 400568
rect 333388 400528 333394 400540
rect 336182 400460 336188 400512
rect 336240 400500 336246 400512
rect 341996 400500 342024 400608
rect 344894 400568 344922 400676
rect 353266 400636 353294 400676
rect 353266 400608 361942 400636
rect 344894 400540 361850 400568
rect 336240 400472 342024 400500
rect 342088 400472 358354 400500
rect 336240 400460 336246 400472
rect 282086 400392 282092 400444
rect 282144 400432 282150 400444
rect 333882 400432 333888 400444
rect 282144 400404 333888 400432
rect 282144 400392 282150 400404
rect 333882 400392 333888 400404
rect 333940 400392 333946 400444
rect 341794 400392 341800 400444
rect 341852 400432 341858 400444
rect 342088 400432 342116 400472
rect 341852 400404 342116 400432
rect 341852 400392 341858 400404
rect 342254 400392 342260 400444
rect 342312 400432 342318 400444
rect 342312 400404 356330 400432
rect 342312 400392 342318 400404
rect 279970 400324 279976 400376
rect 280028 400364 280034 400376
rect 280028 400336 346532 400364
rect 280028 400324 280034 400336
rect 274450 400256 274456 400308
rect 274508 400296 274514 400308
rect 346504 400296 346532 400336
rect 274508 400268 346440 400296
rect 346504 400268 352558 400296
rect 274508 400256 274514 400268
rect 275830 400188 275836 400240
rect 275888 400228 275894 400240
rect 342254 400228 342260 400240
rect 275888 400200 342260 400228
rect 275888 400188 275894 400200
rect 342254 400188 342260 400200
rect 342312 400188 342318 400240
rect 346412 400228 346440 400268
rect 342364 400200 345014 400228
rect 346412 400200 352466 400228
rect 333882 400120 333888 400172
rect 333940 400160 333946 400172
rect 342364 400160 342392 400200
rect 333940 400132 342392 400160
rect 344986 400160 345014 400200
rect 344986 400132 345290 400160
rect 333940 400120 333946 400132
rect 342070 400052 342076 400104
rect 342128 400092 342134 400104
rect 342254 400092 342260 400104
rect 342128 400064 342260 400092
rect 342128 400052 342134 400064
rect 342254 400052 342260 400064
rect 342312 400052 342318 400104
rect 343606 400064 344738 400092
rect 343606 400024 343634 400064
rect 322906 399996 343634 400024
rect 273162 399644 273168 399696
rect 273220 399684 273226 399696
rect 322906 399684 322934 399996
rect 334342 399916 334348 399968
rect 334400 399956 334406 399968
rect 334400 399928 343082 399956
rect 334400 399916 334406 399928
rect 343054 399900 343082 399928
rect 343422 399928 344186 399956
rect 327534 399848 327540 399900
rect 327592 399888 327598 399900
rect 342852 399888 342858 399900
rect 327592 399860 342858 399888
rect 327592 399848 327598 399860
rect 342852 399848 342858 399860
rect 342910 399848 342916 399900
rect 343036 399848 343042 399900
rect 343094 399848 343100 399900
rect 343312 399848 343318 399900
rect 343370 399848 343376 399900
rect 335814 399780 335820 399832
rect 335872 399820 335878 399832
rect 342944 399820 342950 399832
rect 335872 399792 342950 399820
rect 335872 399780 335878 399792
rect 342944 399780 342950 399792
rect 343002 399780 343008 399832
rect 334894 399712 334900 399764
rect 334952 399752 334958 399764
rect 343330 399752 343358 399848
rect 334952 399724 343358 399752
rect 334952 399712 334958 399724
rect 273220 399656 322934 399684
rect 273220 399644 273226 399656
rect 335630 399644 335636 399696
rect 335688 399684 335694 399696
rect 343422 399684 343450 399928
rect 344158 399900 344186 399928
rect 344710 399900 344738 400064
rect 345262 399900 345290 400132
rect 347056 399928 348326 399956
rect 343864 399848 343870 399900
rect 343922 399848 343928 399900
rect 343956 399848 343962 399900
rect 344014 399848 344020 399900
rect 344140 399848 344146 399900
rect 344198 399848 344204 399900
rect 344324 399848 344330 399900
rect 344382 399848 344388 399900
rect 344692 399848 344698 399900
rect 344750 399848 344756 399900
rect 344876 399848 344882 399900
rect 344934 399848 344940 399900
rect 345244 399848 345250 399900
rect 345302 399848 345308 399900
rect 345520 399848 345526 399900
rect 345578 399848 345584 399900
rect 345796 399848 345802 399900
rect 345854 399848 345860 399900
rect 346072 399848 346078 399900
rect 346130 399848 346136 399900
rect 346256 399848 346262 399900
rect 346314 399848 346320 399900
rect 346440 399848 346446 399900
rect 346498 399848 346504 399900
rect 346532 399848 346538 399900
rect 346590 399888 346596 399900
rect 346590 399860 346716 399888
rect 346590 399848 346596 399860
rect 343496 399780 343502 399832
rect 343554 399780 343560 399832
rect 343772 399820 343778 399832
rect 343606 399792 343778 399820
rect 343514 399696 343542 399780
rect 335688 399656 343450 399684
rect 335688 399644 335694 399656
rect 343496 399644 343502 399696
rect 343554 399644 343560 399696
rect 262122 399576 262128 399628
rect 262180 399616 262186 399628
rect 342070 399616 342076 399628
rect 262180 399588 342076 399616
rect 262180 399576 262186 399588
rect 342070 399576 342076 399588
rect 342128 399576 342134 399628
rect 342254 399576 342260 399628
rect 342312 399616 342318 399628
rect 343606 399616 343634 399792
rect 343772 399780 343778 399792
rect 343830 399780 343836 399832
rect 343680 399712 343686 399764
rect 343738 399712 343744 399764
rect 342312 399588 343634 399616
rect 342312 399576 342318 399588
rect 311158 399508 311164 399560
rect 311216 399548 311222 399560
rect 341886 399548 341892 399560
rect 311216 399520 341892 399548
rect 311216 399508 311222 399520
rect 341886 399508 341892 399520
rect 341944 399508 341950 399560
rect 341978 399508 341984 399560
rect 342036 399548 342042 399560
rect 343698 399548 343726 399712
rect 342036 399520 343726 399548
rect 343882 399560 343910 399848
rect 343974 399764 344002 399848
rect 344048 399780 344054 399832
rect 344106 399780 344112 399832
rect 343956 399712 343962 399764
rect 344014 399712 344020 399764
rect 344066 399684 344094 399780
rect 344342 399696 344370 399848
rect 344894 399696 344922 399848
rect 344020 399656 344094 399684
rect 344020 399628 344048 399656
rect 344278 399644 344284 399696
rect 344336 399656 344370 399696
rect 344336 399644 344342 399656
rect 344830 399644 344836 399696
rect 344888 399656 344922 399696
rect 344888 399644 344894 399656
rect 344002 399576 344008 399628
rect 344060 399576 344066 399628
rect 344094 399576 344100 399628
rect 344152 399616 344158 399628
rect 344738 399616 344744 399628
rect 344152 399588 344744 399616
rect 344152 399576 344158 399588
rect 344738 399576 344744 399588
rect 344796 399576 344802 399628
rect 345382 399576 345388 399628
rect 345440 399616 345446 399628
rect 345538 399616 345566 399848
rect 345704 399820 345710 399832
rect 345440 399588 345566 399616
rect 345630 399792 345710 399820
rect 345440 399576 345446 399588
rect 343882 399520 343916 399560
rect 342036 399508 342042 399520
rect 343910 399508 343916 399520
rect 343968 399508 343974 399560
rect 344554 399508 344560 399560
rect 344612 399548 344618 399560
rect 345630 399548 345658 399792
rect 345704 399780 345710 399792
rect 345762 399780 345768 399832
rect 345814 399628 345842 399848
rect 346090 399684 346118 399848
rect 346164 399780 346170 399832
rect 346222 399780 346228 399832
rect 345952 399656 346118 399684
rect 345952 399628 345980 399656
rect 346182 399628 346210 399780
rect 345750 399576 345756 399628
rect 345808 399588 345842 399628
rect 345808 399576 345814 399588
rect 345934 399576 345940 399628
rect 345992 399576 345998 399628
rect 346118 399576 346124 399628
rect 346176 399588 346210 399628
rect 346274 399628 346302 399848
rect 346458 399764 346486 399848
rect 346458 399724 346492 399764
rect 346486 399712 346492 399724
rect 346544 399712 346550 399764
rect 346274 399588 346308 399628
rect 346176 399576 346182 399588
rect 346302 399576 346308 399588
rect 346360 399576 346366 399628
rect 346688 399616 346716 399860
rect 346900 399848 346906 399900
rect 346958 399848 346964 399900
rect 346918 399628 346946 399848
rect 347056 399696 347084 399928
rect 348298 399900 348326 399928
rect 352438 399900 352466 400200
rect 352530 400024 352558 400268
rect 352530 399996 353386 400024
rect 347452 399848 347458 399900
rect 347510 399848 347516 399900
rect 347636 399848 347642 399900
rect 347694 399848 347700 399900
rect 348004 399848 348010 399900
rect 348062 399848 348068 399900
rect 348280 399848 348286 399900
rect 348338 399848 348344 399900
rect 349568 399848 349574 399900
rect 349626 399848 349632 399900
rect 349660 399848 349666 399900
rect 349718 399848 349724 399900
rect 349752 399848 349758 399900
rect 349810 399848 349816 399900
rect 349936 399848 349942 399900
rect 349994 399848 350000 399900
rect 350304 399848 350310 399900
rect 350362 399848 350368 399900
rect 350580 399848 350586 399900
rect 350638 399848 350644 399900
rect 350764 399848 350770 399900
rect 350822 399848 350828 399900
rect 351040 399848 351046 399900
rect 351098 399848 351104 399900
rect 351132 399848 351138 399900
rect 351190 399848 351196 399900
rect 351224 399848 351230 399900
rect 351282 399888 351288 399900
rect 351282 399848 351316 399888
rect 351408 399848 351414 399900
rect 351466 399848 351472 399900
rect 351684 399888 351690 399900
rect 351656 399848 351690 399888
rect 351742 399848 351748 399900
rect 352052 399848 352058 399900
rect 352110 399848 352116 399900
rect 352236 399848 352242 399900
rect 352294 399848 352300 399900
rect 352420 399848 352426 399900
rect 352478 399848 352484 399900
rect 352788 399848 352794 399900
rect 352846 399848 352852 399900
rect 352972 399888 352978 399900
rect 352944 399848 352978 399888
rect 353030 399848 353036 399900
rect 353358 399888 353386 399996
rect 353726 399928 355502 399956
rect 353726 399888 353754 399928
rect 355474 399900 355502 399928
rect 356302 399900 356330 400404
rect 358326 400228 358354 400472
rect 358878 400336 360470 400364
rect 358878 400228 358906 400336
rect 358326 400200 358906 400228
rect 357544 399928 358170 399956
rect 353358 399860 353754 399888
rect 353892 399848 353898 399900
rect 353950 399848 353956 399900
rect 354076 399848 354082 399900
rect 354134 399848 354140 399900
rect 354260 399848 354266 399900
rect 354318 399888 354324 399900
rect 354318 399860 354582 399888
rect 354318 399848 354324 399860
rect 347268 399780 347274 399832
rect 347326 399780 347332 399832
rect 347038 399644 347044 399696
rect 347096 399644 347102 399696
rect 347286 399628 347314 399780
rect 347470 399696 347498 399848
rect 347470 399656 347504 399696
rect 347498 399644 347504 399656
rect 347556 399644 347562 399696
rect 346762 399616 346768 399628
rect 346688 399588 346768 399616
rect 346762 399576 346768 399588
rect 346820 399576 346826 399628
rect 346918 399588 346952 399628
rect 346946 399576 346952 399588
rect 347004 399576 347010 399628
rect 347286 399588 347320 399628
rect 347314 399576 347320 399588
rect 347372 399576 347378 399628
rect 344612 399520 345658 399548
rect 344612 399508 344618 399520
rect 281442 399440 281448 399492
rect 281500 399480 281506 399492
rect 347222 399480 347228 399492
rect 281500 399452 347228 399480
rect 281500 399440 281506 399452
rect 347222 399440 347228 399452
rect 347280 399440 347286 399492
rect 347654 399424 347682 399848
rect 347866 399576 347872 399628
rect 347924 399616 347930 399628
rect 348022 399616 348050 399848
rect 348096 399780 348102 399832
rect 348154 399780 348160 399832
rect 348188 399780 348194 399832
rect 348246 399780 348252 399832
rect 348372 399780 348378 399832
rect 348430 399780 348436 399832
rect 347924 399588 348050 399616
rect 348114 399628 348142 399780
rect 348206 399696 348234 399780
rect 348206 399656 348240 399696
rect 348234 399644 348240 399656
rect 348292 399644 348298 399696
rect 348114 399588 348148 399628
rect 347924 399576 347930 399588
rect 348142 399576 348148 399588
rect 348200 399576 348206 399628
rect 348050 399440 348056 399492
rect 348108 399480 348114 399492
rect 348390 399480 348418 399780
rect 349586 399616 349614 399848
rect 348108 399452 348418 399480
rect 349356 399588 349614 399616
rect 349356 399480 349384 399588
rect 349430 399508 349436 399560
rect 349488 399548 349494 399560
rect 349678 399548 349706 399848
rect 349770 399696 349798 399848
rect 349770 399656 349804 399696
rect 349798 399644 349804 399656
rect 349856 399644 349862 399696
rect 349488 399520 349706 399548
rect 349488 399508 349494 399520
rect 349954 399492 349982 399848
rect 350028 399780 350034 399832
rect 350086 399780 350092 399832
rect 350322 399820 350350 399848
rect 350184 399792 350350 399820
rect 350046 399548 350074 399780
rect 350046 399520 350120 399548
rect 349614 399480 349620 399492
rect 349356 399452 349620 399480
rect 348108 399440 348114 399452
rect 349614 399440 349620 399452
rect 349672 399440 349678 399492
rect 349954 399452 349988 399492
rect 349982 399440 349988 399452
rect 350040 399440 350046 399492
rect 336274 399372 336280 399424
rect 336332 399412 336338 399424
rect 341794 399412 341800 399424
rect 336332 399384 341800 399412
rect 336332 399372 336338 399384
rect 341794 399372 341800 399384
rect 341852 399372 341858 399424
rect 342254 399372 342260 399424
rect 342312 399412 342318 399424
rect 346394 399412 346400 399424
rect 342312 399384 346400 399412
rect 342312 399372 342318 399384
rect 346394 399372 346400 399384
rect 346452 399372 346458 399424
rect 347654 399384 347688 399424
rect 347682 399372 347688 399384
rect 347740 399372 347746 399424
rect 349890 399372 349896 399424
rect 349948 399412 349954 399424
rect 350092 399412 350120 399520
rect 349948 399384 350120 399412
rect 349948 399372 349954 399384
rect 334710 399304 334716 399356
rect 334768 399344 334774 399356
rect 345658 399344 345664 399356
rect 334768 399316 345664 399344
rect 334768 399304 334774 399316
rect 345658 399304 345664 399316
rect 345716 399304 345722 399356
rect 346090 399316 347084 399344
rect 333790 399236 333796 399288
rect 333848 399276 333854 399288
rect 346090 399276 346118 399316
rect 333848 399248 346118 399276
rect 333848 399236 333854 399248
rect 340046 399168 340052 399220
rect 340104 399208 340110 399220
rect 344554 399208 344560 399220
rect 340104 399180 344560 399208
rect 340104 399168 340110 399180
rect 344554 399168 344560 399180
rect 344612 399168 344618 399220
rect 347056 399208 347084 399316
rect 348694 399304 348700 399356
rect 348752 399344 348758 399356
rect 350184 399344 350212 399792
rect 350396 399780 350402 399832
rect 350454 399780 350460 399832
rect 350414 399752 350442 399780
rect 350276 399724 350442 399752
rect 350276 399424 350304 399724
rect 350598 399684 350626 399848
rect 350672 399780 350678 399832
rect 350730 399780 350736 399832
rect 350460 399656 350626 399684
rect 350690 399696 350718 399780
rect 350782 399764 350810 399848
rect 350948 399780 350954 399832
rect 351006 399780 351012 399832
rect 350782 399724 350816 399764
rect 350810 399712 350816 399724
rect 350868 399712 350874 399764
rect 350966 399696 350994 399780
rect 350690 399656 350724 399696
rect 350460 399628 350488 399656
rect 350718 399644 350724 399656
rect 350776 399644 350782 399696
rect 350902 399644 350908 399696
rect 350960 399656 350994 399696
rect 350960 399644 350966 399656
rect 350442 399576 350448 399628
rect 350500 399576 350506 399628
rect 350626 399576 350632 399628
rect 350684 399616 350690 399628
rect 351058 399616 351086 399848
rect 351150 399696 351178 399848
rect 351150 399656 351184 399696
rect 351178 399644 351184 399656
rect 351236 399644 351242 399696
rect 351288 399628 351316 399848
rect 351426 399628 351454 399848
rect 351656 399764 351684 399848
rect 351638 399712 351644 399764
rect 351696 399712 351702 399764
rect 350684 399588 351086 399616
rect 350684 399576 350690 399588
rect 351270 399576 351276 399628
rect 351328 399576 351334 399628
rect 351426 399588 351460 399628
rect 351454 399576 351460 399588
rect 351512 399576 351518 399628
rect 352070 399424 352098 399848
rect 352254 399548 352282 399848
rect 352374 399548 352380 399560
rect 352254 399520 352380 399548
rect 352374 399508 352380 399520
rect 352432 399508 352438 399560
rect 352806 399480 352834 399848
rect 352944 399628 352972 399848
rect 353754 399644 353760 399696
rect 353812 399684 353818 399696
rect 353910 399684 353938 399848
rect 353812 399656 353938 399684
rect 354094 399684 354122 399848
rect 354398 399684 354404 399696
rect 354094 399656 354404 399684
rect 353812 399644 353818 399656
rect 354398 399644 354404 399656
rect 354456 399644 354462 399696
rect 352926 399576 352932 399628
rect 352984 399576 352990 399628
rect 354030 399576 354036 399628
rect 354088 399616 354094 399628
rect 354554 399616 354582 399860
rect 355456 399848 355462 399900
rect 355514 399848 355520 399900
rect 355732 399848 355738 399900
rect 355790 399848 355796 399900
rect 356284 399848 356290 399900
rect 356342 399848 356348 399900
rect 356468 399848 356474 399900
rect 356526 399848 356532 399900
rect 356560 399848 356566 399900
rect 356618 399848 356624 399900
rect 356744 399848 356750 399900
rect 356802 399848 356808 399900
rect 357296 399848 357302 399900
rect 357354 399848 357360 399900
rect 357388 399848 357394 399900
rect 357446 399848 357452 399900
rect 354088 399588 354582 399616
rect 354088 399576 354094 399588
rect 355750 399560 355778 399848
rect 356100 399780 356106 399832
rect 356158 399780 356164 399832
rect 356486 399820 356514 399848
rect 356440 399792 356514 399820
rect 356118 399752 356146 399780
rect 356118 399724 356192 399752
rect 356164 399696 356192 399724
rect 356440 399696 356468 399792
rect 356578 399764 356606 399848
rect 356514 399712 356520 399764
rect 356572 399724 356606 399764
rect 356572 399712 356578 399724
rect 356762 399696 356790 399848
rect 356928 399780 356934 399832
rect 356986 399780 356992 399832
rect 356146 399644 356152 399696
rect 356204 399644 356210 399696
rect 356422 399644 356428 399696
rect 356480 399644 356486 399696
rect 356762 399656 356796 399696
rect 356790 399644 356796 399656
rect 356848 399644 356854 399696
rect 356946 399684 356974 399780
rect 356900 399656 356974 399684
rect 355226 399508 355232 399560
rect 355284 399548 355290 399560
rect 355410 399548 355416 399560
rect 355284 399520 355416 399548
rect 355284 399508 355290 399520
rect 355410 399508 355416 399520
rect 355468 399508 355474 399560
rect 355686 399508 355692 399560
rect 355744 399520 355778 399560
rect 355744 399508 355750 399520
rect 355962 399508 355968 399560
rect 356020 399548 356026 399560
rect 356900 399548 356928 399656
rect 357158 399576 357164 399628
rect 357216 399616 357222 399628
rect 357314 399616 357342 399848
rect 357216 399588 357342 399616
rect 357216 399576 357222 399588
rect 356020 399520 356928 399548
rect 356020 399508 356026 399520
rect 352530 399452 352834 399480
rect 352530 399424 352558 399452
rect 353570 399440 353576 399492
rect 353628 399480 353634 399492
rect 353628 399452 354904 399480
rect 353628 399440 353634 399452
rect 350258 399372 350264 399424
rect 350316 399372 350322 399424
rect 352070 399384 352104 399424
rect 352098 399372 352104 399384
rect 352156 399372 352162 399424
rect 352466 399372 352472 399424
rect 352524 399384 352558 399424
rect 352524 399372 352530 399384
rect 354214 399372 354220 399424
rect 354272 399412 354278 399424
rect 354766 399412 354772 399424
rect 354272 399384 354772 399412
rect 354272 399372 354278 399384
rect 354766 399372 354772 399384
rect 354824 399372 354830 399424
rect 354876 399412 354904 399452
rect 357250 399440 357256 399492
rect 357308 399480 357314 399492
rect 357406 399480 357434 399848
rect 357544 399628 357572 399928
rect 358142 399900 358170 399928
rect 360442 399900 360470 400336
rect 361822 399900 361850 400540
rect 361914 400228 361942 400608
rect 387518 400364 387524 400376
rect 374334 400336 387524 400364
rect 361914 400200 365714 400228
rect 365686 400160 365714 400200
rect 367066 400200 370314 400228
rect 367066 400160 367094 400200
rect 365686 400132 367094 400160
rect 366238 399928 366542 399956
rect 366238 399900 366266 399928
rect 357664 399848 357670 399900
rect 357722 399848 357728 399900
rect 357940 399848 357946 399900
rect 357998 399848 358004 399900
rect 358124 399848 358130 399900
rect 358182 399848 358188 399900
rect 358676 399848 358682 399900
rect 358734 399848 358740 399900
rect 358952 399848 358958 399900
rect 359010 399848 359016 399900
rect 359136 399848 359142 399900
rect 359194 399848 359200 399900
rect 359228 399848 359234 399900
rect 359286 399848 359292 399900
rect 359872 399848 359878 399900
rect 359930 399848 359936 399900
rect 359964 399848 359970 399900
rect 360022 399888 360028 399900
rect 360022 399848 360056 399888
rect 360240 399848 360246 399900
rect 360298 399848 360304 399900
rect 360332 399848 360338 399900
rect 360390 399848 360396 399900
rect 360424 399848 360430 399900
rect 360482 399848 360488 399900
rect 360516 399848 360522 399900
rect 360574 399888 360580 399900
rect 360574 399860 360838 399888
rect 360574 399848 360580 399860
rect 357526 399576 357532 399628
rect 357584 399576 357590 399628
rect 357682 399560 357710 399848
rect 357756 399780 357762 399832
rect 357814 399780 357820 399832
rect 357774 399628 357802 399780
rect 357774 399588 357808 399628
rect 357802 399576 357808 399588
rect 357860 399576 357866 399628
rect 357958 399616 357986 399848
rect 358308 399780 358314 399832
rect 358366 399780 358372 399832
rect 358326 399696 358354 399780
rect 358326 399656 358360 399696
rect 358354 399644 358360 399656
rect 358412 399644 358418 399696
rect 358262 399616 358268 399628
rect 357958 399588 358268 399616
rect 358262 399576 358268 399588
rect 358320 399576 358326 399628
rect 357618 399508 357624 399560
rect 357676 399520 357710 399560
rect 357676 399508 357682 399520
rect 357308 399452 357434 399480
rect 358694 399492 358722 399848
rect 358970 399628 358998 399848
rect 358970 399588 359004 399628
rect 358998 399576 359004 399588
rect 359056 399576 359062 399628
rect 359154 399616 359182 399848
rect 359246 399752 359274 399848
rect 359688 399780 359694 399832
rect 359746 399780 359752 399832
rect 359246 399724 359504 399752
rect 359274 399616 359280 399628
rect 359154 399588 359280 399616
rect 359274 399576 359280 399588
rect 359332 399576 359338 399628
rect 359182 399508 359188 399560
rect 359240 399548 359246 399560
rect 359476 399548 359504 399724
rect 359706 399684 359734 399780
rect 359240 399520 359504 399548
rect 359660 399656 359734 399684
rect 359240 399508 359246 399520
rect 359660 399492 359688 399656
rect 359734 399576 359740 399628
rect 359792 399616 359798 399628
rect 359890 399616 359918 399848
rect 360028 399764 360056 399848
rect 360010 399712 360016 399764
rect 360068 399712 360074 399764
rect 360258 399628 360286 399848
rect 359792 399588 359918 399616
rect 359792 399576 359798 399588
rect 360194 399576 360200 399628
rect 360252 399588 360286 399628
rect 360252 399576 360258 399588
rect 359918 399508 359924 399560
rect 359976 399548 359982 399560
rect 360350 399548 360378 399848
rect 360700 399780 360706 399832
rect 360758 399780 360764 399832
rect 359976 399520 360378 399548
rect 359976 399508 359982 399520
rect 360470 399508 360476 399560
rect 360528 399548 360534 399560
rect 360718 399548 360746 399780
rect 360528 399520 360746 399548
rect 360528 399508 360534 399520
rect 358694 399452 358728 399492
rect 357308 399440 357314 399452
rect 358722 399440 358728 399452
rect 358780 399440 358786 399492
rect 359642 399440 359648 399492
rect 359700 399440 359706 399492
rect 360378 399440 360384 399492
rect 360436 399480 360442 399492
rect 360810 399480 360838 399860
rect 361068 399848 361074 399900
rect 361126 399848 361132 399900
rect 361252 399848 361258 399900
rect 361310 399848 361316 399900
rect 361344 399848 361350 399900
rect 361402 399848 361408 399900
rect 361436 399848 361442 399900
rect 361494 399888 361500 399900
rect 361494 399848 361528 399888
rect 361620 399848 361626 399900
rect 361678 399848 361684 399900
rect 361804 399848 361810 399900
rect 361862 399848 361868 399900
rect 362448 399848 362454 399900
rect 362506 399848 362512 399900
rect 362816 399848 362822 399900
rect 362874 399848 362880 399900
rect 362908 399848 362914 399900
rect 362966 399848 362972 399900
rect 363000 399848 363006 399900
rect 363058 399848 363064 399900
rect 363552 399888 363558 399900
rect 363386 399860 363558 399888
rect 361086 399628 361114 399848
rect 361086 399588 361120 399628
rect 361114 399576 361120 399588
rect 361172 399576 361178 399628
rect 361270 399560 361298 399848
rect 361362 399696 361390 399848
rect 361500 399764 361528 399848
rect 361482 399712 361488 399764
rect 361540 399712 361546 399764
rect 361638 399696 361666 399848
rect 361362 399656 361396 399696
rect 361390 399644 361396 399656
rect 361448 399644 361454 399696
rect 361574 399644 361580 399696
rect 361632 399656 361666 399696
rect 361632 399644 361638 399656
rect 361758 399576 361764 399628
rect 361816 399616 361822 399628
rect 362466 399616 362494 399848
rect 362724 399780 362730 399832
rect 362782 399780 362788 399832
rect 361816 399588 362494 399616
rect 361816 399576 361822 399588
rect 361270 399520 361304 399560
rect 361298 399508 361304 399520
rect 361356 399508 361362 399560
rect 362586 399508 362592 399560
rect 362644 399548 362650 399560
rect 362742 399548 362770 399780
rect 362834 399696 362862 399848
rect 362926 399764 362954 399848
rect 363018 399820 363046 399848
rect 363018 399792 363092 399820
rect 362926 399724 362960 399764
rect 362954 399712 362960 399724
rect 363012 399712 363018 399764
rect 362834 399656 362868 399696
rect 362862 399644 362868 399656
rect 362920 399644 362926 399696
rect 363064 399616 363092 399792
rect 363184 399780 363190 399832
rect 363242 399780 363248 399832
rect 363202 399696 363230 399780
rect 363138 399644 363144 399696
rect 363196 399656 363230 399696
rect 363196 399644 363202 399656
rect 363230 399616 363236 399628
rect 363064 399588 363236 399616
rect 363230 399576 363236 399588
rect 363288 399576 363294 399628
rect 362644 399520 362770 399548
rect 362644 399508 362650 399520
rect 360436 399452 360838 399480
rect 363386 399480 363414 399860
rect 363552 399848 363558 399860
rect 363610 399848 363616 399900
rect 363736 399848 363742 399900
rect 363794 399848 363800 399900
rect 363920 399848 363926 399900
rect 363978 399848 363984 399900
rect 364104 399848 364110 399900
rect 364162 399888 364168 399900
rect 364162 399848 364196 399888
rect 364288 399848 364294 399900
rect 364346 399848 364352 399900
rect 364380 399848 364386 399900
rect 364438 399848 364444 399900
rect 364564 399848 364570 399900
rect 364622 399848 364628 399900
rect 364840 399848 364846 399900
rect 364898 399848 364904 399900
rect 365576 399888 365582 399900
rect 364950 399860 365582 399888
rect 363460 399780 363466 399832
rect 363518 399780 363524 399832
rect 363478 399548 363506 399780
rect 363754 399764 363782 399848
rect 363828 399780 363834 399832
rect 363886 399780 363892 399832
rect 363690 399712 363696 399764
rect 363748 399724 363782 399764
rect 363748 399712 363754 399724
rect 363598 399644 363604 399696
rect 363656 399684 363662 399696
rect 363846 399684 363874 399780
rect 363656 399656 363874 399684
rect 363656 399644 363662 399656
rect 363938 399628 363966 399848
rect 364168 399764 364196 399848
rect 364150 399712 364156 399764
rect 364208 399712 364214 399764
rect 363874 399576 363880 399628
rect 363932 399588 363966 399628
rect 363932 399576 363938 399588
rect 364306 399560 364334 399848
rect 364398 399616 364426 399848
rect 364582 399684 364610 399848
rect 364858 399696 364886 399848
rect 364536 399656 364610 399684
rect 364398 399588 364472 399616
rect 364444 399560 364472 399588
rect 363598 399548 363604 399560
rect 363478 399520 363604 399548
rect 363598 399508 363604 399520
rect 363656 399508 363662 399560
rect 364306 399520 364340 399560
rect 364334 399508 364340 399520
rect 364392 399508 364398 399560
rect 364426 399508 364432 399560
rect 364484 399508 364490 399560
rect 363782 399480 363788 399492
rect 363386 399452 363788 399480
rect 360436 399440 360442 399452
rect 363782 399440 363788 399452
rect 363840 399440 363846 399492
rect 364058 399440 364064 399492
rect 364116 399480 364122 399492
rect 364536 399480 364564 399656
rect 364794 399644 364800 399696
rect 364852 399656 364886 399696
rect 364852 399644 364858 399656
rect 364610 399508 364616 399560
rect 364668 399548 364674 399560
rect 364950 399548 364978 399860
rect 365576 399848 365582 399860
rect 365634 399848 365640 399900
rect 365668 399848 365674 399900
rect 365726 399848 365732 399900
rect 365760 399848 365766 399900
rect 365818 399848 365824 399900
rect 366220 399848 366226 399900
rect 366278 399848 366284 399900
rect 366404 399848 366410 399900
rect 366462 399848 366468 399900
rect 365208 399820 365214 399832
rect 365180 399780 365214 399820
rect 365266 399780 365272 399832
rect 365392 399780 365398 399832
rect 365450 399780 365456 399832
rect 365180 399560 365208 399780
rect 365254 399644 365260 399696
rect 365312 399684 365318 399696
rect 365410 399684 365438 399780
rect 365312 399656 365438 399684
rect 365312 399644 365318 399656
rect 365686 399628 365714 399848
rect 365778 399696 365806 399848
rect 365852 399780 365858 399832
rect 365910 399780 365916 399832
rect 365944 399780 365950 399832
rect 366002 399820 366008 399832
rect 366002 399780 366036 399820
rect 365870 399752 365898 399780
rect 365870 399724 365944 399752
rect 365916 399696 365944 399724
rect 365778 399656 365812 399696
rect 365806 399644 365812 399656
rect 365864 399644 365870 399696
rect 365898 399644 365904 399696
rect 365956 399644 365962 399696
rect 365686 399588 365720 399628
rect 365714 399576 365720 399588
rect 365772 399576 365778 399628
rect 364668 399520 364978 399548
rect 364668 399508 364674 399520
rect 365162 399508 365168 399560
rect 365220 399508 365226 399560
rect 365346 399508 365352 399560
rect 365404 399548 365410 399560
rect 366008 399548 366036 399780
rect 366082 399644 366088 399696
rect 366140 399684 366146 399696
rect 366422 399684 366450 399848
rect 366140 399656 366450 399684
rect 366140 399644 366146 399656
rect 365404 399520 366036 399548
rect 365404 399508 365410 399520
rect 366174 399508 366180 399560
rect 366232 399548 366238 399560
rect 366514 399548 366542 399928
rect 366790 399928 367002 399956
rect 366790 399900 366818 399928
rect 366680 399848 366686 399900
rect 366738 399848 366744 399900
rect 366772 399848 366778 399900
rect 366830 399848 366836 399900
rect 366864 399848 366870 399900
rect 366922 399848 366928 399900
rect 366232 399520 366542 399548
rect 366232 399508 366238 399520
rect 366698 399492 366726 399848
rect 366882 399628 366910 399848
rect 366818 399576 366824 399628
rect 366876 399588 366910 399628
rect 366876 399576 366882 399588
rect 364116 399452 364564 399480
rect 364116 399440 364122 399452
rect 366634 399440 366640 399492
rect 366692 399452 366726 399492
rect 366692 399440 366698 399452
rect 359550 399412 359556 399424
rect 354876 399384 359556 399412
rect 359550 399372 359556 399384
rect 359608 399372 359614 399424
rect 365990 399372 365996 399424
rect 366048 399412 366054 399424
rect 366974 399412 367002 399928
rect 367048 399848 367054 399900
rect 367106 399848 367112 399900
rect 367416 399848 367422 399900
rect 367474 399848 367480 399900
rect 367784 399848 367790 399900
rect 367842 399848 367848 399900
rect 367968 399848 367974 399900
rect 368026 399888 368032 399900
rect 368026 399860 368290 399888
rect 368026 399848 368032 399860
rect 367066 399616 367094 399848
rect 367434 399752 367462 399848
rect 367508 399780 367514 399832
rect 367566 399780 367572 399832
rect 367388 399724 367462 399752
rect 367388 399696 367416 399724
rect 367526 399696 367554 399780
rect 367802 399696 367830 399848
rect 368060 399820 368066 399832
rect 367370 399644 367376 399696
rect 367428 399644 367434 399696
rect 367462 399644 367468 399696
rect 367520 399656 367554 399696
rect 367520 399644 367526 399656
rect 367738 399644 367744 399696
rect 367796 399656 367830 399696
rect 367894 399792 368066 399820
rect 367796 399644 367802 399656
rect 367066 399588 367140 399616
rect 367112 399560 367140 399588
rect 367186 399576 367192 399628
rect 367244 399616 367250 399628
rect 367894 399616 367922 399792
rect 368060 399780 368066 399792
rect 368118 399780 368124 399832
rect 368152 399780 368158 399832
rect 368210 399780 368216 399832
rect 368014 399644 368020 399696
rect 368072 399684 368078 399696
rect 368170 399684 368198 399780
rect 368072 399656 368198 399684
rect 368072 399644 368078 399656
rect 367244 399588 367922 399616
rect 367244 399576 367250 399588
rect 368106 399576 368112 399628
rect 368164 399616 368170 399628
rect 368262 399616 368290 399860
rect 368336 399848 368342 399900
rect 368394 399848 368400 399900
rect 368612 399848 368618 399900
rect 368670 399888 368676 399900
rect 368670 399860 368888 399888
rect 368670 399848 368676 399860
rect 368164 399588 368290 399616
rect 368164 399576 368170 399588
rect 367094 399508 367100 399560
rect 367152 399508 367158 399560
rect 368354 399492 368382 399848
rect 368428 399780 368434 399832
rect 368486 399780 368492 399832
rect 368520 399780 368526 399832
rect 368578 399780 368584 399832
rect 368290 399440 368296 399492
rect 368348 399452 368382 399492
rect 368446 399492 368474 399780
rect 368538 399560 368566 399780
rect 368860 399628 368888 399860
rect 368980 399848 368986 399900
rect 369038 399848 369044 399900
rect 369440 399848 369446 399900
rect 369498 399848 369504 399900
rect 369900 399848 369906 399900
rect 369958 399848 369964 399900
rect 369992 399848 369998 399900
rect 370050 399848 370056 399900
rect 370176 399848 370182 399900
rect 370234 399848 370240 399900
rect 368842 399576 368848 399628
rect 368900 399576 368906 399628
rect 368538 399520 368572 399560
rect 368566 399508 368572 399520
rect 368624 399508 368630 399560
rect 368446 399452 368480 399492
rect 368348 399440 368354 399452
rect 368474 399440 368480 399452
rect 368532 399440 368538 399492
rect 368658 399440 368664 399492
rect 368716 399480 368722 399492
rect 368998 399480 369026 399848
rect 369210 399712 369216 399764
rect 369268 399712 369274 399764
rect 369118 399576 369124 399628
rect 369176 399616 369182 399628
rect 369228 399616 369256 399712
rect 369176 399588 369256 399616
rect 369176 399576 369182 399588
rect 368716 399452 369026 399480
rect 368716 399440 368722 399452
rect 369458 399424 369486 399848
rect 369808 399780 369814 399832
rect 369866 399780 369872 399832
rect 369826 399684 369854 399780
rect 369688 399656 369854 399684
rect 369688 399492 369716 399656
rect 369918 399628 369946 399848
rect 369854 399576 369860 399628
rect 369912 399588 369946 399628
rect 369912 399576 369918 399588
rect 370010 399560 370038 399848
rect 370084 399780 370090 399832
rect 370142 399780 370148 399832
rect 369946 399508 369952 399560
rect 370004 399520 370038 399560
rect 370004 399508 370010 399520
rect 370102 399492 370130 399780
rect 370194 399548 370222 399848
rect 370286 399616 370314 400200
rect 374334 399900 374362 400336
rect 387518 400324 387524 400336
rect 387576 400324 387582 400376
rect 392026 400024 392032 400036
rect 383718 399996 392032 400024
rect 375760 399928 376800 399956
rect 371372 399848 371378 399900
rect 371430 399848 371436 399900
rect 371924 399848 371930 399900
rect 371982 399848 371988 399900
rect 372384 399848 372390 399900
rect 372442 399848 372448 399900
rect 372568 399848 372574 399900
rect 372626 399888 372632 399900
rect 372626 399848 372660 399888
rect 372936 399848 372942 399900
rect 372994 399848 373000 399900
rect 373488 399848 373494 399900
rect 373546 399848 373552 399900
rect 373948 399848 373954 399900
rect 374006 399848 374012 399900
rect 374040 399848 374046 399900
rect 374098 399848 374104 399900
rect 374316 399848 374322 399900
rect 374374 399848 374380 399900
rect 374592 399848 374598 399900
rect 374650 399848 374656 399900
rect 374868 399848 374874 399900
rect 374926 399848 374932 399900
rect 374960 399848 374966 399900
rect 375018 399848 375024 399900
rect 375512 399888 375518 399900
rect 375484 399848 375518 399888
rect 375570 399848 375576 399900
rect 375604 399848 375610 399900
rect 375662 399888 375668 399900
rect 375760 399888 375788 399928
rect 375880 399888 375886 399900
rect 375662 399860 375788 399888
rect 375662 399848 375668 399860
rect 375852 399848 375886 399888
rect 375938 399848 375944 399900
rect 376064 399848 376070 399900
rect 376122 399848 376128 399900
rect 376432 399888 376438 399900
rect 376174 399860 376438 399888
rect 370544 399780 370550 399832
rect 370602 399780 370608 399832
rect 370562 399696 370590 399780
rect 370562 399656 370596 399696
rect 370590 399644 370596 399656
rect 370648 399644 370654 399696
rect 370498 399616 370504 399628
rect 370286 399588 370504 399616
rect 370498 399576 370504 399588
rect 370556 399576 370562 399628
rect 371390 399616 371418 399848
rect 371942 399764 371970 399848
rect 371942 399724 371976 399764
rect 371970 399712 371976 399724
rect 372028 399712 372034 399764
rect 372402 399684 372430 399848
rect 372632 399696 372660 399848
rect 372522 399684 372528 399696
rect 372402 399656 372528 399684
rect 372522 399644 372528 399656
rect 372580 399644 372586 399696
rect 372614 399644 372620 399696
rect 372672 399644 372678 399696
rect 371390 399588 371648 399616
rect 370314 399548 370320 399560
rect 370194 399520 370320 399548
rect 370314 399508 370320 399520
rect 370372 399508 370378 399560
rect 369670 399440 369676 399492
rect 369728 399440 369734 399492
rect 370102 399452 370136 399492
rect 370130 399440 370136 399452
rect 370188 399440 370194 399492
rect 366048 399384 367002 399412
rect 366048 399372 366054 399384
rect 369394 399372 369400 399424
rect 369452 399384 369486 399424
rect 369452 399372 369458 399384
rect 348752 399316 350212 399344
rect 348752 399304 348758 399316
rect 350902 399304 350908 399356
rect 350960 399344 350966 399356
rect 351178 399344 351184 399356
rect 350960 399316 351184 399344
rect 350960 399304 350966 399316
rect 351178 399304 351184 399316
rect 351236 399304 351242 399356
rect 351270 399304 351276 399356
rect 351328 399344 351334 399356
rect 353202 399344 353208 399356
rect 351328 399316 353208 399344
rect 351328 399304 351334 399316
rect 353202 399304 353208 399316
rect 353260 399344 353266 399356
rect 360286 399344 360292 399356
rect 353260 399316 360292 399344
rect 353260 399304 353266 399316
rect 360286 399304 360292 399316
rect 360344 399304 360350 399356
rect 363046 399304 363052 399356
rect 363104 399344 363110 399356
rect 363414 399344 363420 399356
rect 363104 399316 363420 399344
rect 363104 399304 363110 399316
rect 363414 399304 363420 399316
rect 363472 399304 363478 399356
rect 365686 399316 366910 399344
rect 361022 399276 361028 399288
rect 349126 399248 361028 399276
rect 349126 399208 349154 399248
rect 361022 399236 361028 399248
rect 361080 399236 361086 399288
rect 347056 399180 349154 399208
rect 351178 399168 351184 399220
rect 351236 399208 351242 399220
rect 359550 399208 359556 399220
rect 351236 399180 359556 399208
rect 351236 399168 351242 399180
rect 359550 399168 359556 399180
rect 359608 399168 359614 399220
rect 365686 399208 365714 399316
rect 364260 399180 365714 399208
rect 366882 399208 366910 399316
rect 370682 399304 370688 399356
rect 370740 399344 370746 399356
rect 370958 399344 370964 399356
rect 370740 399316 370964 399344
rect 370740 399304 370746 399316
rect 370958 399304 370964 399316
rect 371016 399304 371022 399356
rect 371510 399304 371516 399356
rect 371568 399344 371574 399356
rect 371620 399344 371648 399588
rect 372798 399576 372804 399628
rect 372856 399616 372862 399628
rect 372954 399616 372982 399848
rect 373506 399616 373534 399848
rect 372856 399588 372982 399616
rect 373276 399588 373534 399616
rect 372856 399576 372862 399588
rect 373276 399560 373304 399588
rect 373258 399508 373264 399560
rect 373316 399508 373322 399560
rect 373966 399492 373994 399848
rect 374058 399548 374086 399848
rect 374610 399560 374638 399848
rect 374362 399548 374368 399560
rect 374058 399520 374368 399548
rect 374362 399508 374368 399520
rect 374420 399508 374426 399560
rect 374610 399520 374644 399560
rect 374638 399508 374644 399520
rect 374696 399508 374702 399560
rect 374730 399508 374736 399560
rect 374788 399548 374794 399560
rect 374886 399548 374914 399848
rect 374978 399628 375006 399848
rect 375484 399764 375512 399848
rect 375466 399712 375472 399764
rect 375524 399712 375530 399764
rect 374978 399588 375012 399628
rect 375006 399576 375012 399588
rect 375064 399576 375070 399628
rect 374788 399520 374914 399548
rect 375852 399548 375880 399848
rect 375972 399820 375978 399832
rect 375944 399780 375978 399820
rect 376030 399780 376036 399832
rect 375944 399696 375972 399780
rect 375926 399644 375932 399696
rect 375984 399644 375990 399696
rect 376082 399628 376110 399848
rect 376018 399576 376024 399628
rect 376076 399588 376110 399628
rect 376076 399576 376082 399588
rect 375926 399548 375932 399560
rect 375852 399520 375932 399548
rect 374788 399508 374794 399520
rect 375926 399508 375932 399520
rect 375984 399508 375990 399560
rect 373534 399440 373540 399492
rect 373592 399480 373598 399492
rect 373718 399480 373724 399492
rect 373592 399452 373724 399480
rect 373592 399440 373598 399452
rect 373718 399440 373724 399452
rect 373776 399440 373782 399492
rect 373966 399452 374000 399492
rect 373994 399440 374000 399452
rect 374052 399440 374058 399492
rect 375650 399372 375656 399424
rect 375708 399412 375714 399424
rect 376174 399412 376202 399860
rect 376432 399848 376438 399860
rect 376490 399848 376496 399900
rect 376616 399848 376622 399900
rect 376674 399848 376680 399900
rect 376478 399712 376484 399764
rect 376536 399752 376542 399764
rect 376634 399752 376662 399848
rect 376536 399724 376662 399752
rect 376536 399712 376542 399724
rect 376772 399480 376800 399928
rect 381418 399928 381814 399956
rect 381418 399900 381446 399928
rect 376892 399848 376898 399900
rect 376950 399888 376956 399900
rect 376950 399848 376984 399888
rect 377076 399848 377082 399900
rect 377134 399848 377140 399900
rect 377260 399848 377266 399900
rect 377318 399848 377324 399900
rect 377628 399848 377634 399900
rect 377686 399848 377692 399900
rect 377812 399848 377818 399900
rect 377870 399848 377876 399900
rect 377904 399848 377910 399900
rect 377962 399848 377968 399900
rect 378088 399888 378094 399900
rect 378014 399860 378094 399888
rect 376956 399764 376984 399848
rect 376938 399712 376944 399764
rect 376996 399712 377002 399764
rect 376846 399508 376852 399560
rect 376904 399548 376910 399560
rect 377094 399548 377122 399848
rect 377278 399616 377306 399848
rect 377646 399696 377674 399848
rect 377830 399696 377858 399848
rect 377646 399656 377680 399696
rect 377674 399644 377680 399656
rect 377732 399644 377738 399696
rect 377766 399644 377772 399696
rect 377824 399656 377858 399696
rect 377824 399644 377830 399656
rect 377922 399628 377950 399848
rect 377278 399588 377536 399616
rect 377508 399560 377536 399588
rect 377858 399576 377864 399628
rect 377916 399588 377950 399628
rect 377916 399576 377922 399588
rect 378014 399560 378042 399860
rect 378088 399848 378094 399860
rect 378146 399848 378152 399900
rect 378272 399848 378278 399900
rect 378330 399848 378336 399900
rect 378640 399848 378646 399900
rect 378698 399848 378704 399900
rect 378916 399848 378922 399900
rect 378974 399848 378980 399900
rect 379008 399848 379014 399900
rect 379066 399848 379072 399900
rect 379100 399848 379106 399900
rect 379158 399848 379164 399900
rect 379376 399848 379382 399900
rect 379434 399848 379440 399900
rect 379836 399848 379842 399900
rect 379894 399848 379900 399900
rect 380296 399848 380302 399900
rect 380354 399848 380360 399900
rect 380480 399848 380486 399900
rect 380538 399888 380544 399900
rect 380538 399848 380572 399888
rect 380756 399848 380762 399900
rect 380814 399848 380820 399900
rect 380940 399848 380946 399900
rect 380998 399848 381004 399900
rect 381308 399848 381314 399900
rect 381366 399848 381372 399900
rect 381400 399848 381406 399900
rect 381458 399848 381464 399900
rect 381492 399848 381498 399900
rect 381550 399848 381556 399900
rect 381676 399848 381682 399900
rect 381734 399848 381740 399900
rect 376904 399520 377122 399548
rect 376904 399508 376910 399520
rect 377490 399508 377496 399560
rect 377548 399508 377554 399560
rect 377950 399508 377956 399560
rect 378008 399520 378042 399560
rect 378008 399508 378014 399520
rect 377122 399480 377128 399492
rect 376772 399452 377128 399480
rect 377122 399440 377128 399452
rect 377180 399440 377186 399492
rect 378290 399480 378318 399848
rect 378658 399764 378686 399848
rect 378934 399820 378962 399848
rect 378796 399792 378962 399820
rect 378658 399724 378692 399764
rect 378686 399712 378692 399724
rect 378744 399712 378750 399764
rect 378410 399576 378416 399628
rect 378468 399616 378474 399628
rect 378796 399616 378824 399792
rect 379026 399752 379054 399848
rect 378468 399588 378824 399616
rect 378980 399724 379054 399752
rect 378468 399576 378474 399588
rect 378980 399548 379008 399724
rect 379118 399696 379146 399848
rect 379394 399764 379422 399848
rect 379560 399780 379566 399832
rect 379618 399780 379624 399832
rect 379394 399724 379428 399764
rect 379422 399712 379428 399724
rect 379480 399712 379486 399764
rect 379054 399644 379060 399696
rect 379112 399656 379146 399696
rect 379112 399644 379118 399656
rect 379330 399548 379336 399560
rect 378980 399520 379336 399548
rect 379330 399508 379336 399520
rect 379388 399508 379394 399560
rect 378502 399480 378508 399492
rect 378290 399452 378508 399480
rect 378502 399440 378508 399452
rect 378560 399440 378566 399492
rect 379578 399480 379606 399780
rect 379854 399764 379882 399848
rect 379790 399712 379796 399764
rect 379848 399724 379882 399764
rect 379848 399712 379854 399724
rect 380314 399560 380342 399848
rect 380544 399696 380572 399848
rect 380774 399696 380802 399848
rect 380958 399752 380986 399848
rect 380912 399724 380986 399752
rect 380526 399644 380532 399696
rect 380584 399644 380590 399696
rect 380774 399656 380808 399696
rect 380802 399644 380808 399656
rect 380860 399644 380866 399696
rect 380250 399508 380256 399560
rect 380308 399520 380342 399560
rect 380912 399548 380940 399724
rect 381326 399684 381354 399848
rect 381510 399820 381538 399848
rect 381464 399792 381538 399820
rect 381464 399696 381492 399792
rect 381096 399656 381354 399684
rect 381096 399628 381124 399656
rect 381446 399644 381452 399696
rect 381504 399644 381510 399696
rect 381538 399644 381544 399696
rect 381596 399684 381602 399696
rect 381694 399684 381722 399848
rect 381596 399656 381722 399684
rect 381786 399696 381814 399928
rect 383718 399900 383746 399996
rect 392026 399984 392032 399996
rect 392084 399984 392090 400036
rect 390554 399956 390560 399968
rect 386386 399928 390560 399956
rect 386386 399900 386414 399928
rect 390554 399916 390560 399928
rect 390612 399916 390618 399968
rect 381952 399848 381958 399900
rect 382010 399848 382016 399900
rect 382136 399848 382142 399900
rect 382194 399848 382200 399900
rect 382412 399848 382418 399900
rect 382470 399848 382476 399900
rect 383056 399848 383062 399900
rect 383114 399888 383120 399900
rect 383114 399848 383148 399888
rect 383240 399848 383246 399900
rect 383298 399848 383304 399900
rect 383700 399848 383706 399900
rect 383758 399848 383764 399900
rect 383884 399848 383890 399900
rect 383942 399848 383948 399900
rect 384252 399848 384258 399900
rect 384310 399848 384316 399900
rect 384620 399848 384626 399900
rect 384678 399848 384684 399900
rect 384804 399848 384810 399900
rect 384862 399848 384868 399900
rect 385448 399848 385454 399900
rect 385506 399848 385512 399900
rect 385724 399888 385730 399900
rect 385558 399860 385730 399888
rect 381786 399656 381820 399696
rect 381596 399644 381602 399656
rect 381814 399644 381820 399656
rect 381872 399644 381878 399696
rect 381078 399576 381084 399628
rect 381136 399576 381142 399628
rect 381262 399576 381268 399628
rect 381320 399616 381326 399628
rect 381970 399616 381998 399848
rect 382154 399696 382182 399848
rect 382154 399656 382188 399696
rect 382182 399644 382188 399656
rect 382240 399644 382246 399696
rect 381320 399588 381998 399616
rect 381320 399576 381326 399588
rect 381170 399548 381176 399560
rect 380912 399520 381176 399548
rect 380308 399508 380314 399520
rect 381170 399508 381176 399520
rect 381228 399508 381234 399560
rect 379882 399480 379888 399492
rect 379578 399452 379888 399480
rect 379882 399440 379888 399452
rect 379940 399440 379946 399492
rect 382430 399480 382458 399848
rect 383120 399764 383148 399848
rect 383102 399712 383108 399764
rect 383160 399712 383166 399764
rect 382550 399508 382556 399560
rect 382608 399548 382614 399560
rect 383258 399548 383286 399848
rect 383902 399696 383930 399848
rect 383902 399656 383936 399696
rect 383930 399644 383936 399656
rect 383988 399644 383994 399696
rect 384114 399644 384120 399696
rect 384172 399684 384178 399696
rect 384270 399684 384298 399848
rect 384638 399696 384666 399848
rect 384822 399752 384850 399848
rect 384822 399724 384988 399752
rect 384960 399696 384988 399724
rect 384172 399656 384298 399684
rect 384172 399644 384178 399656
rect 384574 399644 384580 399696
rect 384632 399656 384666 399696
rect 384632 399644 384638 399656
rect 384942 399644 384948 399696
rect 385000 399644 385006 399696
rect 382608 399520 383286 399548
rect 382608 399508 382614 399520
rect 382430 399452 383608 399480
rect 383580 399424 383608 399452
rect 375708 399384 376202 399412
rect 375708 399372 375714 399384
rect 381170 399372 381176 399424
rect 381228 399412 381234 399424
rect 381446 399412 381452 399424
rect 381228 399384 381452 399412
rect 381228 399372 381234 399384
rect 381446 399372 381452 399384
rect 381504 399372 381510 399424
rect 381630 399372 381636 399424
rect 381688 399412 381694 399424
rect 382090 399412 382096 399424
rect 381688 399384 382096 399412
rect 381688 399372 381694 399384
rect 382090 399372 382096 399384
rect 382148 399372 382154 399424
rect 382274 399372 382280 399424
rect 382332 399412 382338 399424
rect 382550 399412 382556 399424
rect 382332 399384 382556 399412
rect 382332 399372 382338 399384
rect 382550 399372 382556 399384
rect 382608 399372 382614 399424
rect 383562 399372 383568 399424
rect 383620 399372 383626 399424
rect 385466 399412 385494 399848
rect 385558 399560 385586 399860
rect 385724 399848 385730 399860
rect 385782 399848 385788 399900
rect 385908 399848 385914 399900
rect 385966 399848 385972 399900
rect 386000 399848 386006 399900
rect 386058 399848 386064 399900
rect 386184 399848 386190 399900
rect 386242 399848 386248 399900
rect 386368 399848 386374 399900
rect 386426 399848 386432 399900
rect 386920 399848 386926 399900
rect 386978 399848 386984 399900
rect 387012 399848 387018 399900
rect 387070 399848 387076 399900
rect 385926 399696 385954 399848
rect 385862 399644 385868 399696
rect 385920 399656 385954 399696
rect 386018 399696 386046 399848
rect 386018 399656 386052 399696
rect 385920 399644 385926 399656
rect 386046 399644 386052 399656
rect 386104 399644 386110 399696
rect 386202 399684 386230 399848
rect 386460 399780 386466 399832
rect 386518 399780 386524 399832
rect 386322 399712 386328 399764
rect 386380 399752 386386 399764
rect 386478 399752 386506 399780
rect 386938 399752 386966 399848
rect 386380 399724 386506 399752
rect 386892 399724 386966 399752
rect 386380 399712 386386 399724
rect 386782 399684 386788 399696
rect 386202 399656 386788 399684
rect 386782 399644 386788 399656
rect 386840 399644 386846 399696
rect 386414 399576 386420 399628
rect 386472 399616 386478 399628
rect 386892 399616 386920 399724
rect 387030 399696 387058 399848
rect 386966 399644 386972 399696
rect 387024 399656 387058 399696
rect 387024 399644 387030 399656
rect 386472 399588 386920 399616
rect 386472 399576 386478 399588
rect 385558 399520 385592 399560
rect 385586 399508 385592 399520
rect 385644 399508 385650 399560
rect 385678 399508 385684 399560
rect 385736 399508 385742 399560
rect 385696 399480 385724 399508
rect 387978 399480 387984 399492
rect 385696 399452 387984 399480
rect 387978 399440 387984 399452
rect 388036 399440 388042 399492
rect 580258 399480 580264 399492
rect 396046 399452 580264 399480
rect 385678 399412 385684 399424
rect 385466 399384 385684 399412
rect 385678 399372 385684 399384
rect 385736 399372 385742 399424
rect 371568 399316 371648 399344
rect 371568 399304 371574 399316
rect 371694 399304 371700 399356
rect 371752 399304 371758 399356
rect 370222 399236 370228 399288
rect 370280 399276 370286 399288
rect 371712 399276 371740 399304
rect 370280 399248 371740 399276
rect 370280 399236 370286 399248
rect 376294 399236 376300 399288
rect 376352 399276 376358 399288
rect 380158 399276 380164 399288
rect 376352 399248 380164 399276
rect 376352 399236 376358 399248
rect 380158 399236 380164 399248
rect 380216 399236 380222 399288
rect 366882 399180 371234 399208
rect 364260 399152 364288 399180
rect 338942 399100 338948 399152
rect 339000 399140 339006 399152
rect 362954 399140 362960 399152
rect 339000 399112 362960 399140
rect 339000 399100 339006 399112
rect 362954 399100 362960 399112
rect 363012 399100 363018 399152
rect 364242 399100 364248 399152
rect 364300 399100 364306 399152
rect 371206 399140 371234 399180
rect 372706 399168 372712 399220
rect 372764 399208 372770 399220
rect 373902 399208 373908 399220
rect 372764 399180 373908 399208
rect 372764 399168 372770 399180
rect 373902 399168 373908 399180
rect 373960 399168 373966 399220
rect 380250 399208 380256 399220
rect 375806 399180 380256 399208
rect 375806 399140 375834 399180
rect 380250 399168 380256 399180
rect 380308 399168 380314 399220
rect 384482 399168 384488 399220
rect 384540 399208 384546 399220
rect 384942 399208 384948 399220
rect 384540 399180 384948 399208
rect 384540 399168 384546 399180
rect 384942 399168 384948 399180
rect 385000 399168 385006 399220
rect 385770 399168 385776 399220
rect 385828 399208 385834 399220
rect 396046 399208 396074 399452
rect 580258 399440 580264 399452
rect 580316 399440 580322 399492
rect 385828 399180 396074 399208
rect 385828 399168 385834 399180
rect 371206 399112 375834 399140
rect 379606 399100 379612 399152
rect 379664 399140 379670 399152
rect 380526 399140 380532 399152
rect 379664 399112 380532 399140
rect 379664 399100 379670 399112
rect 380526 399100 380532 399112
rect 380584 399100 380590 399152
rect 382090 399100 382096 399152
rect 382148 399140 382154 399152
rect 385862 399140 385868 399152
rect 382148 399112 385868 399140
rect 382148 399100 382154 399112
rect 385862 399100 385868 399112
rect 385920 399100 385926 399152
rect 281350 399032 281356 399084
rect 281408 399072 281414 399084
rect 358170 399072 358176 399084
rect 281408 399044 358176 399072
rect 281408 399032 281414 399044
rect 358170 399032 358176 399044
rect 358228 399032 358234 399084
rect 372246 399072 372252 399084
rect 363064 399044 372252 399072
rect 276842 398964 276848 399016
rect 276900 399004 276906 399016
rect 349154 399004 349160 399016
rect 276900 398976 349160 399004
rect 276900 398964 276906 398976
rect 349154 398964 349160 398976
rect 349212 398964 349218 399016
rect 359734 399004 359740 399016
rect 353266 398976 359740 399004
rect 276750 398896 276756 398948
rect 276808 398936 276814 398948
rect 346210 398936 346216 398948
rect 276808 398908 346216 398936
rect 276808 398896 276814 398908
rect 346210 398896 346216 398908
rect 346268 398896 346274 398948
rect 346670 398896 346676 398948
rect 346728 398936 346734 398948
rect 353266 398936 353294 398976
rect 359734 398964 359740 398976
rect 359792 398964 359798 399016
rect 360286 398964 360292 399016
rect 360344 399004 360350 399016
rect 363064 399004 363092 399044
rect 372246 399032 372252 399044
rect 372304 399032 372310 399084
rect 373902 399032 373908 399084
rect 373960 399072 373966 399084
rect 374270 399072 374276 399084
rect 373960 399044 374276 399072
rect 373960 399032 373966 399044
rect 374270 399032 374276 399044
rect 374328 399032 374334 399084
rect 381906 399032 381912 399084
rect 381964 399072 381970 399084
rect 393314 399072 393320 399084
rect 381964 399044 393320 399072
rect 381964 399032 381970 399044
rect 393314 399032 393320 399044
rect 393372 399032 393378 399084
rect 380618 399004 380624 399016
rect 360344 398976 363092 399004
rect 364996 398976 380624 399004
rect 360344 398964 360350 398976
rect 346728 398908 353294 398936
rect 346728 398896 346734 398908
rect 357802 398896 357808 398948
rect 357860 398936 357866 398948
rect 358998 398936 359004 398948
rect 357860 398908 359004 398936
rect 357860 398896 357866 398908
rect 358998 398896 359004 398908
rect 359056 398896 359062 398948
rect 359550 398896 359556 398948
rect 359608 398936 359614 398948
rect 364242 398936 364248 398948
rect 359608 398908 364248 398936
rect 359608 398896 359614 398908
rect 364242 398896 364248 398908
rect 364300 398896 364306 398948
rect 337654 398828 337660 398880
rect 337712 398868 337718 398880
rect 364996 398868 365024 398976
rect 380618 398964 380624 398976
rect 380676 398964 380682 399016
rect 385862 398964 385868 399016
rect 385920 399004 385926 399016
rect 393498 399004 393504 399016
rect 385920 398976 393504 399004
rect 385920 398964 385926 398976
rect 393498 398964 393504 398976
rect 393556 398964 393562 399016
rect 372246 398896 372252 398948
rect 372304 398936 372310 398948
rect 376294 398936 376300 398948
rect 372304 398908 376300 398936
rect 372304 398896 372310 398908
rect 376294 398896 376300 398908
rect 376352 398896 376358 398948
rect 379606 398896 379612 398948
rect 379664 398936 379670 398948
rect 380802 398936 380808 398948
rect 379664 398908 380808 398936
rect 379664 398896 379670 398908
rect 380802 398896 380808 398908
rect 380860 398896 380866 398948
rect 387518 398896 387524 398948
rect 387576 398936 387582 398948
rect 394970 398936 394976 398948
rect 387576 398908 394976 398936
rect 387576 398896 387582 398908
rect 394970 398896 394976 398908
rect 395028 398896 395034 398948
rect 337712 398840 365024 398868
rect 337712 398828 337718 398840
rect 368934 398828 368940 398880
rect 368992 398868 368998 398880
rect 369302 398868 369308 398880
rect 368992 398840 369308 398868
rect 368992 398828 368998 398840
rect 369302 398828 369308 398840
rect 369360 398828 369366 398880
rect 373810 398828 373816 398880
rect 373868 398868 373874 398880
rect 373868 398840 375236 398868
rect 373868 398828 373874 398840
rect 327718 398760 327724 398812
rect 327776 398800 327782 398812
rect 344646 398800 344652 398812
rect 327776 398772 344652 398800
rect 327776 398760 327782 398772
rect 344646 398760 344652 398772
rect 344704 398760 344710 398812
rect 346394 398800 346400 398812
rect 344756 398772 346400 398800
rect 343450 398692 343456 398744
rect 343508 398732 343514 398744
rect 344756 398732 344784 398772
rect 346394 398760 346400 398772
rect 346452 398760 346458 398812
rect 360470 398800 360476 398812
rect 346734 398772 349752 398800
rect 343508 398704 344784 398732
rect 343508 398692 343514 398704
rect 345106 398692 345112 398744
rect 345164 398732 345170 398744
rect 346734 398732 346762 398772
rect 345164 398704 346762 398732
rect 349724 398732 349752 398772
rect 357176 398772 360476 398800
rect 357176 398732 357204 398772
rect 360470 398760 360476 398772
rect 360528 398760 360534 398812
rect 360838 398760 360844 398812
rect 360896 398800 360902 398812
rect 366542 398800 366548 398812
rect 360896 398772 366548 398800
rect 360896 398760 360902 398772
rect 366542 398760 366548 398772
rect 366600 398760 366606 398812
rect 367020 398772 375144 398800
rect 360654 398732 360660 398744
rect 349724 398704 357204 398732
rect 357268 398704 360660 398732
rect 345164 398692 345170 398704
rect 300394 398624 300400 398676
rect 300452 398664 300458 398676
rect 344278 398664 344284 398676
rect 300452 398636 344284 398664
rect 300452 398624 300458 398636
rect 344278 398624 344284 398636
rect 344336 398624 344342 398676
rect 344462 398624 344468 398676
rect 344520 398664 344526 398676
rect 345474 398664 345480 398676
rect 344520 398636 345480 398664
rect 344520 398624 344526 398636
rect 345474 398624 345480 398636
rect 345532 398624 345538 398676
rect 346210 398624 346216 398676
rect 346268 398664 346274 398676
rect 350442 398664 350448 398676
rect 346268 398636 350448 398664
rect 346268 398624 346274 398636
rect 350442 398624 350448 398636
rect 350500 398624 350506 398676
rect 351822 398624 351828 398676
rect 351880 398664 351886 398676
rect 357268 398664 357296 398704
rect 360654 398692 360660 398704
rect 360712 398692 360718 398744
rect 361482 398692 361488 398744
rect 361540 398732 361546 398744
rect 367020 398732 367048 398772
rect 361540 398704 367048 398732
rect 361540 398692 361546 398704
rect 351880 398636 357296 398664
rect 351880 398624 351886 398636
rect 366542 398624 366548 398676
rect 366600 398664 366606 398676
rect 368934 398664 368940 398676
rect 366600 398636 368940 398664
rect 366600 398624 366606 398636
rect 368934 398624 368940 398636
rect 368992 398624 368998 398676
rect 329190 398556 329196 398608
rect 329248 398596 329254 398608
rect 362402 398596 362408 398608
rect 329248 398568 362408 398596
rect 329248 398556 329254 398568
rect 362402 398556 362408 398568
rect 362460 398556 362466 398608
rect 362862 398556 362868 398608
rect 362920 398596 362926 398608
rect 373902 398596 373908 398608
rect 362920 398568 373908 398596
rect 362920 398556 362926 398568
rect 373902 398556 373908 398568
rect 373960 398556 373966 398608
rect 309962 398488 309968 398540
rect 310020 398528 310026 398540
rect 344462 398528 344468 398540
rect 310020 398500 344468 398528
rect 310020 398488 310026 398500
rect 344462 398488 344468 398500
rect 344520 398488 344526 398540
rect 354766 398528 354772 398540
rect 345308 398500 354772 398528
rect 305086 398420 305092 398472
rect 305144 398460 305150 398472
rect 343634 398460 343640 398472
rect 305144 398432 343640 398460
rect 305144 398420 305150 398432
rect 343634 398420 343640 398432
rect 343692 398420 343698 398472
rect 304994 398352 305000 398404
rect 305052 398392 305058 398404
rect 343818 398392 343824 398404
rect 305052 398364 343824 398392
rect 305052 398352 305058 398364
rect 343818 398352 343824 398364
rect 343876 398352 343882 398404
rect 345308 398392 345336 398500
rect 354766 398488 354772 398500
rect 354824 398488 354830 398540
rect 358170 398488 358176 398540
rect 358228 398528 358234 398540
rect 362310 398528 362316 398540
rect 358228 398500 362316 398528
rect 358228 398488 358234 398500
rect 362310 398488 362316 398500
rect 362368 398488 362374 398540
rect 369762 398488 369768 398540
rect 369820 398528 369826 398540
rect 373442 398528 373448 398540
rect 369820 398500 373448 398528
rect 369820 398488 369826 398500
rect 373442 398488 373448 398500
rect 373500 398488 373506 398540
rect 375116 398528 375144 398772
rect 375208 398596 375236 398840
rect 379882 398828 379888 398880
rect 379940 398868 379946 398880
rect 393406 398868 393412 398880
rect 379940 398840 393412 398868
rect 379940 398828 379946 398840
rect 393406 398828 393412 398840
rect 393464 398828 393470 398880
rect 379790 398760 379796 398812
rect 379848 398800 379854 398812
rect 379974 398800 379980 398812
rect 379848 398772 379980 398800
rect 379848 398760 379854 398772
rect 379974 398760 379980 398772
rect 380032 398760 380038 398812
rect 380158 398760 380164 398812
rect 380216 398800 380222 398812
rect 385770 398800 385776 398812
rect 380216 398772 385776 398800
rect 380216 398760 380222 398772
rect 385770 398760 385776 398772
rect 385828 398760 385834 398812
rect 377950 398692 377956 398744
rect 378008 398732 378014 398744
rect 378008 398704 380894 398732
rect 378008 398692 378014 398704
rect 379974 398664 379980 398676
rect 377968 398636 379980 398664
rect 377968 398596 377996 398636
rect 379974 398624 379980 398636
rect 380032 398624 380038 398676
rect 375208 398568 377996 398596
rect 380866 398596 380894 398704
rect 382642 398692 382648 398744
rect 382700 398732 382706 398744
rect 389266 398732 389272 398744
rect 382700 398704 389272 398732
rect 382700 398692 382706 398704
rect 389266 398692 389272 398704
rect 389324 398692 389330 398744
rect 382826 398624 382832 398676
rect 382884 398664 382890 398676
rect 383010 398664 383016 398676
rect 382884 398636 383016 398664
rect 382884 398624 382890 398636
rect 383010 398624 383016 398636
rect 383068 398624 383074 398676
rect 389174 398596 389180 398608
rect 380866 398568 389180 398596
rect 389174 398556 389180 398568
rect 389232 398556 389238 398608
rect 380894 398528 380900 398540
rect 375116 398500 380900 398528
rect 380894 398488 380900 398500
rect 380952 398488 380958 398540
rect 381446 398488 381452 398540
rect 381504 398528 381510 398540
rect 392210 398528 392216 398540
rect 381504 398500 392216 398528
rect 381504 398488 381510 398500
rect 392210 398488 392216 398500
rect 392268 398488 392274 398540
rect 348326 398420 348332 398472
rect 348384 398460 348390 398472
rect 357342 398460 357348 398472
rect 348384 398432 357348 398460
rect 348384 398420 348390 398432
rect 357342 398420 357348 398432
rect 357400 398420 357406 398472
rect 377582 398420 377588 398472
rect 377640 398460 377646 398472
rect 377950 398460 377956 398472
rect 377640 398432 377956 398460
rect 377640 398420 377646 398432
rect 377950 398420 377956 398432
rect 378008 398420 378014 398472
rect 382366 398420 382372 398472
rect 382424 398460 382430 398472
rect 389634 398460 389640 398472
rect 382424 398432 389640 398460
rect 382424 398420 382430 398432
rect 389634 398420 389640 398432
rect 389692 398420 389698 398472
rect 344204 398364 345336 398392
rect 342070 398284 342076 398336
rect 342128 398324 342134 398336
rect 344204 398324 344232 398364
rect 349154 398352 349160 398404
rect 349212 398392 349218 398404
rect 352190 398392 352196 398404
rect 349212 398364 352196 398392
rect 349212 398352 349218 398364
rect 352190 398352 352196 398364
rect 352248 398352 352254 398404
rect 357066 398352 357072 398404
rect 357124 398392 357130 398404
rect 357618 398392 357624 398404
rect 357124 398364 357624 398392
rect 357124 398352 357130 398364
rect 357618 398352 357624 398364
rect 357676 398352 357682 398404
rect 357986 398352 357992 398404
rect 358044 398392 358050 398404
rect 371142 398392 371148 398404
rect 358044 398364 371148 398392
rect 358044 398352 358050 398364
rect 371142 398352 371148 398364
rect 371200 398352 371206 398404
rect 373258 398352 373264 398404
rect 373316 398392 373322 398404
rect 382826 398392 382832 398404
rect 373316 398364 382832 398392
rect 373316 398352 373322 398364
rect 382826 398352 382832 398364
rect 382884 398352 382890 398404
rect 383654 398352 383660 398404
rect 383712 398392 383718 398404
rect 388162 398392 388168 398404
rect 383712 398364 388168 398392
rect 383712 398352 383718 398364
rect 388162 398352 388168 398364
rect 388220 398352 388226 398404
rect 342128 398296 344232 398324
rect 342128 398284 342134 398296
rect 344278 398284 344284 398336
rect 344336 398324 344342 398336
rect 352006 398324 352012 398336
rect 344336 398296 352012 398324
rect 344336 398284 344342 398296
rect 352006 398284 352012 398296
rect 352064 398284 352070 398336
rect 360654 398284 360660 398336
rect 360712 398324 360718 398336
rect 374546 398324 374552 398336
rect 360712 398296 374552 398324
rect 360712 398284 360718 398296
rect 374546 398284 374552 398296
rect 374604 398284 374610 398336
rect 374656 398296 379514 398324
rect 282914 398216 282920 398268
rect 282972 398256 282978 398268
rect 327534 398256 327540 398268
rect 282972 398228 327540 398256
rect 282972 398216 282978 398228
rect 327534 398216 327540 398228
rect 327592 398216 327598 398268
rect 344554 398216 344560 398268
rect 344612 398256 344618 398268
rect 351178 398256 351184 398268
rect 344612 398228 351184 398256
rect 344612 398216 344618 398228
rect 351178 398216 351184 398228
rect 351236 398216 351242 398268
rect 352282 398216 352288 398268
rect 352340 398256 352346 398268
rect 352650 398256 352656 398268
rect 352340 398228 352656 398256
rect 352340 398216 352346 398228
rect 352650 398216 352656 398228
rect 352708 398216 352714 398268
rect 353386 398216 353392 398268
rect 353444 398256 353450 398268
rect 355318 398256 355324 398268
rect 353444 398228 355324 398256
rect 353444 398216 353450 398228
rect 355318 398216 355324 398228
rect 355376 398216 355382 398268
rect 357618 398216 357624 398268
rect 357676 398256 357682 398268
rect 358814 398256 358820 398268
rect 357676 398228 358820 398256
rect 357676 398216 357682 398228
rect 358814 398216 358820 398228
rect 358872 398216 358878 398268
rect 362218 398216 362224 398268
rect 362276 398256 362282 398268
rect 369670 398256 369676 398268
rect 362276 398228 369676 398256
rect 362276 398216 362282 398228
rect 369670 398216 369676 398228
rect 369728 398216 369734 398268
rect 372246 398216 372252 398268
rect 372304 398256 372310 398268
rect 374656 398256 374684 398296
rect 372304 398228 374684 398256
rect 372304 398216 372310 398228
rect 376754 398216 376760 398268
rect 376812 398256 376818 398268
rect 377582 398256 377588 398268
rect 376812 398228 377588 398256
rect 376812 398216 376818 398228
rect 377582 398216 377588 398228
rect 377640 398216 377646 398268
rect 379486 398256 379514 398296
rect 383654 398256 383660 398268
rect 379486 398228 383660 398256
rect 383654 398216 383660 398228
rect 383712 398216 383718 398268
rect 276934 398148 276940 398200
rect 276992 398188 276998 398200
rect 335630 398188 335636 398200
rect 276992 398160 335636 398188
rect 276992 398148 276998 398160
rect 335630 398148 335636 398160
rect 335688 398148 335694 398200
rect 342530 398148 342536 398200
rect 342588 398188 342594 398200
rect 342714 398188 342720 398200
rect 342588 398160 342720 398188
rect 342588 398148 342594 398160
rect 342714 398148 342720 398160
rect 342772 398148 342778 398200
rect 344094 398148 344100 398200
rect 344152 398188 344158 398200
rect 355410 398188 355416 398200
rect 344152 398160 355416 398188
rect 344152 398148 344158 398160
rect 355410 398148 355416 398160
rect 355468 398148 355474 398200
rect 377122 398148 377128 398200
rect 377180 398188 377186 398200
rect 387794 398188 387800 398200
rect 377180 398160 387800 398188
rect 377180 398148 377186 398160
rect 387794 398148 387800 398160
rect 387852 398148 387858 398200
rect 389358 398188 389364 398200
rect 389146 398160 389364 398188
rect 341886 398080 341892 398132
rect 341944 398120 341950 398132
rect 345106 398120 345112 398132
rect 341944 398092 345112 398120
rect 341944 398080 341950 398092
rect 345106 398080 345112 398092
rect 345164 398080 345170 398132
rect 346394 398080 346400 398132
rect 346452 398120 346458 398132
rect 349154 398120 349160 398132
rect 346452 398092 349160 398120
rect 346452 398080 346458 398092
rect 349154 398080 349160 398092
rect 349212 398080 349218 398132
rect 358814 398080 358820 398132
rect 358872 398120 358878 398132
rect 376754 398120 376760 398132
rect 358872 398092 376760 398120
rect 358872 398080 358878 398092
rect 376754 398080 376760 398092
rect 376812 398080 376818 398132
rect 347038 398012 347044 398064
rect 347096 398052 347102 398064
rect 347682 398052 347688 398064
rect 347096 398024 347688 398052
rect 347096 398012 347102 398024
rect 347682 398012 347688 398024
rect 347740 398012 347746 398064
rect 352006 398012 352012 398064
rect 352064 398052 352070 398064
rect 356238 398052 356244 398064
rect 352064 398024 356244 398052
rect 352064 398012 352070 398024
rect 356238 398012 356244 398024
rect 356296 398012 356302 398064
rect 357158 398012 357164 398064
rect 357216 398052 357222 398064
rect 357342 398052 357348 398064
rect 357216 398024 357348 398052
rect 357216 398012 357222 398024
rect 357342 398012 357348 398024
rect 357400 398012 357406 398064
rect 372522 398012 372528 398064
rect 372580 398052 372586 398064
rect 372706 398052 372712 398064
rect 372580 398024 372712 398052
rect 372580 398012 372586 398024
rect 372706 398012 372712 398024
rect 372764 398012 372770 398064
rect 373350 398012 373356 398064
rect 373408 398052 373414 398064
rect 373994 398052 374000 398064
rect 373408 398024 374000 398052
rect 373408 398012 373414 398024
rect 373994 398012 374000 398024
rect 374052 398012 374058 398064
rect 382550 398012 382556 398064
rect 382608 398052 382614 398064
rect 388070 398052 388076 398064
rect 382608 398024 388076 398052
rect 382608 398012 382614 398024
rect 388070 398012 388076 398024
rect 388128 398012 388134 398064
rect 324222 397944 324228 397996
rect 324280 397984 324286 397996
rect 343910 397984 343916 397996
rect 324280 397956 343916 397984
rect 324280 397944 324286 397956
rect 343910 397944 343916 397956
rect 343968 397944 343974 397996
rect 352650 397944 352656 397996
rect 352708 397984 352714 397996
rect 355594 397984 355600 397996
rect 352708 397956 355600 397984
rect 352708 397944 352714 397956
rect 355594 397944 355600 397956
rect 355652 397944 355658 397996
rect 375374 397944 375380 397996
rect 375432 397984 375438 397996
rect 389146 397984 389174 398160
rect 389358 398148 389364 398160
rect 389416 398148 389422 398200
rect 375432 397956 389174 397984
rect 375432 397944 375438 397956
rect 345658 397876 345664 397928
rect 345716 397916 345722 397928
rect 356514 397916 356520 397928
rect 345716 397888 356520 397916
rect 345716 397876 345722 397888
rect 356514 397876 356520 397888
rect 356572 397876 356578 397928
rect 367830 397876 367836 397928
rect 367888 397916 367894 397928
rect 369026 397916 369032 397928
rect 367888 397888 369032 397916
rect 367888 397876 367894 397888
rect 369026 397876 369032 397888
rect 369084 397876 369090 397928
rect 376570 397876 376576 397928
rect 376628 397916 376634 397928
rect 381446 397916 381452 397928
rect 376628 397888 381452 397916
rect 376628 397876 376634 397888
rect 381446 397876 381452 397888
rect 381504 397876 381510 397928
rect 383286 397876 383292 397928
rect 383344 397916 383350 397928
rect 383562 397916 383568 397928
rect 383344 397888 383568 397916
rect 383344 397876 383350 397888
rect 383562 397876 383568 397888
rect 383620 397876 383626 397928
rect 383930 397876 383936 397928
rect 383988 397916 383994 397928
rect 389450 397916 389456 397928
rect 383988 397888 389456 397916
rect 383988 397876 383994 397888
rect 389450 397876 389456 397888
rect 389508 397876 389514 397928
rect 343726 397808 343732 397860
rect 343784 397848 343790 397860
rect 346578 397848 346584 397860
rect 343784 397820 346584 397848
rect 343784 397808 343790 397820
rect 346578 397808 346584 397820
rect 346636 397808 346642 397860
rect 352742 397808 352748 397860
rect 352800 397848 352806 397860
rect 352926 397848 352932 397860
rect 352800 397820 352932 397848
rect 352800 397808 352806 397820
rect 352926 397808 352932 397820
rect 352984 397808 352990 397860
rect 359366 397848 359372 397860
rect 353266 397820 359372 397848
rect 337746 397740 337752 397792
rect 337804 397780 337810 397792
rect 353266 397780 353294 397820
rect 359366 397808 359372 397820
rect 359424 397808 359430 397860
rect 362862 397808 362868 397860
rect 362920 397848 362926 397860
rect 365806 397848 365812 397860
rect 362920 397820 365812 397848
rect 362920 397808 362926 397820
rect 365806 397808 365812 397820
rect 365864 397808 365870 397860
rect 376202 397808 376208 397860
rect 376260 397848 376266 397860
rect 376260 397820 380894 397848
rect 376260 397808 376266 397820
rect 362034 397780 362040 397792
rect 337804 397752 353294 397780
rect 356256 397752 362040 397780
rect 337804 397740 337810 397752
rect 339126 397672 339132 397724
rect 339184 397712 339190 397724
rect 345658 397712 345664 397724
rect 339184 397684 345664 397712
rect 339184 397672 339190 397684
rect 345658 397672 345664 397684
rect 345716 397672 345722 397724
rect 345842 397672 345848 397724
rect 345900 397712 345906 397724
rect 346210 397712 346216 397724
rect 345900 397684 346216 397712
rect 345900 397672 345906 397684
rect 346210 397672 346216 397684
rect 346268 397672 346274 397724
rect 346578 397672 346584 397724
rect 346636 397712 346642 397724
rect 356256 397712 356284 397752
rect 362034 397740 362040 397752
rect 362092 397740 362098 397792
rect 380866 397780 380894 397820
rect 384482 397808 384488 397860
rect 384540 397848 384546 397860
rect 390922 397848 390928 397860
rect 384540 397820 390928 397848
rect 384540 397808 384546 397820
rect 390922 397808 390928 397820
rect 390980 397808 390986 397860
rect 383562 397780 383568 397792
rect 380866 397752 383568 397780
rect 383562 397740 383568 397752
rect 383620 397740 383626 397792
rect 384206 397740 384212 397792
rect 384264 397780 384270 397792
rect 387886 397780 387892 397792
rect 384264 397752 387892 397780
rect 384264 397740 384270 397752
rect 387886 397740 387892 397752
rect 387944 397740 387950 397792
rect 346636 397684 356284 397712
rect 346636 397672 346642 397684
rect 356330 397672 356336 397724
rect 356388 397712 356394 397724
rect 363690 397712 363696 397724
rect 356388 397684 363696 397712
rect 356388 397672 356394 397684
rect 363690 397672 363696 397684
rect 363748 397672 363754 397724
rect 364150 397672 364156 397724
rect 364208 397712 364214 397724
rect 368658 397712 368664 397724
rect 364208 397684 368664 397712
rect 364208 397672 364214 397684
rect 368658 397672 368664 397684
rect 368716 397672 368722 397724
rect 384666 397672 384672 397724
rect 384724 397712 384730 397724
rect 392302 397712 392308 397724
rect 384724 397684 392308 397712
rect 384724 397672 384730 397684
rect 392302 397672 392308 397684
rect 392360 397672 392366 397724
rect 278498 397604 278504 397656
rect 278556 397644 278562 397656
rect 356606 397644 356612 397656
rect 278556 397616 356612 397644
rect 278556 397604 278562 397616
rect 356606 397604 356612 397616
rect 356664 397604 356670 397656
rect 356790 397604 356796 397656
rect 356848 397644 356854 397656
rect 357158 397644 357164 397656
rect 356848 397616 357164 397644
rect 356848 397604 356854 397616
rect 357158 397604 357164 397616
rect 357216 397604 357222 397656
rect 366542 397604 366548 397656
rect 366600 397644 366606 397656
rect 370406 397644 370412 397656
rect 366600 397616 370412 397644
rect 366600 397604 366606 397616
rect 370406 397604 370412 397616
rect 370464 397604 370470 397656
rect 386690 397604 386696 397656
rect 386748 397644 386754 397656
rect 393130 397644 393136 397656
rect 386748 397616 393136 397644
rect 386748 397604 386754 397616
rect 393130 397604 393136 397616
rect 393188 397604 393194 397656
rect 343818 397536 343824 397588
rect 343876 397576 343882 397588
rect 343876 397548 345060 397576
rect 343876 397536 343882 397548
rect 3418 397468 3424 397520
rect 3476 397508 3482 397520
rect 256878 397508 256884 397520
rect 3476 397480 256884 397508
rect 3476 397468 3482 397480
rect 256878 397468 256884 397480
rect 256936 397508 256942 397520
rect 307662 397508 307668 397520
rect 256936 397480 307668 397508
rect 256936 397468 256942 397480
rect 307662 397468 307668 397480
rect 307720 397468 307726 397520
rect 345032 397508 345060 397548
rect 347866 397536 347872 397588
rect 347924 397576 347930 397588
rect 348878 397576 348884 397588
rect 347924 397548 348884 397576
rect 347924 397536 347930 397548
rect 348878 397536 348884 397548
rect 348936 397536 348942 397588
rect 350810 397536 350816 397588
rect 350868 397576 350874 397588
rect 351270 397576 351276 397588
rect 350868 397548 351276 397576
rect 350868 397536 350874 397548
rect 351270 397536 351276 397548
rect 351328 397536 351334 397588
rect 351914 397536 351920 397588
rect 351972 397576 351978 397588
rect 352190 397576 352196 397588
rect 351972 397548 352196 397576
rect 351972 397536 351978 397548
rect 352190 397536 352196 397548
rect 352248 397536 352254 397588
rect 356882 397536 356888 397588
rect 356940 397576 356946 397588
rect 357342 397576 357348 397588
rect 356940 397548 357348 397576
rect 356940 397536 356946 397548
rect 357342 397536 357348 397548
rect 357400 397536 357406 397588
rect 365806 397536 365812 397588
rect 365864 397576 365870 397588
rect 365864 397548 367094 397576
rect 365864 397536 365870 397548
rect 346578 397508 346584 397520
rect 345032 397480 346584 397508
rect 346578 397468 346584 397480
rect 346636 397468 346642 397520
rect 348142 397468 348148 397520
rect 348200 397508 348206 397520
rect 348602 397508 348608 397520
rect 348200 397480 348608 397508
rect 348200 397468 348206 397480
rect 348602 397468 348608 397480
rect 348660 397468 348666 397520
rect 351178 397468 351184 397520
rect 351236 397508 351242 397520
rect 352374 397508 352380 397520
rect 351236 397480 352380 397508
rect 351236 397468 351242 397480
rect 352374 397468 352380 397480
rect 352432 397468 352438 397520
rect 352742 397468 352748 397520
rect 352800 397508 352806 397520
rect 354582 397508 354588 397520
rect 352800 397480 354588 397508
rect 352800 397468 352806 397480
rect 354582 397468 354588 397480
rect 354640 397468 354646 397520
rect 356606 397468 356612 397520
rect 356664 397508 356670 397520
rect 360194 397508 360200 397520
rect 356664 397480 360200 397508
rect 356664 397468 356670 397480
rect 360194 397468 360200 397480
rect 360252 397468 360258 397520
rect 367066 397508 367094 397548
rect 386782 397536 386788 397588
rect 386840 397576 386846 397588
rect 391934 397576 391940 397588
rect 386840 397548 391940 397576
rect 386840 397536 386846 397548
rect 391934 397536 391940 397548
rect 391992 397536 391998 397588
rect 369118 397508 369124 397520
rect 367066 397480 369124 397508
rect 369118 397468 369124 397480
rect 369176 397468 369182 397520
rect 370774 397468 370780 397520
rect 370832 397508 370838 397520
rect 372614 397508 372620 397520
rect 370832 397480 372620 397508
rect 370832 397468 370838 397480
rect 372614 397468 372620 397480
rect 372672 397468 372678 397520
rect 383654 397468 383660 397520
rect 383712 397508 383718 397520
rect 384390 397508 384396 397520
rect 383712 397480 384396 397508
rect 383712 397468 383718 397480
rect 384390 397468 384396 397480
rect 384448 397468 384454 397520
rect 385862 397468 385868 397520
rect 385920 397508 385926 397520
rect 390738 397508 390744 397520
rect 385920 397480 390744 397508
rect 385920 397468 385926 397480
rect 390738 397468 390744 397480
rect 390796 397468 390802 397520
rect 343082 397400 343088 397452
rect 343140 397440 343146 397452
rect 346946 397440 346952 397452
rect 343140 397412 346952 397440
rect 343140 397400 343146 397412
rect 346946 397400 346952 397412
rect 347004 397400 347010 397452
rect 348510 397400 348516 397452
rect 348568 397440 348574 397452
rect 348878 397440 348884 397452
rect 348568 397412 348884 397440
rect 348568 397400 348574 397412
rect 348878 397400 348884 397412
rect 348936 397400 348942 397452
rect 350166 397400 350172 397452
rect 350224 397440 350230 397452
rect 360746 397440 360752 397452
rect 350224 397412 360752 397440
rect 350224 397400 350230 397412
rect 360746 397400 360752 397412
rect 360804 397400 360810 397452
rect 369486 397400 369492 397452
rect 369544 397440 369550 397452
rect 374546 397440 374552 397452
rect 369544 397412 374552 397440
rect 369544 397400 369550 397412
rect 374546 397400 374552 397412
rect 374604 397400 374610 397452
rect 377306 397400 377312 397452
rect 377364 397440 377370 397452
rect 386046 397440 386052 397452
rect 377364 397412 386052 397440
rect 377364 397400 377370 397412
rect 386046 397400 386052 397412
rect 386104 397400 386110 397452
rect 341150 397332 341156 397384
rect 341208 397372 341214 397384
rect 344002 397372 344008 397384
rect 341208 397344 344008 397372
rect 341208 397332 341214 397344
rect 344002 397332 344008 397344
rect 344060 397332 344066 397384
rect 345658 397332 345664 397384
rect 345716 397372 345722 397384
rect 356606 397372 356612 397384
rect 345716 397344 356612 397372
rect 345716 397332 345722 397344
rect 356606 397332 356612 397344
rect 356664 397332 356670 397384
rect 357342 397332 357348 397384
rect 357400 397372 357406 397384
rect 358446 397372 358452 397384
rect 357400 397344 358452 397372
rect 357400 397332 357406 397344
rect 358446 397332 358452 397344
rect 358504 397332 358510 397384
rect 364978 397332 364984 397384
rect 365036 397372 365042 397384
rect 366266 397372 366272 397384
rect 365036 397344 366272 397372
rect 365036 397332 365042 397344
rect 366266 397332 366272 397344
rect 366324 397332 366330 397384
rect 366450 397332 366456 397384
rect 366508 397372 366514 397384
rect 366726 397372 366732 397384
rect 366508 397344 366732 397372
rect 366508 397332 366514 397344
rect 366726 397332 366732 397344
rect 366784 397332 366790 397384
rect 367002 397332 367008 397384
rect 367060 397372 367066 397384
rect 369854 397372 369860 397384
rect 367060 397344 369860 397372
rect 367060 397332 367066 397344
rect 369854 397332 369860 397344
rect 369912 397332 369918 397384
rect 386690 397332 386696 397384
rect 386748 397372 386754 397384
rect 387334 397372 387340 397384
rect 386748 397344 387340 397372
rect 386748 397332 386754 397344
rect 387334 397332 387340 397344
rect 387392 397332 387398 397384
rect 334802 397264 334808 397316
rect 334860 397304 334866 397316
rect 356146 397304 356152 397316
rect 334860 397276 356152 397304
rect 334860 397264 334866 397276
rect 356146 397264 356152 397276
rect 356204 397264 356210 397316
rect 356790 397264 356796 397316
rect 356848 397304 356854 397316
rect 359458 397304 359464 397316
rect 356848 397276 359464 397304
rect 356848 397264 356854 397276
rect 359458 397264 359464 397276
rect 359516 397264 359522 397316
rect 382274 397264 382280 397316
rect 382332 397304 382338 397316
rect 383194 397304 383200 397316
rect 382332 397276 383200 397304
rect 382332 397264 382338 397276
rect 383194 397264 383200 397276
rect 383252 397264 383258 397316
rect 333422 397196 333428 397248
rect 333480 397236 333486 397248
rect 358906 397236 358912 397248
rect 333480 397208 358912 397236
rect 333480 397196 333486 397208
rect 358906 397196 358912 397208
rect 358964 397196 358970 397248
rect 360470 397196 360476 397248
rect 360528 397236 360534 397248
rect 361206 397236 361212 397248
rect 360528 397208 361212 397236
rect 360528 397196 360534 397208
rect 361206 397196 361212 397208
rect 361264 397196 361270 397248
rect 337470 397128 337476 397180
rect 337528 397168 337534 397180
rect 364426 397168 364432 397180
rect 337528 397140 364432 397168
rect 337528 397128 337534 397140
rect 364426 397128 364432 397140
rect 364484 397128 364490 397180
rect 337562 397060 337568 397112
rect 337620 397100 337626 397112
rect 370130 397100 370136 397112
rect 337620 397072 370136 397100
rect 337620 397060 337626 397072
rect 370130 397060 370136 397072
rect 370188 397060 370194 397112
rect 333238 396992 333244 397044
rect 333296 397032 333302 397044
rect 366818 397032 366824 397044
rect 333296 397004 366824 397032
rect 333296 396992 333302 397004
rect 366818 396992 366824 397004
rect 366876 396992 366882 397044
rect 329098 396924 329104 396976
rect 329156 396964 329162 396976
rect 368106 396964 368112 396976
rect 329156 396936 368112 396964
rect 329156 396924 329162 396936
rect 368106 396924 368112 396936
rect 368164 396924 368170 396976
rect 381538 396964 381544 396976
rect 369826 396936 381544 396964
rect 336642 396856 336648 396908
rect 336700 396896 336706 396908
rect 369826 396896 369854 396936
rect 381538 396924 381544 396936
rect 381596 396924 381602 396976
rect 336700 396868 369854 396896
rect 336700 396856 336706 396868
rect 281534 396788 281540 396840
rect 281592 396828 281598 396840
rect 295334 396828 295340 396840
rect 281592 396800 295340 396828
rect 281592 396788 281598 396800
rect 295334 396788 295340 396800
rect 295392 396788 295398 396840
rect 340414 396788 340420 396840
rect 340472 396828 340478 396840
rect 385402 396828 385408 396840
rect 340472 396800 385408 396828
rect 340472 396788 340478 396800
rect 385402 396788 385408 396800
rect 385460 396788 385466 396840
rect 270126 396720 270132 396772
rect 270184 396760 270190 396772
rect 346118 396760 346124 396772
rect 270184 396732 346124 396760
rect 270184 396720 270190 396732
rect 346118 396720 346124 396732
rect 346176 396720 346182 396772
rect 348510 396720 348516 396772
rect 348568 396760 348574 396772
rect 349890 396760 349896 396772
rect 348568 396732 349896 396760
rect 348568 396720 348574 396732
rect 349890 396720 349896 396732
rect 349948 396720 349954 396772
rect 359458 396720 359464 396772
rect 359516 396760 359522 396772
rect 362678 396760 362684 396772
rect 359516 396732 362684 396760
rect 359516 396720 359522 396732
rect 362678 396720 362684 396732
rect 362736 396720 362742 396772
rect 375558 396720 375564 396772
rect 375616 396760 375622 396772
rect 376570 396760 376576 396772
rect 375616 396732 376576 396760
rect 375616 396720 375622 396732
rect 376570 396720 376576 396732
rect 376628 396720 376634 396772
rect 341978 396652 341984 396704
rect 342036 396692 342042 396704
rect 357250 396692 357256 396704
rect 342036 396664 357256 396692
rect 342036 396652 342042 396664
rect 357250 396652 357256 396664
rect 357308 396652 357314 396704
rect 360286 396652 360292 396704
rect 360344 396692 360350 396704
rect 361574 396692 361580 396704
rect 360344 396664 361580 396692
rect 360344 396652 360350 396664
rect 361574 396652 361580 396664
rect 361632 396652 361638 396704
rect 362034 396652 362040 396704
rect 362092 396692 362098 396704
rect 362494 396692 362500 396704
rect 362092 396664 362500 396692
rect 362092 396652 362098 396664
rect 362494 396652 362500 396664
rect 362552 396652 362558 396704
rect 341702 396584 341708 396636
rect 341760 396624 341766 396636
rect 350166 396624 350172 396636
rect 341760 396596 350172 396624
rect 341760 396584 341766 396596
rect 350166 396584 350172 396596
rect 350224 396584 350230 396636
rect 363598 396584 363604 396636
rect 363656 396624 363662 396636
rect 364242 396624 364248 396636
rect 363656 396596 364248 396624
rect 363656 396584 363662 396596
rect 364242 396584 364248 396596
rect 364300 396584 364306 396636
rect 343358 396516 343364 396568
rect 343416 396556 343422 396568
rect 345934 396556 345940 396568
rect 343416 396528 345940 396556
rect 343416 396516 343422 396528
rect 345934 396516 345940 396528
rect 345992 396516 345998 396568
rect 360562 396516 360568 396568
rect 360620 396556 360626 396568
rect 361390 396556 361396 396568
rect 360620 396528 361396 396556
rect 360620 396516 360626 396528
rect 361390 396516 361396 396528
rect 361448 396516 361454 396568
rect 343634 396448 343640 396500
rect 343692 396488 343698 396500
rect 346762 396488 346768 396500
rect 343692 396460 346768 396488
rect 343692 396448 343698 396460
rect 346762 396448 346768 396460
rect 346820 396448 346826 396500
rect 359734 396448 359740 396500
rect 359792 396488 359798 396500
rect 360102 396488 360108 396500
rect 359792 396460 360108 396488
rect 359792 396448 359798 396460
rect 360102 396448 360108 396460
rect 360160 396448 360166 396500
rect 339034 396380 339040 396432
rect 339092 396420 339098 396432
rect 357434 396420 357440 396432
rect 339092 396392 357440 396420
rect 339092 396380 339098 396392
rect 357434 396380 357440 396392
rect 357492 396380 357498 396432
rect 361666 396380 361672 396432
rect 361724 396420 361730 396432
rect 362586 396420 362592 396432
rect 361724 396392 362592 396420
rect 361724 396380 361730 396392
rect 362586 396380 362592 396392
rect 362644 396380 362650 396432
rect 336366 396312 336372 396364
rect 336424 396352 336430 396364
rect 356238 396352 356244 396364
rect 336424 396324 356244 396352
rect 336424 396312 336430 396324
rect 356238 396312 356244 396324
rect 356296 396312 356302 396364
rect 363690 396312 363696 396364
rect 363748 396352 363754 396364
rect 365346 396352 365352 396364
rect 363748 396324 365352 396352
rect 363748 396312 363754 396324
rect 365346 396312 365352 396324
rect 365404 396312 365410 396364
rect 355502 396176 355508 396228
rect 355560 396216 355566 396228
rect 358262 396216 358268 396228
rect 355560 396188 358268 396216
rect 355560 396176 355566 396188
rect 358262 396176 358268 396188
rect 358320 396176 358326 396228
rect 377306 396176 377312 396228
rect 377364 396216 377370 396228
rect 378226 396216 378232 396228
rect 377364 396188 378232 396216
rect 377364 396176 377370 396188
rect 378226 396176 378232 396188
rect 378284 396176 378290 396228
rect 340230 396108 340236 396160
rect 340288 396148 340294 396160
rect 345658 396148 345664 396160
rect 340288 396120 345664 396148
rect 340288 396108 340294 396120
rect 345658 396108 345664 396120
rect 345716 396108 345722 396160
rect 345842 396040 345848 396092
rect 345900 396080 345906 396092
rect 346026 396080 346032 396092
rect 345900 396052 346032 396080
rect 345900 396040 345906 396052
rect 346026 396040 346032 396052
rect 346084 396040 346090 396092
rect 355594 396040 355600 396092
rect 355652 396080 355658 396092
rect 356974 396080 356980 396092
rect 355652 396052 356980 396080
rect 355652 396040 355658 396052
rect 356974 396040 356980 396052
rect 357032 396040 357038 396092
rect 358262 396040 358268 396092
rect 358320 396080 358326 396092
rect 359090 396080 359096 396092
rect 358320 396052 359096 396080
rect 358320 396040 358326 396052
rect 359090 396040 359096 396052
rect 359148 396040 359154 396092
rect 377398 396040 377404 396092
rect 377456 396080 377462 396092
rect 384666 396080 384672 396092
rect 377456 396052 384672 396080
rect 377456 396040 377462 396052
rect 384666 396040 384672 396052
rect 384724 396040 384730 396092
rect 338758 395972 338764 396024
rect 338816 396012 338822 396024
rect 362862 396012 362868 396024
rect 338816 395984 362868 396012
rect 338816 395972 338822 395984
rect 362862 395972 362868 395984
rect 362920 395972 362926 396024
rect 341794 395904 341800 395956
rect 341852 395944 341858 395956
rect 343542 395944 343548 395956
rect 341852 395916 343548 395944
rect 341852 395904 341858 395916
rect 343542 395904 343548 395916
rect 343600 395904 343606 395956
rect 345842 395904 345848 395956
rect 345900 395944 345906 395956
rect 364886 395944 364892 395956
rect 345900 395916 364892 395944
rect 345900 395904 345906 395916
rect 364886 395904 364892 395916
rect 364944 395904 364950 395956
rect 377858 395904 377864 395956
rect 377916 395944 377922 395956
rect 384206 395944 384212 395956
rect 377916 395916 384212 395944
rect 377916 395904 377922 395916
rect 384206 395904 384212 395916
rect 384264 395904 384270 395956
rect 341334 395836 341340 395888
rect 341392 395876 341398 395888
rect 370682 395876 370688 395888
rect 341392 395848 370688 395876
rect 341392 395836 341398 395848
rect 370682 395836 370688 395848
rect 370740 395836 370746 395888
rect 340322 395768 340328 395820
rect 340380 395808 340386 395820
rect 370958 395808 370964 395820
rect 340380 395780 370964 395808
rect 340380 395768 340386 395780
rect 370958 395768 370964 395780
rect 371016 395768 371022 395820
rect 331858 395700 331864 395752
rect 331916 395740 331922 395752
rect 360838 395740 360844 395752
rect 331916 395712 360844 395740
rect 331916 395700 331922 395712
rect 360838 395700 360844 395712
rect 360896 395700 360902 395752
rect 330938 395632 330944 395684
rect 330996 395672 331002 395684
rect 368014 395672 368020 395684
rect 330996 395644 368020 395672
rect 330996 395632 331002 395644
rect 368014 395632 368020 395644
rect 368072 395632 368078 395684
rect 374730 395632 374736 395684
rect 374788 395672 374794 395684
rect 378686 395672 378692 395684
rect 374788 395644 378692 395672
rect 374788 395632 374794 395644
rect 378686 395632 378692 395644
rect 378744 395632 378750 395684
rect 344186 395564 344192 395616
rect 344244 395604 344250 395616
rect 345014 395604 345020 395616
rect 344244 395576 345020 395604
rect 344244 395564 344250 395576
rect 345014 395564 345020 395576
rect 345072 395564 345078 395616
rect 345290 395564 345296 395616
rect 345348 395604 345354 395616
rect 345566 395604 345572 395616
rect 345348 395576 345572 395604
rect 345348 395564 345354 395576
rect 345566 395564 345572 395576
rect 345624 395564 345630 395616
rect 345658 395564 345664 395616
rect 345716 395604 345722 395616
rect 385310 395604 385316 395616
rect 345716 395576 385316 395604
rect 345716 395564 345722 395576
rect 385310 395564 385316 395576
rect 385368 395564 385374 395616
rect 272978 395496 272984 395548
rect 273036 395536 273042 395548
rect 334894 395536 334900 395548
rect 273036 395508 334900 395536
rect 273036 395496 273042 395508
rect 334894 395496 334900 395508
rect 334952 395496 334958 395548
rect 271598 395428 271604 395480
rect 271656 395468 271662 395480
rect 343358 395468 343364 395480
rect 271656 395440 343364 395468
rect 271656 395428 271662 395440
rect 343358 395428 343364 395440
rect 343416 395428 343422 395480
rect 376386 395428 376392 395480
rect 376444 395468 376450 395480
rect 378686 395468 378692 395480
rect 376444 395440 378692 395468
rect 376444 395428 376450 395440
rect 378686 395428 378692 395440
rect 378744 395428 378750 395480
rect 379054 395428 379060 395480
rect 379112 395468 379118 395480
rect 379790 395468 379796 395480
rect 379112 395440 379796 395468
rect 379112 395428 379118 395440
rect 379790 395428 379796 395440
rect 379848 395428 379854 395480
rect 268470 395360 268476 395412
rect 268528 395400 268534 395412
rect 334342 395400 334348 395412
rect 268528 395372 334348 395400
rect 268528 395360 268534 395372
rect 334342 395360 334348 395372
rect 334400 395360 334406 395412
rect 343910 395360 343916 395412
rect 343968 395400 343974 395412
rect 344370 395400 344376 395412
rect 343968 395372 344376 395400
rect 343968 395360 343974 395372
rect 344370 395360 344376 395372
rect 344428 395360 344434 395412
rect 345198 395360 345204 395412
rect 345256 395400 345262 395412
rect 345750 395400 345756 395412
rect 345256 395372 345756 395400
rect 345256 395360 345262 395372
rect 345750 395360 345756 395372
rect 345808 395360 345814 395412
rect 357710 395360 357716 395412
rect 357768 395400 357774 395412
rect 357894 395400 357900 395412
rect 357768 395372 357900 395400
rect 357768 395360 357774 395372
rect 357894 395360 357900 395372
rect 357952 395360 357958 395412
rect 361114 395360 361120 395412
rect 361172 395400 361178 395412
rect 369946 395400 369952 395412
rect 361172 395372 369952 395400
rect 361172 395360 361178 395372
rect 369946 395360 369952 395372
rect 370004 395360 370010 395412
rect 376662 395360 376668 395412
rect 376720 395400 376726 395412
rect 376938 395400 376944 395412
rect 376720 395372 376944 395400
rect 376720 395360 376726 395372
rect 376938 395360 376944 395372
rect 376996 395360 377002 395412
rect 378318 395360 378324 395412
rect 378376 395400 378382 395412
rect 380250 395400 380256 395412
rect 378376 395372 380256 395400
rect 378376 395360 378382 395372
rect 380250 395360 380256 395372
rect 380308 395360 380314 395412
rect 274358 395292 274364 395344
rect 274416 395332 274422 395344
rect 367646 395332 367652 395344
rect 274416 395304 367652 395332
rect 274416 395292 274422 395304
rect 367646 395292 367652 395304
rect 367704 395292 367710 395344
rect 371786 395292 371792 395344
rect 371844 395332 371850 395344
rect 376754 395332 376760 395344
rect 371844 395304 376760 395332
rect 371844 395292 371850 395304
rect 376754 395292 376760 395304
rect 376812 395292 376818 395344
rect 378502 395292 378508 395344
rect 378560 395332 378566 395344
rect 379422 395332 379428 395344
rect 378560 395304 379428 395332
rect 378560 395292 378566 395304
rect 379422 395292 379428 395304
rect 379480 395292 379486 395344
rect 379790 395292 379796 395344
rect 379848 395332 379854 395344
rect 380342 395332 380348 395344
rect 379848 395304 380348 395332
rect 379848 395292 379854 395304
rect 380342 395292 380348 395304
rect 380400 395292 380406 395344
rect 383286 395292 383292 395344
rect 383344 395332 383350 395344
rect 394786 395332 394792 395344
rect 383344 395304 394792 395332
rect 383344 395292 383350 395304
rect 394786 395292 394792 395304
rect 394844 395292 394850 395344
rect 338666 395224 338672 395276
rect 338724 395264 338730 395276
rect 345658 395264 345664 395276
rect 338724 395236 345664 395264
rect 338724 395224 338730 395236
rect 345658 395224 345664 395236
rect 345716 395224 345722 395276
rect 348234 395224 348240 395276
rect 348292 395264 348298 395276
rect 348786 395264 348792 395276
rect 348292 395236 348792 395264
rect 348292 395224 348298 395236
rect 348786 395224 348792 395236
rect 348844 395224 348850 395276
rect 376386 395224 376392 395276
rect 376444 395264 376450 395276
rect 378134 395264 378140 395276
rect 376444 395236 378140 395264
rect 376444 395224 376450 395236
rect 378134 395224 378140 395236
rect 378192 395224 378198 395276
rect 339954 395156 339960 395208
rect 340012 395196 340018 395208
rect 353478 395196 353484 395208
rect 340012 395168 353484 395196
rect 340012 395156 340018 395168
rect 353478 395156 353484 395168
rect 353536 395156 353542 395208
rect 356790 395156 356796 395208
rect 356848 395196 356854 395208
rect 358630 395196 358636 395208
rect 356848 395168 358636 395196
rect 356848 395156 356854 395168
rect 358630 395156 358636 395168
rect 358688 395156 358694 395208
rect 281626 395088 281632 395140
rect 281684 395128 281690 395140
rect 282914 395128 282920 395140
rect 281684 395100 282920 395128
rect 281684 395088 281690 395100
rect 282914 395088 282920 395100
rect 282972 395088 282978 395140
rect 336090 395088 336096 395140
rect 336148 395128 336154 395140
rect 353754 395128 353760 395140
rect 336148 395100 353760 395128
rect 336148 395088 336154 395100
rect 353754 395088 353760 395100
rect 353812 395088 353818 395140
rect 362126 395088 362132 395140
rect 362184 395128 362190 395140
rect 365714 395128 365720 395140
rect 362184 395100 365720 395128
rect 362184 395088 362190 395100
rect 365714 395088 365720 395100
rect 365772 395088 365778 395140
rect 375650 395088 375656 395140
rect 375708 395088 375714 395140
rect 378134 395088 378140 395140
rect 378192 395128 378198 395140
rect 378778 395128 378784 395140
rect 378192 395100 378784 395128
rect 378192 395088 378198 395100
rect 378778 395088 378784 395100
rect 378836 395088 378842 395140
rect 335998 395020 336004 395072
rect 336056 395060 336062 395072
rect 345842 395060 345848 395072
rect 336056 395032 345848 395060
rect 336056 395020 336062 395032
rect 345842 395020 345848 395032
rect 345900 395020 345906 395072
rect 346486 395020 346492 395072
rect 346544 395060 346550 395072
rect 346670 395060 346676 395072
rect 346544 395032 346676 395060
rect 346544 395020 346550 395032
rect 346670 395020 346676 395032
rect 346728 395020 346734 395072
rect 346762 395020 346768 395072
rect 346820 395060 346826 395072
rect 347590 395060 347596 395072
rect 346820 395032 347596 395060
rect 346820 395020 346826 395032
rect 347590 395020 347596 395032
rect 347648 395020 347654 395072
rect 345382 394952 345388 395004
rect 345440 394992 345446 395004
rect 346302 394992 346308 395004
rect 345440 394964 346308 394992
rect 345440 394952 345446 394964
rect 346302 394952 346308 394964
rect 346360 394952 346366 395004
rect 375668 394936 375696 395088
rect 375650 394884 375656 394936
rect 375708 394884 375714 394936
rect 386322 394884 386328 394936
rect 386380 394924 386386 394936
rect 394878 394924 394884 394936
rect 386380 394896 394884 394924
rect 386380 394884 386386 394896
rect 394878 394884 394884 394896
rect 394936 394884 394942 394936
rect 342898 394816 342904 394868
rect 342956 394856 342962 394868
rect 349154 394856 349160 394868
rect 342956 394828 349160 394856
rect 342956 394816 342962 394828
rect 349154 394816 349160 394828
rect 349212 394816 349218 394868
rect 393130 394748 393136 394800
rect 393188 394788 393194 394800
rect 394694 394788 394700 394800
rect 393188 394760 394700 394788
rect 393188 394748 393194 394760
rect 394694 394748 394700 394760
rect 394752 394748 394758 394800
rect 366450 394680 366456 394732
rect 366508 394720 366514 394732
rect 367094 394720 367100 394732
rect 366508 394692 367100 394720
rect 366508 394680 366514 394692
rect 367094 394680 367100 394692
rect 367152 394680 367158 394732
rect 370498 394680 370504 394732
rect 370556 394720 370562 394732
rect 371234 394720 371240 394732
rect 370556 394692 371240 394720
rect 370556 394680 370562 394692
rect 371234 394680 371240 394692
rect 371292 394680 371298 394732
rect 381538 394680 381544 394732
rect 381596 394720 381602 394732
rect 384298 394720 384304 394732
rect 381596 394692 384304 394720
rect 381596 394680 381602 394692
rect 384298 394680 384304 394692
rect 384356 394680 384362 394732
rect 307662 394612 307668 394664
rect 307720 394652 307726 394664
rect 316310 394652 316316 394664
rect 307720 394624 316316 394652
rect 307720 394612 307726 394624
rect 316310 394612 316316 394624
rect 316368 394652 316374 394664
rect 316678 394652 316684 394664
rect 316368 394624 316684 394652
rect 316368 394612 316374 394624
rect 316678 394612 316684 394624
rect 316736 394612 316742 394664
rect 363230 394612 363236 394664
rect 363288 394652 363294 394664
rect 364702 394652 364708 394664
rect 363288 394624 364708 394652
rect 363288 394612 363294 394624
rect 364702 394612 364708 394624
rect 364760 394612 364766 394664
rect 342530 394544 342536 394596
rect 342588 394584 342594 394596
rect 342990 394584 342996 394596
rect 342588 394556 342996 394584
rect 342588 394544 342594 394556
rect 342990 394544 342996 394556
rect 343048 394544 343054 394596
rect 363138 394544 363144 394596
rect 363196 394584 363202 394596
rect 363322 394584 363328 394596
rect 363196 394556 363328 394584
rect 363196 394544 363202 394556
rect 363322 394544 363328 394556
rect 363380 394544 363386 394596
rect 355870 394408 355876 394460
rect 355928 394448 355934 394460
rect 375282 394448 375288 394460
rect 355928 394420 375288 394448
rect 355928 394408 355934 394420
rect 375282 394408 375288 394420
rect 375340 394408 375346 394460
rect 347682 394340 347688 394392
rect 347740 394380 347746 394392
rect 349062 394380 349068 394392
rect 347740 394352 349068 394380
rect 347740 394340 347746 394352
rect 349062 394340 349068 394352
rect 349120 394340 349126 394392
rect 350810 394340 350816 394392
rect 350868 394380 350874 394392
rect 352834 394380 352840 394392
rect 350868 394352 352840 394380
rect 350868 394340 350874 394352
rect 352834 394340 352840 394352
rect 352892 394340 352898 394392
rect 353662 394340 353668 394392
rect 353720 394380 353726 394392
rect 354490 394380 354496 394392
rect 353720 394352 354496 394380
rect 353720 394340 353726 394352
rect 354490 394340 354496 394352
rect 354548 394340 354554 394392
rect 354582 394340 354588 394392
rect 354640 394380 354646 394392
rect 377030 394380 377036 394392
rect 354640 394352 377036 394380
rect 354640 394340 354646 394352
rect 377030 394340 377036 394352
rect 377088 394340 377094 394392
rect 340598 394272 340604 394324
rect 340656 394312 340662 394324
rect 366726 394312 366732 394324
rect 340656 394284 366732 394312
rect 340656 394272 340662 394284
rect 366726 394272 366732 394284
rect 366784 394272 366790 394324
rect 374270 394272 374276 394324
rect 374328 394312 374334 394324
rect 374638 394312 374644 394324
rect 374328 394284 374644 394312
rect 374328 394272 374334 394284
rect 374638 394272 374644 394284
rect 374696 394272 374702 394324
rect 332134 394204 332140 394256
rect 332192 394244 332198 394256
rect 367922 394244 367928 394256
rect 332192 394216 367928 394244
rect 332192 394204 332198 394216
rect 367922 394204 367928 394216
rect 367980 394204 367986 394256
rect 371234 394204 371240 394256
rect 371292 394244 371298 394256
rect 371510 394244 371516 394256
rect 371292 394216 371516 394244
rect 371292 394204 371298 394216
rect 371510 394204 371516 394216
rect 371568 394204 371574 394256
rect 374362 394204 374368 394256
rect 374420 394244 374426 394256
rect 375282 394244 375288 394256
rect 374420 394216 375288 394244
rect 374420 394204 374426 394216
rect 375282 394204 375288 394216
rect 375340 394204 375346 394256
rect 321370 394136 321376 394188
rect 321428 394176 321434 394188
rect 381078 394176 381084 394188
rect 321428 394148 381084 394176
rect 321428 394136 321434 394148
rect 381078 394136 381084 394148
rect 381136 394136 381142 394188
rect 383838 394136 383844 394188
rect 383896 394136 383902 394188
rect 268838 394068 268844 394120
rect 268896 394108 268902 394120
rect 350810 394108 350816 394120
rect 268896 394080 350816 394108
rect 268896 394068 268902 394080
rect 350810 394068 350816 394080
rect 350868 394068 350874 394120
rect 350994 394068 351000 394120
rect 351052 394108 351058 394120
rect 351638 394108 351644 394120
rect 351052 394080 351644 394108
rect 351052 394068 351058 394080
rect 351638 394068 351644 394080
rect 351696 394068 351702 394120
rect 359550 394068 359556 394120
rect 359608 394108 359614 394120
rect 383102 394108 383108 394120
rect 359608 394080 383108 394108
rect 359608 394068 359614 394080
rect 383102 394068 383108 394080
rect 383160 394068 383166 394120
rect 268746 394000 268752 394052
rect 268804 394040 268810 394052
rect 358170 394040 358176 394052
rect 268804 394012 358176 394040
rect 268804 394000 268810 394012
rect 358170 394000 358176 394012
rect 358228 394000 358234 394052
rect 370222 394000 370228 394052
rect 370280 394040 370286 394052
rect 370866 394040 370872 394052
rect 370280 394012 370872 394040
rect 370280 394000 370286 394012
rect 370866 394000 370872 394012
rect 370924 394000 370930 394052
rect 371510 394000 371516 394052
rect 371568 394040 371574 394052
rect 371878 394040 371884 394052
rect 371568 394012 371884 394040
rect 371568 394000 371574 394012
rect 371878 394000 371884 394012
rect 371936 394000 371942 394052
rect 377214 394000 377220 394052
rect 377272 394040 377278 394052
rect 377858 394040 377864 394052
rect 377272 394012 377864 394040
rect 377272 394000 377278 394012
rect 377858 394000 377864 394012
rect 377916 394000 377922 394052
rect 382550 394000 382556 394052
rect 382608 394040 382614 394052
rect 383378 394040 383384 394052
rect 382608 394012 383384 394040
rect 382608 394000 382614 394012
rect 383378 394000 383384 394012
rect 383436 394000 383442 394052
rect 267366 393932 267372 393984
rect 267424 393972 267430 393984
rect 267424 393944 350534 393972
rect 267424 393932 267430 393944
rect 343174 393864 343180 393916
rect 343232 393904 343238 393916
rect 343450 393904 343456 393916
rect 343232 393876 343456 393904
rect 343232 393864 343238 393876
rect 343450 393864 343456 393876
rect 343508 393864 343514 393916
rect 350506 393904 350534 393944
rect 350810 393932 350816 393984
rect 350868 393972 350874 393984
rect 351362 393972 351368 393984
rect 350868 393944 351368 393972
rect 350868 393932 350874 393944
rect 351362 393932 351368 393944
rect 351420 393932 351426 393984
rect 353386 393932 353392 393984
rect 353444 393972 353450 393984
rect 354122 393972 354128 393984
rect 353444 393944 354128 393972
rect 353444 393932 353450 393944
rect 354122 393932 354128 393944
rect 354180 393932 354186 393984
rect 355410 393932 355416 393984
rect 355468 393972 355474 393984
rect 356054 393972 356060 393984
rect 355468 393944 356060 393972
rect 355468 393932 355474 393944
rect 356054 393932 356060 393944
rect 356112 393932 356118 393984
rect 365898 393932 365904 393984
rect 365956 393972 365962 393984
rect 366266 393972 366272 393984
rect 365956 393944 366272 393972
rect 365956 393932 365962 393944
rect 366266 393932 366272 393944
rect 366324 393932 366330 393984
rect 367278 393932 367284 393984
rect 367336 393972 367342 393984
rect 367922 393972 367928 393984
rect 367336 393944 367928 393972
rect 367336 393932 367342 393944
rect 367922 393932 367928 393944
rect 367980 393932 367986 393984
rect 368566 393932 368572 393984
rect 368624 393972 368630 393984
rect 369118 393972 369124 393984
rect 368624 393944 369124 393972
rect 368624 393932 368630 393944
rect 369118 393932 369124 393944
rect 369176 393932 369182 393984
rect 370130 393932 370136 393984
rect 370188 393972 370194 393984
rect 370590 393972 370596 393984
rect 370188 393944 370596 393972
rect 370188 393932 370194 393944
rect 370590 393932 370596 393944
rect 370648 393932 370654 393984
rect 371786 393932 371792 393984
rect 371844 393972 371850 393984
rect 372338 393972 372344 393984
rect 371844 393944 372344 393972
rect 371844 393932 371850 393944
rect 372338 393932 372344 393944
rect 372396 393932 372402 393984
rect 377030 393932 377036 393984
rect 377088 393972 377094 393984
rect 377766 393972 377772 393984
rect 377088 393944 377772 393972
rect 377088 393932 377094 393944
rect 377766 393932 377772 393944
rect 377824 393932 377830 393984
rect 381078 393932 381084 393984
rect 381136 393972 381142 393984
rect 381998 393972 382004 393984
rect 381136 393944 382004 393972
rect 381136 393932 381142 393944
rect 381998 393932 382004 393944
rect 382056 393932 382062 393984
rect 383856 393916 383884 394136
rect 385126 393932 385132 393984
rect 385184 393972 385190 393984
rect 385310 393972 385316 393984
rect 385184 393944 385316 393972
rect 385184 393932 385190 393944
rect 385310 393932 385316 393944
rect 385368 393932 385374 393984
rect 386598 393932 386604 393984
rect 386656 393972 386662 393984
rect 387334 393972 387340 393984
rect 386656 393944 387340 393972
rect 386656 393932 386662 393944
rect 387334 393932 387340 393944
rect 387392 393932 387398 393984
rect 359918 393904 359924 393916
rect 350506 393876 359924 393904
rect 359918 393864 359924 393876
rect 359976 393864 359982 393916
rect 372706 393864 372712 393916
rect 372764 393904 372770 393916
rect 372982 393904 372988 393916
rect 372764 393876 372988 393904
rect 372764 393864 372770 393876
rect 372982 393864 372988 393876
rect 373040 393864 373046 393916
rect 374362 393864 374368 393916
rect 374420 393904 374426 393916
rect 375006 393904 375012 393916
rect 374420 393876 375012 393904
rect 374420 393864 374426 393876
rect 375006 393864 375012 393876
rect 375064 393864 375070 393916
rect 383838 393864 383844 393916
rect 383896 393864 383902 393916
rect 347958 393796 347964 393848
rect 348016 393836 348022 393848
rect 348326 393836 348332 393848
rect 348016 393808 348332 393836
rect 348016 393796 348022 393808
rect 348326 393796 348332 393808
rect 348384 393796 348390 393848
rect 351086 393796 351092 393848
rect 351144 393836 351150 393848
rect 351638 393836 351644 393848
rect 351144 393808 351644 393836
rect 351144 393796 351150 393808
rect 351638 393796 351644 393808
rect 351696 393796 351702 393848
rect 358170 393796 358176 393848
rect 358228 393836 358234 393848
rect 363506 393836 363512 393848
rect 358228 393808 363512 393836
rect 358228 393796 358234 393808
rect 363506 393796 363512 393808
rect 363564 393796 363570 393848
rect 370590 393796 370596 393848
rect 370648 393836 370654 393848
rect 370774 393836 370780 393848
rect 370648 393808 370780 393836
rect 370648 393796 370654 393808
rect 370774 393796 370780 393808
rect 370832 393796 370838 393848
rect 382734 393796 382740 393848
rect 382792 393836 382798 393848
rect 383286 393836 383292 393848
rect 382792 393808 383292 393836
rect 382792 393796 382798 393808
rect 383286 393796 383292 393808
rect 383344 393796 383350 393848
rect 383746 393796 383752 393848
rect 383804 393836 383810 393848
rect 384758 393836 384764 393848
rect 383804 393808 384764 393836
rect 383804 393796 383810 393808
rect 384758 393796 384764 393808
rect 384816 393796 384822 393848
rect 385034 393796 385040 393848
rect 385092 393836 385098 393848
rect 385770 393836 385776 393848
rect 385092 393808 385776 393836
rect 385092 393796 385098 393808
rect 385770 393796 385776 393808
rect 385828 393796 385834 393848
rect 350718 393728 350724 393780
rect 350776 393768 350782 393780
rect 351730 393768 351736 393780
rect 350776 393740 351736 393768
rect 350776 393728 350782 393740
rect 351730 393728 351736 393740
rect 351788 393728 351794 393780
rect 357066 393728 357072 393780
rect 357124 393768 357130 393780
rect 359550 393768 359556 393780
rect 357124 393740 359556 393768
rect 357124 393728 357130 393740
rect 359550 393728 359556 393740
rect 359608 393728 359614 393780
rect 360838 393728 360844 393780
rect 360896 393768 360902 393780
rect 365622 393768 365628 393780
rect 360896 393740 365628 393768
rect 360896 393728 360902 393740
rect 365622 393728 365628 393740
rect 365680 393728 365686 393780
rect 372982 393728 372988 393780
rect 373040 393768 373046 393780
rect 373534 393768 373540 393780
rect 373040 393740 373540 393768
rect 373040 393728 373046 393740
rect 373534 393728 373540 393740
rect 373592 393728 373598 393780
rect 347774 393660 347780 393712
rect 347832 393700 347838 393712
rect 347958 393700 347964 393712
rect 347832 393672 347964 393700
rect 347832 393660 347838 393672
rect 347958 393660 347964 393672
rect 348016 393660 348022 393712
rect 351270 393660 351276 393712
rect 351328 393700 351334 393712
rect 353570 393700 353576 393712
rect 351328 393672 353576 393700
rect 351328 393660 351334 393672
rect 353570 393660 353576 393672
rect 353628 393660 353634 393712
rect 363690 393660 363696 393712
rect 363748 393700 363754 393712
rect 364150 393700 364156 393712
rect 363748 393672 364156 393700
rect 363748 393660 363754 393672
rect 364150 393660 364156 393672
rect 364208 393660 364214 393712
rect 366910 393660 366916 393712
rect 366968 393700 366974 393712
rect 367462 393700 367468 393712
rect 366968 393672 367468 393700
rect 366968 393660 366974 393672
rect 367462 393660 367468 393672
rect 367520 393660 367526 393712
rect 374086 393660 374092 393712
rect 374144 393700 374150 393712
rect 374822 393700 374828 393712
rect 374144 393672 374828 393700
rect 374144 393660 374150 393672
rect 374822 393660 374828 393672
rect 374880 393660 374886 393712
rect 344646 393592 344652 393644
rect 344704 393632 344710 393644
rect 349430 393632 349436 393644
rect 344704 393604 349436 393632
rect 344704 393592 344710 393604
rect 349430 393592 349436 393604
rect 349488 393592 349494 393644
rect 352650 393592 352656 393644
rect 352708 393632 352714 393644
rect 359642 393632 359648 393644
rect 352708 393604 359648 393632
rect 352708 393592 352714 393604
rect 359642 393592 359648 393604
rect 359700 393592 359706 393644
rect 367186 393592 367192 393644
rect 367244 393632 367250 393644
rect 367554 393632 367560 393644
rect 367244 393604 367560 393632
rect 367244 393592 367250 393604
rect 367554 393592 367560 393604
rect 367612 393592 367618 393644
rect 384206 393524 384212 393576
rect 384264 393564 384270 393576
rect 384666 393564 384672 393576
rect 384264 393536 384672 393564
rect 384264 393524 384270 393536
rect 384666 393524 384672 393536
rect 384724 393524 384730 393576
rect 342990 393456 342996 393508
rect 343048 393496 343054 393508
rect 350626 393496 350632 393508
rect 343048 393468 350632 393496
rect 343048 393456 343054 393468
rect 350626 393456 350632 393468
rect 350684 393456 350690 393508
rect 363506 393456 363512 393508
rect 363564 393496 363570 393508
rect 363966 393496 363972 393508
rect 363564 393468 363972 393496
rect 363564 393456 363570 393468
rect 363966 393456 363972 393468
rect 364024 393456 364030 393508
rect 321278 393388 321284 393440
rect 321336 393428 321342 393440
rect 380894 393428 380900 393440
rect 321336 393400 380900 393428
rect 321336 393388 321342 393400
rect 380894 393388 380900 393400
rect 380952 393388 380958 393440
rect 267550 393320 267556 393372
rect 267608 393360 267614 393372
rect 349338 393360 349344 393372
rect 267608 393332 349344 393360
rect 267608 393320 267614 393332
rect 349338 393320 349344 393332
rect 349396 393320 349402 393372
rect 349430 393320 349436 393372
rect 349488 393360 349494 393372
rect 349614 393360 349620 393372
rect 349488 393332 349620 393360
rect 349488 393320 349494 393332
rect 349614 393320 349620 393332
rect 349672 393320 349678 393372
rect 353938 393320 353944 393372
rect 353996 393360 354002 393372
rect 354582 393360 354588 393372
rect 353996 393332 354588 393360
rect 353996 393320 354002 393332
rect 354582 393320 354588 393332
rect 354640 393320 354646 393372
rect 355318 393320 355324 393372
rect 355376 393360 355382 393372
rect 355870 393360 355876 393372
rect 355376 393332 355876 393360
rect 355376 393320 355382 393332
rect 355870 393320 355876 393332
rect 355928 393320 355934 393372
rect 350442 393156 350448 393168
rect 340846 393128 350448 393156
rect 338850 393048 338856 393100
rect 338908 393088 338914 393100
rect 340846 393088 340874 393128
rect 350442 393116 350448 393128
rect 350500 393116 350506 393168
rect 338908 393060 340874 393088
rect 338908 393048 338914 393060
rect 343174 393048 343180 393100
rect 343232 393088 343238 393100
rect 343232 393060 350534 393088
rect 343232 393048 343238 393060
rect 350506 393020 350534 393060
rect 364242 393020 364248 393032
rect 350506 392992 364248 393020
rect 364242 392980 364248 392992
rect 364300 392980 364306 393032
rect 333606 392912 333612 392964
rect 333664 392952 333670 392964
rect 373718 392952 373724 392964
rect 333664 392924 373724 392952
rect 333664 392912 333670 392924
rect 373718 392912 373724 392924
rect 373776 392912 373782 392964
rect 386414 392952 386420 392964
rect 379486 392924 386420 392952
rect 332318 392844 332324 392896
rect 332376 392884 332382 392896
rect 379486 392884 379514 392924
rect 386414 392912 386420 392924
rect 386472 392912 386478 392964
rect 332376 392856 379514 392884
rect 332376 392844 332382 392856
rect 381262 392844 381268 392896
rect 381320 392884 381326 392896
rect 381722 392884 381728 392896
rect 381320 392856 381728 392884
rect 381320 392844 381326 392856
rect 381722 392844 381728 392856
rect 381780 392844 381786 392896
rect 302142 392776 302148 392828
rect 302200 392816 302206 392828
rect 361574 392816 361580 392828
rect 302200 392788 361580 392816
rect 302200 392776 302206 392788
rect 361574 392776 361580 392788
rect 361632 392776 361638 392828
rect 375374 392776 375380 392828
rect 375432 392816 375438 392828
rect 375926 392816 375932 392828
rect 375432 392788 375932 392816
rect 375432 392776 375438 392788
rect 375926 392776 375932 392788
rect 375984 392776 375990 392828
rect 379330 392776 379336 392828
rect 379388 392816 379394 392828
rect 380066 392816 380072 392828
rect 379388 392788 380072 392816
rect 379388 392776 379394 392788
rect 380066 392776 380072 392788
rect 380124 392776 380130 392828
rect 303338 392708 303344 392760
rect 303396 392748 303402 392760
rect 363138 392748 363144 392760
rect 303396 392720 363144 392748
rect 303396 392708 303402 392720
rect 363138 392708 363144 392720
rect 363196 392708 363202 392760
rect 280982 392640 280988 392692
rect 281040 392680 281046 392692
rect 344922 392680 344928 392692
rect 281040 392652 344928 392680
rect 281040 392640 281046 392652
rect 344922 392640 344928 392652
rect 344980 392640 344986 392692
rect 359090 392640 359096 392692
rect 359148 392680 359154 392692
rect 360010 392680 360016 392692
rect 359148 392652 360016 392680
rect 359148 392640 359154 392652
rect 360010 392640 360016 392652
rect 360068 392640 360074 392692
rect 374178 392640 374184 392692
rect 374236 392680 374242 392692
rect 375098 392680 375104 392692
rect 374236 392652 375104 392680
rect 374236 392640 374242 392652
rect 375098 392640 375104 392652
rect 375156 392640 375162 392692
rect 269850 392572 269856 392624
rect 269908 392612 269914 392624
rect 341150 392612 341156 392624
rect 269908 392584 341156 392612
rect 269908 392572 269914 392584
rect 341150 392572 341156 392584
rect 341208 392572 341214 392624
rect 352834 392572 352840 392624
rect 352892 392612 352898 392624
rect 363046 392612 363052 392624
rect 352892 392584 363052 392612
rect 352892 392572 352898 392584
rect 363046 392572 363052 392584
rect 363104 392572 363110 392624
rect 343818 392504 343824 392556
rect 343876 392544 343882 392556
rect 344554 392544 344560 392556
rect 343876 392516 344560 392544
rect 343876 392504 343882 392516
rect 344554 392504 344560 392516
rect 344612 392504 344618 392556
rect 367370 392504 367376 392556
rect 367428 392544 367434 392556
rect 367738 392544 367744 392556
rect 367428 392516 367744 392544
rect 367428 392504 367434 392516
rect 367738 392504 367744 392516
rect 367796 392504 367802 392556
rect 374546 392504 374552 392556
rect 374604 392544 374610 392556
rect 375190 392544 375196 392556
rect 374604 392516 375196 392544
rect 374604 392504 374610 392516
rect 375190 392504 375196 392516
rect 375248 392504 375254 392556
rect 344094 392436 344100 392488
rect 344152 392476 344158 392488
rect 344738 392476 344744 392488
rect 344152 392448 344744 392476
rect 344152 392436 344158 392448
rect 344738 392436 344744 392448
rect 344796 392436 344802 392488
rect 346486 392368 346492 392420
rect 346544 392408 346550 392420
rect 347130 392408 347136 392420
rect 346544 392380 347136 392408
rect 346544 392368 346550 392380
rect 347130 392368 347136 392380
rect 347188 392368 347194 392420
rect 314286 392096 314292 392148
rect 314344 392136 314350 392148
rect 373994 392136 374000 392148
rect 314344 392108 374000 392136
rect 314344 392096 314350 392108
rect 373994 392096 374000 392108
rect 374052 392096 374058 392148
rect 268930 392028 268936 392080
rect 268988 392068 268994 392080
rect 343082 392068 343088 392080
rect 268988 392040 343088 392068
rect 268988 392028 268994 392040
rect 343082 392028 343088 392040
rect 343140 392028 343146 392080
rect 345934 392028 345940 392080
rect 345992 392068 345998 392080
rect 348694 392068 348700 392080
rect 345992 392040 348700 392068
rect 345992 392028 345998 392040
rect 348694 392028 348700 392040
rect 348752 392028 348758 392080
rect 277026 391960 277032 392012
rect 277084 392000 277090 392012
rect 368474 392000 368480 392012
rect 277084 391972 368480 392000
rect 277084 391960 277090 391972
rect 368474 391960 368480 391972
rect 368532 391960 368538 392012
rect 307938 391892 307944 391944
rect 307996 391932 308002 391944
rect 368198 391932 368204 391944
rect 307996 391904 368204 391932
rect 307996 391892 308002 391904
rect 368198 391892 368204 391904
rect 368256 391892 368262 391944
rect 379882 391824 379888 391876
rect 379940 391864 379946 391876
rect 380710 391864 380716 391876
rect 379940 391836 380716 391864
rect 379940 391824 379946 391836
rect 380710 391824 380716 391836
rect 380768 391824 380774 391876
rect 337378 391756 337384 391808
rect 337436 391796 337442 391808
rect 350350 391796 350356 391808
rect 337436 391768 350356 391796
rect 337436 391756 337442 391768
rect 350350 391756 350356 391768
rect 350408 391756 350414 391808
rect 345658 391688 345664 391740
rect 345716 391728 345722 391740
rect 365530 391728 365536 391740
rect 345716 391700 365536 391728
rect 345716 391688 345722 391700
rect 365530 391688 365536 391700
rect 365588 391688 365594 391740
rect 338574 391620 338580 391672
rect 338632 391660 338638 391672
rect 376110 391660 376116 391672
rect 338632 391632 376116 391660
rect 338632 391620 338638 391632
rect 376110 391620 376116 391632
rect 376168 391620 376174 391672
rect 329282 391552 329288 391604
rect 329340 391592 329346 391604
rect 368566 391592 368572 391604
rect 329340 391564 368572 391592
rect 329340 391552 329346 391564
rect 368566 391552 368572 391564
rect 368624 391552 368630 391604
rect 314378 391484 314384 391536
rect 314436 391524 314442 391536
rect 372614 391524 372620 391536
rect 314436 391496 372620 391524
rect 314436 391484 314442 391496
rect 372614 391484 372620 391496
rect 372672 391484 372678 391536
rect 313182 391416 313188 391468
rect 313240 391456 313246 391468
rect 372706 391456 372712 391468
rect 313240 391428 372712 391456
rect 313240 391416 313246 391428
rect 372706 391416 372712 391428
rect 372764 391416 372770 391468
rect 311802 391348 311808 391400
rect 311860 391388 311866 391400
rect 371234 391388 371240 391400
rect 311860 391360 371240 391388
rect 311860 391348 311866 391360
rect 371234 391348 371240 391360
rect 371292 391348 371298 391400
rect 315850 391280 315856 391332
rect 315908 391320 315914 391332
rect 375466 391320 375472 391332
rect 315908 391292 375472 391320
rect 315908 391280 315914 391292
rect 375466 391280 375472 391292
rect 375524 391280 375530 391332
rect 311710 391212 311716 391264
rect 311768 391252 311774 391264
rect 371326 391252 371332 391264
rect 311768 391224 371332 391252
rect 311768 391212 311774 391224
rect 371326 391212 371332 391224
rect 371384 391212 371390 391264
rect 354214 391144 354220 391196
rect 354272 391184 354278 391196
rect 354398 391184 354404 391196
rect 354272 391156 354404 391184
rect 354272 391144 354278 391156
rect 354398 391144 354404 391156
rect 354456 391144 354462 391196
rect 356882 391144 356888 391196
rect 356940 391184 356946 391196
rect 357342 391184 357348 391196
rect 356940 391156 357348 391184
rect 356940 391144 356946 391156
rect 357342 391144 357348 391156
rect 357400 391144 357406 391196
rect 344370 390736 344376 390788
rect 344428 390776 344434 390788
rect 348970 390776 348976 390788
rect 344428 390748 348976 390776
rect 344428 390736 344434 390748
rect 348970 390736 348976 390748
rect 349028 390736 349034 390788
rect 360654 390736 360660 390788
rect 360712 390776 360718 390788
rect 361298 390776 361304 390788
rect 360712 390748 361304 390776
rect 360712 390736 360718 390748
rect 361298 390736 361304 390748
rect 361356 390736 361362 390788
rect 368750 390736 368756 390788
rect 368808 390776 368814 390788
rect 369578 390776 369584 390788
rect 368808 390748 369584 390776
rect 368808 390736 368814 390748
rect 369578 390736 369584 390748
rect 369636 390736 369642 390788
rect 386598 390736 386604 390788
rect 386656 390776 386662 390788
rect 386874 390776 386880 390788
rect 386656 390748 386880 390776
rect 386656 390736 386662 390748
rect 386874 390736 386880 390748
rect 386932 390736 386938 390788
rect 386874 390600 386880 390652
rect 386932 390640 386938 390652
rect 387426 390640 387432 390652
rect 386932 390612 387432 390640
rect 386932 390600 386938 390612
rect 387426 390600 387432 390612
rect 387484 390600 387490 390652
rect 349614 390464 349620 390516
rect 349672 390504 349678 390516
rect 350074 390504 350080 390516
rect 349672 390476 350080 390504
rect 349672 390464 349678 390476
rect 350074 390464 350080 390476
rect 350132 390464 350138 390516
rect 354214 390192 354220 390244
rect 354272 390232 354278 390244
rect 356330 390232 356336 390244
rect 354272 390204 356336 390232
rect 354272 390192 354278 390204
rect 356330 390192 356336 390204
rect 356388 390192 356394 390244
rect 319806 390056 319812 390108
rect 319864 390096 319870 390108
rect 378134 390096 378140 390108
rect 319864 390068 378140 390096
rect 319864 390056 319870 390068
rect 378134 390056 378140 390068
rect 378192 390056 378198 390108
rect 319898 389988 319904 390040
rect 319956 390028 319962 390040
rect 378962 390028 378968 390040
rect 319956 390000 378968 390028
rect 319956 389988 319962 390000
rect 378962 389988 378968 390000
rect 379020 389988 379026 390040
rect 318702 389920 318708 389972
rect 318760 389960 318766 389972
rect 379422 389960 379428 389972
rect 318760 389932 379428 389960
rect 318760 389920 318766 389932
rect 379422 389920 379428 389932
rect 379480 389920 379486 389972
rect 281718 389852 281724 389904
rect 281776 389892 281782 389904
rect 342438 389892 342444 389904
rect 281776 389864 342444 389892
rect 281776 389852 281782 389864
rect 342438 389852 342444 389864
rect 342496 389852 342502 389904
rect 345750 389852 345756 389904
rect 345808 389892 345814 389904
rect 366174 389892 366180 389904
rect 345808 389864 366180 389892
rect 345808 389852 345814 389864
rect 366174 389852 366180 389864
rect 366232 389852 366238 389904
rect 265986 389784 265992 389836
rect 266044 389824 266050 389836
rect 350534 389824 350540 389836
rect 266044 389796 350540 389824
rect 266044 389784 266050 389796
rect 350534 389784 350540 389796
rect 350592 389784 350598 389836
rect 354122 389784 354128 389836
rect 354180 389824 354186 389836
rect 380986 389824 380992 389836
rect 354180 389796 380992 389824
rect 354180 389784 354186 389796
rect 380986 389784 380992 389796
rect 381044 389784 381050 389836
rect 377950 389716 377956 389768
rect 378008 389756 378014 389768
rect 378134 389756 378140 389768
rect 378008 389728 378140 389756
rect 378008 389716 378014 389728
rect 378134 389716 378140 389728
rect 378192 389716 378198 389768
rect 377674 389648 377680 389700
rect 377732 389688 377738 389700
rect 378042 389688 378048 389700
rect 377732 389660 378048 389688
rect 377732 389648 377738 389660
rect 378042 389648 378048 389660
rect 378100 389648 378106 389700
rect 340138 389104 340144 389156
rect 340196 389144 340202 389156
rect 346762 389144 346768 389156
rect 340196 389116 346768 389144
rect 340196 389104 340202 389116
rect 346762 389104 346768 389116
rect 346820 389104 346826 389156
rect 327994 388968 328000 389020
rect 328052 389008 328058 389020
rect 349706 389008 349712 389020
rect 328052 388980 349712 389008
rect 328052 388968 328058 388980
rect 349706 388968 349712 388980
rect 349764 388968 349770 389020
rect 344922 388900 344928 388952
rect 344980 388940 344986 388952
rect 370130 388940 370136 388952
rect 344980 388912 370136 388940
rect 344980 388900 344986 388912
rect 370130 388900 370136 388912
rect 370188 388900 370194 388952
rect 335262 388832 335268 388884
rect 335320 388872 335326 388884
rect 370222 388872 370228 388884
rect 335320 388844 370228 388872
rect 335320 388832 335326 388844
rect 370222 388832 370228 388844
rect 370280 388832 370286 388884
rect 324590 388764 324596 388816
rect 324648 388804 324654 388816
rect 384850 388804 384856 388816
rect 324648 388776 384856 388804
rect 324648 388764 324654 388776
rect 384850 388764 384856 388776
rect 384908 388764 384914 388816
rect 279602 388696 279608 388748
rect 279660 388736 279666 388748
rect 342530 388736 342536 388748
rect 279660 388708 342536 388736
rect 279660 388696 279666 388708
rect 342530 388696 342536 388708
rect 342588 388696 342594 388748
rect 343082 388696 343088 388748
rect 343140 388736 343146 388748
rect 370038 388736 370044 388748
rect 343140 388708 370044 388736
rect 343140 388696 343146 388708
rect 370038 388696 370044 388708
rect 370096 388696 370102 388748
rect 271506 388628 271512 388680
rect 271564 388668 271570 388680
rect 345290 388668 345296 388680
rect 271564 388640 345296 388668
rect 271564 388628 271570 388640
rect 345290 388628 345296 388640
rect 345348 388628 345354 388680
rect 347406 388628 347412 388680
rect 347464 388668 347470 388680
rect 360562 388668 360568 388680
rect 347464 388640 360568 388668
rect 347464 388628 347470 388640
rect 360562 388628 360568 388640
rect 360620 388628 360626 388680
rect 261938 388560 261944 388612
rect 261996 388600 262002 388612
rect 342254 388600 342260 388612
rect 261996 388572 342260 388600
rect 261996 388560 262002 388572
rect 342254 388560 342260 388572
rect 342312 388560 342318 388612
rect 347130 388560 347136 388612
rect 347188 388600 347194 388612
rect 375374 388600 375380 388612
rect 347188 388572 375380 388600
rect 347188 388560 347194 388572
rect 375374 388560 375380 388572
rect 375432 388560 375438 388612
rect 267642 388492 267648 388544
rect 267700 388532 267706 388544
rect 349338 388532 349344 388544
rect 267700 388504 349344 388532
rect 267700 388492 267706 388504
rect 349338 388492 349344 388504
rect 349396 388492 349402 388544
rect 263410 388424 263416 388476
rect 263468 388464 263474 388476
rect 347866 388464 347872 388476
rect 263468 388436 347872 388464
rect 263468 388424 263474 388436
rect 347866 388424 347872 388436
rect 347924 388424 347930 388476
rect 351362 388424 351368 388476
rect 351420 388464 351426 388476
rect 361206 388464 361212 388476
rect 351420 388436 361212 388464
rect 351420 388424 351426 388436
rect 361206 388424 361212 388436
rect 361264 388424 361270 388476
rect 351270 388152 351276 388204
rect 351328 388192 351334 388204
rect 355042 388192 355048 388204
rect 351328 388164 355048 388192
rect 351328 388152 351334 388164
rect 355042 388152 355048 388164
rect 355100 388152 355106 388204
rect 357618 387472 357624 387524
rect 357676 387512 357682 387524
rect 358538 387512 358544 387524
rect 357676 387484 358544 387512
rect 357676 387472 357682 387484
rect 358538 387472 358544 387484
rect 358596 387472 358602 387524
rect 263318 387336 263324 387388
rect 263376 387376 263382 387388
rect 344830 387376 344836 387388
rect 263376 387348 344836 387376
rect 263376 387336 263382 387348
rect 344830 387336 344836 387348
rect 344888 387336 344894 387388
rect 347314 387336 347320 387388
rect 347372 387376 347378 387388
rect 354950 387376 354956 387388
rect 347372 387348 354956 387376
rect 347372 387336 347378 387348
rect 354950 387336 354956 387348
rect 355008 387336 355014 387388
rect 330846 387268 330852 387320
rect 330904 387308 330910 387320
rect 380250 387308 380256 387320
rect 330904 387280 380256 387308
rect 330904 387268 330910 387280
rect 380250 387268 380256 387280
rect 380308 387268 380314 387320
rect 278406 387200 278412 387252
rect 278464 387240 278470 387252
rect 345198 387240 345204 387252
rect 278464 387212 345204 387240
rect 278464 387200 278470 387212
rect 345198 387200 345204 387212
rect 345256 387200 345262 387252
rect 346026 387200 346032 387252
rect 346084 387240 346090 387252
rect 379882 387240 379888 387252
rect 346084 387212 379888 387240
rect 346084 387200 346090 387212
rect 379882 387200 379888 387212
rect 379940 387200 379946 387252
rect 344094 387132 344100 387184
rect 344152 387172 344158 387184
rect 382274 387172 382280 387184
rect 344152 387144 382280 387172
rect 344152 387132 344158 387144
rect 382274 387132 382280 387144
rect 382332 387132 382338 387184
rect 264882 387064 264888 387116
rect 264940 387104 264946 387116
rect 346394 387104 346400 387116
rect 264940 387076 346400 387104
rect 264940 387064 264946 387076
rect 346394 387064 346400 387076
rect 346452 387064 346458 387116
rect 349798 387064 349804 387116
rect 349856 387104 349862 387116
rect 357710 387104 357716 387116
rect 349856 387076 357716 387104
rect 349856 387064 349862 387076
rect 357710 387064 357716 387076
rect 357768 387064 357774 387116
rect 350074 386520 350080 386572
rect 350132 386560 350138 386572
rect 355686 386560 355692 386572
rect 350132 386532 355692 386560
rect 350132 386520 350138 386532
rect 355686 386520 355692 386532
rect 355744 386520 355750 386572
rect 320174 386316 320180 386368
rect 320232 386356 320238 386368
rect 321002 386356 321008 386368
rect 320232 386328 321008 386356
rect 320232 386316 320238 386328
rect 321002 386316 321008 386328
rect 321060 386316 321066 386368
rect 322934 386316 322940 386368
rect 322992 386356 322998 386368
rect 323762 386356 323768 386368
rect 322992 386328 323768 386356
rect 322992 386316 322998 386328
rect 323762 386316 323768 386328
rect 323820 386316 323826 386368
rect 330662 386112 330668 386164
rect 330720 386152 330726 386164
rect 374730 386152 374736 386164
rect 330720 386124 374736 386152
rect 330720 386112 330726 386124
rect 374730 386112 374736 386124
rect 374788 386112 374794 386164
rect 329466 386044 329472 386096
rect 329524 386084 329530 386096
rect 377950 386084 377956 386096
rect 329524 386056 377956 386084
rect 329524 386044 329530 386056
rect 377950 386044 377956 386056
rect 378008 386044 378014 386096
rect 333698 385976 333704 386028
rect 333756 386016 333762 386028
rect 385954 386016 385960 386028
rect 333756 385988 385960 386016
rect 333756 385976 333762 385988
rect 385954 385976 385960 385988
rect 386012 385976 386018 386028
rect 282730 385908 282736 385960
rect 282788 385948 282794 385960
rect 339954 385948 339960 385960
rect 282788 385920 339960 385948
rect 282788 385908 282794 385920
rect 339954 385908 339960 385920
rect 340012 385908 340018 385960
rect 265894 385840 265900 385892
rect 265952 385880 265958 385892
rect 346670 385880 346676 385892
rect 265952 385852 346676 385880
rect 265952 385840 265958 385852
rect 346670 385840 346676 385852
rect 346728 385840 346734 385892
rect 276658 385772 276664 385824
rect 276716 385812 276722 385824
rect 363506 385812 363512 385824
rect 276716 385784 363512 385812
rect 276716 385772 276722 385784
rect 363506 385772 363512 385784
rect 363564 385772 363570 385824
rect 280890 385704 280896 385756
rect 280948 385744 280954 385756
rect 369762 385744 369768 385756
rect 280948 385716 369768 385744
rect 280948 385704 280954 385716
rect 369762 385704 369768 385716
rect 369820 385704 369826 385756
rect 273806 385636 273812 385688
rect 273864 385676 273870 385688
rect 365898 385676 365904 385688
rect 273864 385648 365904 385676
rect 273864 385636 273870 385648
rect 365898 385636 365904 385648
rect 365956 385636 365962 385688
rect 271138 385160 271144 385212
rect 271196 385200 271202 385212
rect 320174 385200 320180 385212
rect 271196 385172 320180 385200
rect 271196 385160 271202 385172
rect 320174 385160 320180 385172
rect 320232 385160 320238 385212
rect 262950 385092 262956 385144
rect 263008 385132 263014 385144
rect 322934 385132 322940 385144
rect 263008 385104 322940 385132
rect 263008 385092 263014 385104
rect 322934 385092 322940 385104
rect 322992 385092 322998 385144
rect 264330 385024 264336 385076
rect 264388 385064 264394 385076
rect 324590 385064 324596 385076
rect 264388 385036 324596 385064
rect 264388 385024 264394 385036
rect 324590 385024 324596 385036
rect 324648 385024 324654 385076
rect 319070 384956 319076 385008
rect 319128 384996 319134 385008
rect 319714 384996 319720 385008
rect 319128 384968 319720 384996
rect 319128 384956 319134 384968
rect 319714 384956 319720 384968
rect 319772 384956 319778 385008
rect 321738 384956 321744 385008
rect 321796 384996 321802 385008
rect 322382 384996 322388 385008
rect 321796 384968 322388 384996
rect 321796 384956 321802 384968
rect 322382 384956 322388 384968
rect 322440 384956 322446 385008
rect 259178 384276 259184 384328
rect 259236 384316 259242 384328
rect 348234 384316 348240 384328
rect 259236 384288 348240 384316
rect 259236 384276 259242 384288
rect 348234 384276 348240 384288
rect 348292 384276 348298 384328
rect 265618 383800 265624 383852
rect 265676 383840 265682 383852
rect 324314 383840 324320 383852
rect 265676 383812 324320 383840
rect 265676 383800 265682 383812
rect 324314 383800 324320 383812
rect 324372 383800 324378 383852
rect 261478 383732 261484 383784
rect 261536 383772 261542 383784
rect 321738 383772 321744 383784
rect 261536 383744 321744 383772
rect 261536 383732 261542 383744
rect 321738 383732 321744 383744
rect 321796 383732 321802 383784
rect 258718 383664 258724 383716
rect 258776 383704 258782 383716
rect 319070 383704 319076 383716
rect 258776 383676 319076 383704
rect 258776 383664 258782 383676
rect 319070 383664 319076 383676
rect 319128 383664 319134 383716
rect 343542 383460 343548 383512
rect 343600 383500 343606 383512
rect 359090 383500 359096 383512
rect 343600 383472 359096 383500
rect 343600 383460 343606 383472
rect 359090 383460 359096 383472
rect 359148 383460 359154 383512
rect 343450 383392 343456 383444
rect 343508 383432 343514 383444
rect 367738 383432 367744 383444
rect 343508 383404 367744 383432
rect 343508 383392 343514 383404
rect 367738 383392 367744 383404
rect 367796 383392 367802 383444
rect 331030 383324 331036 383376
rect 331088 383364 331094 383376
rect 379790 383364 379796 383376
rect 331088 383336 379796 383364
rect 331088 383324 331094 383336
rect 379790 383324 379796 383336
rect 379848 383324 379854 383376
rect 332410 383256 332416 383308
rect 332468 383296 332474 383308
rect 382550 383296 382556 383308
rect 332468 383268 382556 383296
rect 332468 383256 332474 383268
rect 382550 383256 382556 383268
rect 382608 383256 382614 383308
rect 274082 383188 274088 383240
rect 274140 383228 274146 383240
rect 348602 383228 348608 383240
rect 274140 383200 348608 383228
rect 274140 383188 274146 383200
rect 348602 383188 348608 383200
rect 348660 383188 348666 383240
rect 349890 383188 349896 383240
rect 349948 383228 349954 383240
rect 361850 383228 361856 383240
rect 349948 383200 361856 383228
rect 349948 383188 349954 383200
rect 361850 383188 361856 383200
rect 361908 383188 361914 383240
rect 277762 383120 277768 383172
rect 277820 383160 277826 383172
rect 360470 383160 360476 383172
rect 277820 383132 360476 383160
rect 277820 383120 277826 383132
rect 360470 383120 360476 383132
rect 360528 383120 360534 383172
rect 269942 383052 269948 383104
rect 270000 383092 270006 383104
rect 354490 383092 354496 383104
rect 270000 383064 354496 383092
rect 270000 383052 270006 383064
rect 354490 383052 354496 383064
rect 354548 383052 354554 383104
rect 263226 382984 263232 383036
rect 263284 383024 263290 383036
rect 348142 383024 348148 383036
rect 263284 382996 348148 383024
rect 263284 382984 263290 382996
rect 348142 382984 348148 382996
rect 348200 382984 348206 383036
rect 348602 382984 348608 383036
rect 348660 383024 348666 383036
rect 360194 383024 360200 383036
rect 348660 382996 360200 383024
rect 348660 382984 348666 382996
rect 360194 382984 360200 382996
rect 360252 382984 360258 383036
rect 280798 382916 280804 382968
rect 280856 382956 280862 382968
rect 372982 382956 372988 382968
rect 280856 382928 372988 382956
rect 280856 382916 280862 382928
rect 372982 382916 372988 382928
rect 373040 382916 373046 382968
rect 321646 382644 321652 382696
rect 321704 382684 321710 382696
rect 322474 382684 322480 382696
rect 321704 382656 322480 382684
rect 321704 382644 321710 382656
rect 322474 382644 322480 382656
rect 322532 382644 322538 382696
rect 321646 382480 321652 382492
rect 316006 382452 321652 382480
rect 271230 382372 271236 382424
rect 271288 382412 271294 382424
rect 316006 382412 316034 382452
rect 321646 382440 321652 382452
rect 321704 382440 321710 382492
rect 271288 382384 316034 382412
rect 271288 382372 271294 382384
rect 318886 382372 318892 382424
rect 318944 382412 318950 382424
rect 319622 382412 319628 382424
rect 318944 382384 319628 382412
rect 318944 382372 318950 382384
rect 319622 382372 319628 382384
rect 319680 382372 319686 382424
rect 260098 382304 260104 382356
rect 260156 382344 260162 382356
rect 260156 382316 319024 382344
rect 260156 382304 260162 382316
rect 318996 382288 319024 382316
rect 257338 382236 257344 382288
rect 257396 382276 257402 382288
rect 318886 382276 318892 382288
rect 257396 382248 318892 382276
rect 257396 382236 257402 382248
rect 318886 382236 318892 382248
rect 318944 382236 318950 382288
rect 318978 382236 318984 382288
rect 319036 382276 319042 382288
rect 319438 382276 319444 382288
rect 319036 382248 319444 382276
rect 319036 382236 319042 382248
rect 319438 382236 319444 382248
rect 319496 382236 319502 382288
rect 323026 381692 323032 381744
rect 323084 381732 323090 381744
rect 323670 381732 323676 381744
rect 323084 381704 323676 381732
rect 323084 381692 323090 381704
rect 323670 381692 323676 381704
rect 323728 381692 323734 381744
rect 320266 381284 320272 381336
rect 320324 381324 320330 381336
rect 320818 381324 320824 381336
rect 320324 381296 320824 381324
rect 320324 381284 320330 381296
rect 320818 381284 320824 381296
rect 320876 381284 320882 381336
rect 272610 381012 272616 381064
rect 272668 381052 272674 381064
rect 320266 381052 320272 381064
rect 272668 381024 320272 381052
rect 272668 381012 272674 381024
rect 320266 381012 320272 381024
rect 320324 381012 320330 381064
rect 253842 380944 253848 380996
rect 253900 380984 253906 380996
rect 313366 380984 313372 380996
rect 253900 380956 313372 380984
rect 253900 380944 253906 380956
rect 313366 380944 313372 380956
rect 313424 380944 313430 380996
rect 262858 380876 262864 380928
rect 262916 380916 262922 380928
rect 323026 380916 323032 380928
rect 262916 380888 323032 380916
rect 262916 380876 262922 380888
rect 323026 380876 323032 380888
rect 323084 380876 323090 380928
rect 314838 380332 314844 380384
rect 314896 380372 314902 380384
rect 315298 380372 315304 380384
rect 314896 380344 315304 380372
rect 314896 380332 314902 380344
rect 315298 380332 315304 380344
rect 315356 380332 315362 380384
rect 281810 380196 281816 380248
rect 281868 380236 281874 380248
rect 342714 380236 342720 380248
rect 281868 380208 342720 380236
rect 281868 380196 281874 380208
rect 342714 380196 342720 380208
rect 342772 380196 342778 380248
rect 261846 380128 261852 380180
rect 261904 380168 261910 380180
rect 348050 380168 348056 380180
rect 261904 380140 348056 380168
rect 261904 380128 261910 380140
rect 348050 380128 348056 380140
rect 348108 380128 348114 380180
rect 272702 379856 272708 379908
rect 272760 379896 272766 379908
rect 314838 379896 314844 379908
rect 272760 379868 314844 379896
rect 272760 379856 272766 379868
rect 314838 379856 314844 379868
rect 314896 379856 314902 379908
rect 244918 379788 244924 379840
rect 244976 379828 244982 379840
rect 303614 379828 303620 379840
rect 244976 379800 303620 379828
rect 244976 379788 244982 379800
rect 303614 379788 303620 379800
rect 303672 379828 303678 379840
rect 304258 379828 304264 379840
rect 303672 379800 304264 379828
rect 303672 379788 303678 379800
rect 304258 379788 304264 379800
rect 304316 379788 304322 379840
rect 249058 379720 249064 379772
rect 249116 379760 249122 379772
rect 309134 379760 309140 379772
rect 249116 379732 309140 379760
rect 249116 379720 249122 379732
rect 309134 379720 309140 379732
rect 309192 379720 309198 379772
rect 264698 379652 264704 379704
rect 264756 379692 264762 379704
rect 264756 379664 324544 379692
rect 264756 379652 264762 379664
rect 324516 379636 324544 379664
rect 264422 379584 264428 379636
rect 264480 379624 264486 379636
rect 264480 379596 324360 379624
rect 264480 379584 264486 379596
rect 324332 379568 324360 379596
rect 324498 379584 324504 379636
rect 324556 379624 324562 379636
rect 325142 379624 325148 379636
rect 324556 379596 325148 379624
rect 324556 379584 324562 379596
rect 325142 379584 325148 379596
rect 325200 379584 325206 379636
rect 259362 379516 259368 379568
rect 259420 379556 259426 379568
rect 320910 379556 320916 379568
rect 259420 379528 320916 379556
rect 259420 379516 259426 379528
rect 320910 379516 320916 379528
rect 320968 379516 320974 379568
rect 324314 379516 324320 379568
rect 324372 379556 324378 379568
rect 325050 379556 325056 379568
rect 324372 379528 325056 379556
rect 324372 379516 324378 379528
rect 325050 379516 325056 379528
rect 325108 379516 325114 379568
rect 345842 379516 345848 379568
rect 345900 379556 345906 379568
rect 353570 379556 353576 379568
rect 345900 379528 353576 379556
rect 345900 379516 345906 379528
rect 353570 379516 353576 379528
rect 353628 379516 353634 379568
rect 313918 378468 313924 378480
rect 311866 378440 313924 378468
rect 254118 378292 254124 378344
rect 254176 378332 254182 378344
rect 311866 378332 311894 378440
rect 313918 378428 313924 378440
rect 313976 378428 313982 378480
rect 319530 378400 319536 378412
rect 254176 378304 311894 378332
rect 313844 378372 319536 378400
rect 254176 378292 254182 378304
rect 259730 378224 259736 378276
rect 259788 378264 259794 378276
rect 313844 378264 313872 378372
rect 319530 378360 319536 378372
rect 319588 378360 319594 378412
rect 259788 378236 313872 378264
rect 259788 378224 259794 378236
rect 313918 378224 313924 378276
rect 313976 378264 313982 378276
rect 314194 378264 314200 378276
rect 313976 378236 314200 378264
rect 313976 378224 313982 378236
rect 314194 378224 314200 378236
rect 314252 378224 314258 378276
rect 263502 378156 263508 378208
rect 263560 378196 263566 378208
rect 323854 378196 323860 378208
rect 263560 378168 323860 378196
rect 263560 378156 263566 378168
rect 323854 378156 323860 378168
rect 323912 378156 323918 378208
rect 348694 378020 348700 378072
rect 348752 378060 348758 378072
rect 357250 378060 357256 378072
rect 348752 378032 357256 378060
rect 348752 378020 348758 378032
rect 357250 378020 357256 378032
rect 357308 378020 357314 378072
rect 348786 377544 348792 377596
rect 348844 377584 348850 377596
rect 358998 377584 359004 377596
rect 348844 377556 359004 377584
rect 348844 377544 348850 377556
rect 358998 377544 359004 377556
rect 359056 377544 359062 377596
rect 350166 377476 350172 377528
rect 350224 377516 350230 377528
rect 363230 377516 363236 377528
rect 350224 377488 363236 377516
rect 350224 377476 350230 377488
rect 363230 377476 363236 377488
rect 363288 377476 363294 377528
rect 281902 377408 281908 377460
rect 281960 377448 281966 377460
rect 342622 377448 342628 377460
rect 281960 377420 342628 377448
rect 281960 377408 281966 377420
rect 342622 377408 342628 377420
rect 342680 377408 342686 377460
rect 348510 377408 348516 377460
rect 348568 377448 348574 377460
rect 367370 377448 367376 377460
rect 348568 377420 367376 377448
rect 348568 377408 348574 377420
rect 367370 377408 367376 377420
rect 367428 377408 367434 377460
rect 264238 376932 264244 376984
rect 264296 376972 264302 376984
rect 311986 376972 311992 376984
rect 264296 376944 311992 376972
rect 264296 376932 264302 376944
rect 311986 376932 311992 376944
rect 312044 376972 312050 376984
rect 312538 376972 312544 376984
rect 312044 376944 312544 376972
rect 312044 376932 312050 376944
rect 312538 376932 312544 376944
rect 312596 376932 312602 376984
rect 242158 376864 242164 376916
rect 242216 376904 242222 376916
rect 301590 376904 301596 376916
rect 242216 376876 301596 376904
rect 242216 376864 242222 376876
rect 301590 376864 301596 376876
rect 301648 376864 301654 376916
rect 255498 376796 255504 376848
rect 255556 376836 255562 376848
rect 316126 376836 316132 376848
rect 255556 376808 316132 376836
rect 255556 376796 255562 376808
rect 316126 376796 316132 376808
rect 316184 376796 316190 376848
rect 245010 376728 245016 376780
rect 245068 376768 245074 376780
rect 307846 376768 307852 376780
rect 245068 376740 307852 376768
rect 245068 376728 245074 376740
rect 307846 376728 307852 376740
rect 307904 376728 307910 376780
rect 291286 376116 291292 376168
rect 291344 376156 291350 376168
rect 291930 376156 291936 376168
rect 291344 376128 291936 376156
rect 291344 376116 291350 376128
rect 291930 376116 291936 376128
rect 291988 376156 291994 376168
rect 292298 376156 292304 376168
rect 291988 376128 292304 376156
rect 291988 376116 291994 376128
rect 292298 376116 292304 376128
rect 292356 376116 292362 376168
rect 275370 376048 275376 376100
rect 275428 376088 275434 376100
rect 293034 376088 293040 376100
rect 275428 376060 293040 376088
rect 275428 376048 275434 376060
rect 293034 376048 293040 376060
rect 293092 376048 293098 376100
rect 274174 375980 274180 376032
rect 274232 376020 274238 376032
rect 292206 376020 292212 376032
rect 274232 375992 292212 376020
rect 274232 375980 274238 375992
rect 292206 375980 292212 375992
rect 292264 375980 292270 376032
rect 275646 375912 275652 375964
rect 275704 375952 275710 375964
rect 298554 375952 298560 375964
rect 275704 375924 298560 375952
rect 275704 375912 275710 375924
rect 298554 375912 298560 375924
rect 298612 375912 298618 375964
rect 274266 375844 274272 375896
rect 274324 375884 274330 375896
rect 302602 375884 302608 375896
rect 274324 375856 302608 375884
rect 274324 375844 274330 375856
rect 302602 375844 302608 375856
rect 302660 375844 302666 375896
rect 279694 375776 279700 375828
rect 279752 375816 279758 375828
rect 312906 375816 312912 375828
rect 279752 375788 312912 375816
rect 279752 375776 279758 375788
rect 312906 375776 312912 375788
rect 312964 375776 312970 375828
rect 264514 375708 264520 375760
rect 264572 375748 264578 375760
rect 300210 375748 300216 375760
rect 264572 375720 300216 375748
rect 264572 375708 264578 375720
rect 300210 375708 300216 375720
rect 300268 375708 300274 375760
rect 267090 375640 267096 375692
rect 267148 375680 267154 375692
rect 311066 375680 311072 375692
rect 267148 375652 311072 375680
rect 267148 375640 267154 375652
rect 311066 375640 311072 375652
rect 311124 375640 311130 375692
rect 232498 375572 232504 375624
rect 232556 375612 232562 375624
rect 291286 375612 291292 375624
rect 232556 375584 291292 375612
rect 232556 375572 232562 375584
rect 291286 375572 291292 375584
rect 291344 375572 291350 375624
rect 298554 375572 298560 375624
rect 298612 375612 298618 375624
rect 298922 375612 298928 375624
rect 298612 375584 298928 375612
rect 298612 375572 298618 375584
rect 298922 375572 298928 375584
rect 298980 375572 298986 375624
rect 236638 375504 236644 375556
rect 236696 375544 236702 375556
rect 297450 375544 297456 375556
rect 236696 375516 297456 375544
rect 236696 375504 236702 375516
rect 297450 375504 297456 375516
rect 297508 375544 297514 375556
rect 301498 375544 301504 375556
rect 297508 375516 301504 375544
rect 297508 375504 297514 375516
rect 301498 375504 301504 375516
rect 301556 375504 301562 375556
rect 238662 375436 238668 375488
rect 238720 375476 238726 375488
rect 298830 375476 298836 375488
rect 238720 375448 298836 375476
rect 238720 375436 238726 375448
rect 298830 375436 298836 375448
rect 298888 375436 298894 375488
rect 261294 375368 261300 375420
rect 261352 375408 261358 375420
rect 321830 375408 321836 375420
rect 261352 375380 321836 375408
rect 261352 375368 261358 375380
rect 321830 375368 321836 375380
rect 321888 375408 321894 375420
rect 322290 375408 322296 375420
rect 321888 375380 322296 375408
rect 321888 375368 321894 375380
rect 322290 375368 322296 375380
rect 322348 375368 322354 375420
rect 268378 374756 268384 374808
rect 268436 374796 268442 374808
rect 293310 374796 293316 374808
rect 268436 374768 293316 374796
rect 268436 374756 268442 374768
rect 293310 374756 293316 374768
rect 293368 374756 293374 374808
rect 294322 374756 294328 374808
rect 294380 374796 294386 374808
rect 294782 374796 294788 374808
rect 294380 374768 294788 374796
rect 294380 374756 294386 374768
rect 294782 374756 294788 374768
rect 294840 374756 294846 374808
rect 318426 374756 318432 374808
rect 318484 374796 318490 374808
rect 318484 374768 321554 374796
rect 318484 374756 318490 374768
rect 267182 374688 267188 374740
rect 267240 374728 267246 374740
rect 275278 374728 275284 374740
rect 267240 374700 275284 374728
rect 267240 374688 267246 374700
rect 275278 374688 275284 374700
rect 275336 374728 275342 374740
rect 306190 374728 306196 374740
rect 275336 374700 306196 374728
rect 275336 374688 275342 374700
rect 306190 374688 306196 374700
rect 306248 374688 306254 374740
rect 318886 374688 318892 374740
rect 318944 374728 318950 374740
rect 319162 374728 319168 374740
rect 318944 374700 319168 374728
rect 318944 374688 318950 374700
rect 319162 374688 319168 374700
rect 319220 374688 319226 374740
rect 320174 374688 320180 374740
rect 320232 374728 320238 374740
rect 321002 374728 321008 374740
rect 320232 374700 321008 374728
rect 320232 374688 320238 374700
rect 321002 374688 321008 374700
rect 321060 374688 321066 374740
rect 321526 374728 321554 374768
rect 324314 374756 324320 374808
rect 324372 374796 324378 374808
rect 324958 374796 324964 374808
rect 324372 374768 324964 374796
rect 324372 374756 324378 374768
rect 324958 374756 324964 374768
rect 325016 374756 325022 374808
rect 332042 374728 332048 374740
rect 321526 374700 332048 374728
rect 332042 374688 332048 374700
rect 332100 374688 332106 374740
rect 219250 374620 219256 374672
rect 219308 374660 219314 374672
rect 282822 374660 282828 374672
rect 219308 374632 282828 374660
rect 219308 374620 219314 374632
rect 282822 374620 282828 374632
rect 282880 374620 282886 374672
rect 299382 374620 299388 374672
rect 299440 374660 299446 374672
rect 340782 374660 340788 374672
rect 299440 374632 340788 374660
rect 299440 374620 299446 374632
rect 340782 374620 340788 374632
rect 340840 374620 340846 374672
rect 267274 374552 267280 374604
rect 267332 374592 267338 374604
rect 295794 374592 295800 374604
rect 267332 374564 295800 374592
rect 267332 374552 267338 374564
rect 295794 374552 295800 374564
rect 295852 374552 295858 374604
rect 321646 374552 321652 374604
rect 321704 374592 321710 374604
rect 322382 374592 322388 374604
rect 321704 374564 322388 374592
rect 321704 374552 321710 374564
rect 322382 374552 322388 374564
rect 322440 374552 322446 374604
rect 324498 374552 324504 374604
rect 324556 374592 324562 374604
rect 324682 374592 324688 374604
rect 324556 374564 324688 374592
rect 324556 374552 324562 374564
rect 324682 374552 324688 374564
rect 324740 374552 324746 374604
rect 277302 374484 277308 374536
rect 277360 374524 277366 374536
rect 308398 374524 308404 374536
rect 277360 374496 308404 374524
rect 277360 374484 277366 374496
rect 308398 374484 308404 374496
rect 308456 374484 308462 374536
rect 324406 374484 324412 374536
rect 324464 374524 324470 374536
rect 325326 374524 325332 374536
rect 324464 374496 325332 374524
rect 324464 374484 324470 374496
rect 325326 374484 325332 374496
rect 325384 374484 325390 374536
rect 272334 374416 272340 374468
rect 272392 374456 272398 374468
rect 303246 374456 303252 374468
rect 272392 374428 303252 374456
rect 272392 374416 272398 374428
rect 303246 374416 303252 374428
rect 303304 374416 303310 374468
rect 273070 374348 273076 374400
rect 273128 374388 273134 374400
rect 304350 374388 304356 374400
rect 273128 374360 304356 374388
rect 273128 374348 273134 374360
rect 304350 374348 304356 374360
rect 304408 374348 304414 374400
rect 269758 374280 269764 374332
rect 269816 374320 269822 374332
rect 305362 374320 305368 374332
rect 269816 374292 305368 374320
rect 269816 374280 269822 374292
rect 305362 374280 305368 374292
rect 305420 374280 305426 374332
rect 277854 374212 277860 374264
rect 277912 374252 277918 374264
rect 317966 374252 317972 374264
rect 277912 374224 317972 374252
rect 277912 374212 277918 374224
rect 317966 374212 317972 374224
rect 318024 374252 318030 374264
rect 318426 374252 318432 374264
rect 318024 374224 318432 374252
rect 318024 374212 318030 374224
rect 318426 374212 318432 374224
rect 318484 374212 318490 374264
rect 245102 374144 245108 374196
rect 245160 374184 245166 374196
rect 297082 374184 297088 374196
rect 245160 374156 297088 374184
rect 245160 374144 245166 374156
rect 297082 374144 297088 374156
rect 297140 374144 297146 374196
rect 238846 374076 238852 374128
rect 238904 374116 238910 374128
rect 298830 374116 298836 374128
rect 238904 374088 298836 374116
rect 238904 374076 238910 374088
rect 298830 374076 298836 374088
rect 298888 374076 298894 374128
rect 219342 374008 219348 374060
rect 219400 374048 219406 374060
rect 294322 374048 294328 374060
rect 219400 374020 294328 374048
rect 219400 374008 219406 374020
rect 294322 374008 294328 374020
rect 294380 374008 294386 374060
rect 153194 373940 153200 373992
rect 153252 373980 153258 373992
rect 280154 373980 280160 373992
rect 153252 373952 280160 373980
rect 153252 373940 153258 373952
rect 280154 373940 280160 373952
rect 280212 373940 280218 373992
rect 220078 373872 220084 373924
rect 220136 373912 220142 373924
rect 282270 373912 282276 373924
rect 220136 373884 282276 373912
rect 220136 373872 220142 373884
rect 282270 373872 282276 373884
rect 282328 373872 282334 373924
rect 297358 373872 297364 373924
rect 297416 373912 297422 373924
rect 307110 373912 307116 373924
rect 297416 373884 307116 373912
rect 297416 373872 297422 373884
rect 307110 373872 307116 373884
rect 307168 373872 307174 373924
rect 314930 373600 314936 373652
rect 314988 373640 314994 373652
rect 315482 373640 315488 373652
rect 314988 373612 315488 373640
rect 314988 373600 314994 373612
rect 315482 373600 315488 373612
rect 315540 373600 315546 373652
rect 304166 373464 304172 373516
rect 304224 373504 304230 373516
rect 304350 373504 304356 373516
rect 304224 373476 304356 373504
rect 304224 373464 304230 373476
rect 304350 373464 304356 373476
rect 304408 373464 304414 373516
rect 300854 373396 300860 373448
rect 300912 373436 300918 373448
rect 338022 373436 338028 373448
rect 300912 373408 338028 373436
rect 300912 373396 300918 373408
rect 338022 373396 338028 373408
rect 338080 373396 338086 373448
rect 294506 373328 294512 373380
rect 294564 373368 294570 373380
rect 332226 373368 332232 373380
rect 294564 373340 332232 373368
rect 294564 373328 294570 373340
rect 332226 373328 332232 373340
rect 332284 373328 332290 373380
rect 220722 373260 220728 373312
rect 220780 373300 220786 373312
rect 281258 373300 281264 373312
rect 220780 373272 281264 373300
rect 220780 373260 220786 373272
rect 281258 373260 281264 373272
rect 281316 373300 281322 373312
rect 287422 373300 287428 373312
rect 281316 373272 287428 373300
rect 281316 373260 281322 373272
rect 287422 373260 287428 373272
rect 287480 373260 287486 373312
rect 296622 373260 296628 373312
rect 296680 373300 296686 373312
rect 340690 373300 340696 373312
rect 296680 373272 340696 373300
rect 296680 373260 296686 373272
rect 340690 373260 340696 373272
rect 340748 373260 340754 373312
rect 233878 373192 233884 373244
rect 233936 373232 233942 373244
rect 294506 373232 294512 373244
rect 233936 373204 294512 373232
rect 233936 373192 233942 373204
rect 294506 373192 294512 373204
rect 294564 373192 294570 373244
rect 278130 373124 278136 373176
rect 278188 373164 278194 373176
rect 294598 373164 294604 373176
rect 278188 373136 294604 373164
rect 278188 373124 278194 373136
rect 294598 373124 294604 373136
rect 294656 373164 294662 373176
rect 295334 373164 295340 373176
rect 294656 373136 295340 373164
rect 294656 373124 294662 373136
rect 295334 373124 295340 373136
rect 295392 373124 295398 373176
rect 275186 373056 275192 373108
rect 275244 373096 275250 373108
rect 297818 373096 297824 373108
rect 275244 373068 297824 373096
rect 275244 373056 275250 373068
rect 297818 373056 297824 373068
rect 297876 373096 297882 373108
rect 299382 373096 299388 373108
rect 297876 373068 299388 373096
rect 297876 373056 297882 373068
rect 299382 373056 299388 373068
rect 299440 373056 299446 373108
rect 279050 372988 279056 373040
rect 279108 373028 279114 373040
rect 299934 373028 299940 373040
rect 279108 373000 299940 373028
rect 279108 372988 279114 373000
rect 299934 372988 299940 373000
rect 299992 373028 299998 373040
rect 300302 373028 300308 373040
rect 299992 373000 300308 373028
rect 299992 372988 299998 373000
rect 300302 372988 300308 373000
rect 300360 372988 300366 373040
rect 313366 372988 313372 373040
rect 313424 373028 313430 373040
rect 314654 373028 314660 373040
rect 313424 373000 314660 373028
rect 313424 372988 313430 373000
rect 314654 372988 314660 373000
rect 314712 372988 314718 373040
rect 322842 372988 322848 373040
rect 322900 373028 322906 373040
rect 323026 373028 323032 373040
rect 322900 373000 323032 373028
rect 322900 372988 322906 373000
rect 323026 372988 323032 373000
rect 323084 372988 323090 373040
rect 275094 372920 275100 372972
rect 275152 372960 275158 372972
rect 298738 372960 298744 372972
rect 275152 372932 298744 372960
rect 275152 372920 275158 372932
rect 298738 372920 298744 372932
rect 298796 372920 298802 372972
rect 275738 372852 275744 372904
rect 275796 372892 275802 372904
rect 300854 372892 300860 372904
rect 275796 372864 300860 372892
rect 275796 372852 275802 372864
rect 300854 372852 300860 372864
rect 300912 372852 300918 372904
rect 277210 372784 277216 372836
rect 277268 372824 277274 372836
rect 303522 372824 303528 372836
rect 277268 372796 303528 372824
rect 277268 372784 277274 372796
rect 303522 372784 303528 372796
rect 303580 372784 303586 372836
rect 272426 372716 272432 372768
rect 272484 372756 272490 372768
rect 301038 372756 301044 372768
rect 272484 372728 301044 372756
rect 272484 372716 272490 372728
rect 301038 372716 301044 372728
rect 301096 372716 301102 372768
rect 274542 372648 274548 372700
rect 274600 372688 274606 372700
rect 274600 372660 302234 372688
rect 274600 372648 274606 372660
rect 278222 372580 278228 372632
rect 278280 372620 278286 372632
rect 296622 372620 296628 372632
rect 278280 372592 296628 372620
rect 278280 372580 278286 372592
rect 296622 372580 296628 372592
rect 296680 372580 296686 372632
rect 302206 372620 302234 372660
rect 302206 372592 304994 372620
rect 304966 372552 304994 372592
rect 307294 372552 307300 372564
rect 304966 372524 307300 372552
rect 307294 372512 307300 372524
rect 307352 372512 307358 372564
rect 314930 372512 314936 372564
rect 314988 372552 314994 372564
rect 358354 372552 358360 372564
rect 314988 372524 358360 372552
rect 314988 372512 314994 372524
rect 358354 372512 358360 372524
rect 358412 372512 358418 372564
rect 298830 372444 298836 372496
rect 298888 372484 298894 372496
rect 335078 372484 335084 372496
rect 298888 372456 335084 372484
rect 298888 372444 298894 372456
rect 335078 372444 335084 372456
rect 335136 372444 335142 372496
rect 303246 372376 303252 372428
rect 303304 372416 303310 372428
rect 337930 372416 337936 372428
rect 303304 372388 337936 372416
rect 303304 372376 303310 372388
rect 337930 372376 337936 372388
rect 337988 372376 337994 372428
rect 303522 372308 303528 372360
rect 303580 372348 303586 372360
rect 334618 372348 334624 372360
rect 303580 372320 334624 372348
rect 303580 372308 303586 372320
rect 334618 372308 334624 372320
rect 334676 372308 334682 372360
rect 278038 372240 278044 372292
rect 278096 372280 278102 372292
rect 288250 372280 288256 372292
rect 278096 372252 288256 372280
rect 278096 372240 278102 372252
rect 288250 372240 288256 372252
rect 288308 372240 288314 372292
rect 280154 372104 280160 372156
rect 280212 372144 280218 372156
rect 287698 372144 287704 372156
rect 280212 372116 287704 372144
rect 280212 372104 280218 372116
rect 287698 372104 287704 372116
rect 287756 372104 287762 372156
rect 288250 372104 288256 372156
rect 288308 372144 288314 372156
rect 288308 372116 292574 372144
rect 288308 372104 288314 372116
rect 273898 372036 273904 372088
rect 273956 372076 273962 372088
rect 282730 372076 282736 372088
rect 273956 372048 282736 372076
rect 273956 372036 273962 372048
rect 282730 372036 282736 372048
rect 282788 372036 282794 372088
rect 282914 372036 282920 372088
rect 282972 372076 282978 372088
rect 288526 372076 288532 372088
rect 282972 372048 288532 372076
rect 282972 372036 282978 372048
rect 288526 372036 288532 372048
rect 288584 372036 288590 372088
rect 292546 372076 292574 372116
rect 293862 372104 293868 372156
rect 293920 372144 293926 372156
rect 294782 372144 294788 372156
rect 293920 372116 294788 372144
rect 293920 372104 293926 372116
rect 294782 372104 294788 372116
rect 294840 372144 294846 372156
rect 329650 372144 329656 372156
rect 294840 372116 329656 372144
rect 294840 372104 294846 372116
rect 329650 372104 329656 372116
rect 329708 372104 329714 372156
rect 328362 372076 328368 372088
rect 292546 372048 328368 372076
rect 328362 372036 328368 372048
rect 328420 372036 328426 372088
rect 279878 371968 279884 372020
rect 279936 372008 279942 372020
rect 294782 372008 294788 372020
rect 279936 371980 294788 372008
rect 279936 371968 279942 371980
rect 294782 371968 294788 371980
rect 294840 371968 294846 372020
rect 229738 371900 229744 371952
rect 229796 371940 229802 371952
rect 281074 371940 281080 371952
rect 229796 371912 281080 371940
rect 229796 371900 229802 371912
rect 281074 371900 281080 371912
rect 281132 371940 281138 371952
rect 286318 371940 286324 371952
rect 281132 371912 286324 371940
rect 281132 371900 281138 371912
rect 286318 371900 286324 371912
rect 286376 371900 286382 371952
rect 220630 371832 220636 371884
rect 220688 371872 220694 371884
rect 281166 371872 281172 371884
rect 220688 371844 281172 371872
rect 220688 371832 220694 371844
rect 281166 371832 281172 371844
rect 281224 371832 281230 371884
rect 282730 371832 282736 371884
rect 282788 371872 282794 371884
rect 283650 371872 283656 371884
rect 282788 371844 283656 371872
rect 282788 371832 282794 371844
rect 283650 371832 283656 371844
rect 283708 371832 283714 371884
rect 287606 371832 287612 371884
rect 287664 371872 287670 371884
rect 293862 371872 293868 371884
rect 287664 371844 293868 371872
rect 287664 371832 287670 371844
rect 293862 371832 293868 371844
rect 293920 371832 293926 371884
rect 304074 371872 304080 371884
rect 299446 371844 304080 371872
rect 282270 371764 282276 371816
rect 282328 371804 282334 371816
rect 299446 371804 299474 371844
rect 304074 371832 304080 371844
rect 304132 371872 304138 371884
rect 322198 371872 322204 371884
rect 304132 371844 322204 371872
rect 304132 371832 304138 371844
rect 322198 371832 322204 371844
rect 322256 371832 322262 371884
rect 332778 371832 332784 371884
rect 332836 371872 332842 371884
rect 346210 371872 346216 371884
rect 332836 371844 346216 371872
rect 332836 371832 332842 371844
rect 346210 371832 346216 371844
rect 346268 371832 346274 371884
rect 282328 371776 299474 371804
rect 282328 371764 282334 371776
rect 282178 371696 282184 371748
rect 282236 371736 282242 371748
rect 305822 371736 305828 371748
rect 282236 371708 305828 371736
rect 282236 371696 282242 371708
rect 305822 371696 305828 371708
rect 305880 371696 305886 371748
rect 308306 371736 308312 371748
rect 306300 371708 308312 371736
rect 280706 371628 280712 371680
rect 280764 371668 280770 371680
rect 285214 371668 285220 371680
rect 280764 371640 285220 371668
rect 280764 371628 280770 371640
rect 285214 371628 285220 371640
rect 285272 371628 285278 371680
rect 287698 371628 287704 371680
rect 287756 371668 287762 371680
rect 306300 371668 306328 371708
rect 308306 371696 308312 371708
rect 308364 371696 308370 371748
rect 287756 371640 306328 371668
rect 287756 371628 287762 371640
rect 307754 371628 307760 371680
rect 307812 371668 307818 371680
rect 318058 371668 318064 371680
rect 307812 371640 318064 371668
rect 307812 371628 307818 371640
rect 318058 371628 318064 371640
rect 318116 371628 318122 371680
rect 281258 371560 281264 371612
rect 281316 371600 281322 371612
rect 312630 371600 312636 371612
rect 281316 371572 312636 371600
rect 281316 371560 281322 371572
rect 312630 371560 312636 371572
rect 312688 371600 312694 371612
rect 312814 371600 312820 371612
rect 312688 371572 312820 371600
rect 312688 371560 312694 371572
rect 312814 371560 312820 371572
rect 312872 371560 312878 371612
rect 316218 371560 316224 371612
rect 316276 371600 316282 371612
rect 316862 371600 316868 371612
rect 316276 371572 316868 371600
rect 316276 371560 316282 371572
rect 316862 371560 316868 371572
rect 316920 371560 316926 371612
rect 280614 371492 280620 371544
rect 280672 371532 280678 371544
rect 314010 371532 314016 371544
rect 280672 371504 314016 371532
rect 280672 371492 280678 371504
rect 314010 371492 314016 371504
rect 314068 371492 314074 371544
rect 277946 371424 277952 371476
rect 278004 371464 278010 371476
rect 279878 371464 279884 371476
rect 278004 371436 279884 371464
rect 278004 371424 278010 371436
rect 279878 371424 279884 371436
rect 279936 371424 279942 371476
rect 280706 371424 280712 371476
rect 280764 371464 280770 371476
rect 316236 371464 316264 371560
rect 332594 371492 332600 371544
rect 332652 371532 332658 371544
rect 333514 371532 333520 371544
rect 332652 371504 333520 371532
rect 332652 371492 332658 371504
rect 333514 371492 333520 371504
rect 333572 371492 333578 371544
rect 280764 371436 316264 371464
rect 280764 371424 280770 371436
rect 279234 371356 279240 371408
rect 279292 371396 279298 371408
rect 315758 371396 315764 371408
rect 279292 371368 315764 371396
rect 279292 371356 279298 371368
rect 315758 371356 315764 371368
rect 315816 371356 315822 371408
rect 320634 371356 320640 371408
rect 320692 371396 320698 371408
rect 332594 371396 332600 371408
rect 320692 371368 332600 371396
rect 320692 371356 320698 371368
rect 332594 371356 332600 371368
rect 332652 371356 332658 371408
rect 279510 371288 279516 371340
rect 279568 371328 279574 371340
rect 287606 371328 287612 371340
rect 279568 371300 287612 371328
rect 279568 371288 279574 371300
rect 287606 371288 287612 371300
rect 287664 371288 287670 371340
rect 288342 371288 288348 371340
rect 288400 371328 288406 371340
rect 291838 371328 291844 371340
rect 288400 371300 291844 371328
rect 288400 371288 288406 371300
rect 291838 371288 291844 371300
rect 291896 371288 291902 371340
rect 323578 371288 323584 371340
rect 323636 371328 323642 371340
rect 333974 371328 333980 371340
rect 323636 371300 333980 371328
rect 323636 371288 323642 371300
rect 333974 371288 333980 371300
rect 334032 371288 334038 371340
rect 3418 371220 3424 371272
rect 3476 371260 3482 371272
rect 257062 371260 257068 371272
rect 3476 371232 257068 371260
rect 3476 371220 3482 371232
rect 257062 371220 257068 371232
rect 257120 371260 257126 371272
rect 257120 371232 258074 371260
rect 257120 371220 257126 371232
rect 258046 371192 258074 371232
rect 279326 371220 279332 371272
rect 279384 371260 279390 371272
rect 287146 371260 287152 371272
rect 279384 371232 287152 371260
rect 279384 371220 279390 371232
rect 287146 371220 287152 371232
rect 287204 371220 287210 371272
rect 289722 371220 289728 371272
rect 289780 371260 289786 371272
rect 290734 371260 290740 371272
rect 289780 371232 290740 371260
rect 289780 371220 289786 371232
rect 290734 371220 290740 371232
rect 290792 371220 290798 371272
rect 326246 371220 326252 371272
rect 326304 371260 326310 371272
rect 332778 371260 332784 371272
rect 326304 371232 332784 371260
rect 326304 371220 326310 371232
rect 332778 371220 332784 371232
rect 332836 371220 332842 371272
rect 307754 371192 307760 371204
rect 258046 371164 307760 371192
rect 307754 371152 307760 371164
rect 307812 371152 307818 371204
rect 278590 371084 278596 371136
rect 278648 371124 278654 371136
rect 289722 371124 289728 371136
rect 278648 371096 289728 371124
rect 278648 371084 278654 371096
rect 289722 371084 289728 371096
rect 289780 371084 289786 371136
rect 278682 371056 278688 371068
rect 258046 371028 278688 371056
rect 233142 370676 233148 370728
rect 233200 370716 233206 370728
rect 258046 370716 258074 371028
rect 278682 371016 278688 371028
rect 278740 371056 278746 371068
rect 288342 371056 288348 371068
rect 278740 371028 288348 371056
rect 278740 371016 278746 371028
rect 288342 371016 288348 371028
rect 288400 371016 288406 371068
rect 300302 370880 300308 370932
rect 300360 370920 300366 370932
rect 327810 370920 327816 370932
rect 300360 370892 327816 370920
rect 300360 370880 300366 370892
rect 327810 370880 327816 370892
rect 327868 370880 327874 370932
rect 305086 370812 305092 370864
rect 305144 370852 305150 370864
rect 336458 370852 336464 370864
rect 305144 370824 336464 370852
rect 305144 370812 305150 370824
rect 336458 370812 336464 370824
rect 336516 370812 336522 370864
rect 271322 370744 271328 370796
rect 271380 370784 271386 370796
rect 305454 370784 305460 370796
rect 271380 370756 305460 370784
rect 271380 370744 271386 370756
rect 305454 370744 305460 370756
rect 305512 370744 305518 370796
rect 233200 370688 258074 370716
rect 233200 370676 233206 370688
rect 301498 370676 301504 370728
rect 301556 370716 301562 370728
rect 341518 370716 341524 370728
rect 301556 370688 341524 370716
rect 301556 370676 301562 370688
rect 341518 370676 341524 370688
rect 341576 370676 341582 370728
rect 231762 370608 231768 370660
rect 231820 370648 231826 370660
rect 278590 370648 278596 370660
rect 231820 370620 278596 370648
rect 231820 370608 231826 370620
rect 278590 370608 278596 370620
rect 278648 370608 278654 370660
rect 298094 370608 298100 370660
rect 298152 370648 298158 370660
rect 337838 370648 337844 370660
rect 298152 370620 337844 370648
rect 298152 370608 298158 370620
rect 337838 370608 337844 370620
rect 337896 370608 337902 370660
rect 245746 370540 245752 370592
rect 245804 370580 245810 370592
rect 271322 370580 271328 370592
rect 245804 370552 271328 370580
rect 245804 370540 245810 370552
rect 271322 370540 271328 370552
rect 271380 370540 271386 370592
rect 276566 370540 276572 370592
rect 276624 370580 276630 370592
rect 333790 370580 333796 370592
rect 276624 370552 333796 370580
rect 276624 370540 276630 370552
rect 333790 370540 333796 370552
rect 333848 370540 333854 370592
rect 258810 370472 258816 370524
rect 258868 370512 258874 370524
rect 318334 370512 318340 370524
rect 258868 370484 318340 370512
rect 258868 370472 258874 370484
rect 318334 370472 318340 370484
rect 318392 370472 318398 370524
rect 278314 370404 278320 370456
rect 278372 370444 278378 370456
rect 285122 370444 285128 370456
rect 278372 370416 285128 370444
rect 278372 370404 278378 370416
rect 285122 370404 285128 370416
rect 285180 370404 285186 370456
rect 235258 370336 235264 370388
rect 235316 370376 235322 370388
rect 295886 370376 295892 370388
rect 235316 370348 295892 370376
rect 235316 370336 235322 370348
rect 295886 370336 295892 370348
rect 295944 370336 295950 370388
rect 264606 370268 264612 370320
rect 264664 370308 264670 370320
rect 300302 370308 300308 370320
rect 264664 370280 300308 370308
rect 264664 370268 264670 370280
rect 300302 370268 300308 370280
rect 300360 370268 300366 370320
rect 279878 370200 279884 370252
rect 279936 370240 279942 370252
rect 306558 370240 306564 370252
rect 279936 370212 306564 370240
rect 279936 370200 279942 370212
rect 306558 370200 306564 370212
rect 306616 370200 306622 370252
rect 245194 370132 245200 370184
rect 245252 370172 245258 370184
rect 305086 370172 305092 370184
rect 245252 370144 305092 370172
rect 245252 370132 245258 370144
rect 305086 370132 305092 370144
rect 305144 370132 305150 370184
rect 281074 370064 281080 370116
rect 281132 370104 281138 370116
rect 317598 370104 317604 370116
rect 281132 370076 317604 370104
rect 281132 370064 281138 370076
rect 317598 370064 317604 370076
rect 317656 370064 317662 370116
rect 318978 370064 318984 370116
rect 319036 370104 319042 370116
rect 320036 370104 320042 370116
rect 319036 370076 320042 370104
rect 319036 370064 319042 370076
rect 320036 370064 320042 370076
rect 320094 370064 320100 370116
rect 320266 370064 320272 370116
rect 320324 370104 320330 370116
rect 321508 370104 321514 370116
rect 320324 370076 321514 370104
rect 320324 370064 320330 370076
rect 321508 370064 321514 370076
rect 321566 370064 321572 370116
rect 238018 369996 238024 370048
rect 238076 370036 238082 370048
rect 298094 370036 298100 370048
rect 238076 370008 298100 370036
rect 238076 369996 238082 370008
rect 298094 369996 298100 370008
rect 298152 369996 298158 370048
rect 301038 369996 301044 370048
rect 301096 370036 301102 370048
rect 301866 370036 301872 370048
rect 301096 370008 301872 370036
rect 301096 369996 301102 370008
rect 301866 369996 301872 370008
rect 301924 370036 301930 370048
rect 340506 370036 340512 370048
rect 301924 370008 340512 370036
rect 301924 369996 301930 370008
rect 340506 369996 340512 370008
rect 340564 369996 340570 370048
rect 293034 369928 293040 369980
rect 293092 369968 293098 369980
rect 534718 369968 534724 369980
rect 293092 369940 534724 369968
rect 293092 369928 293098 369940
rect 534718 369928 534724 369940
rect 534776 369928 534782 369980
rect 292574 369860 292580 369912
rect 292632 369900 292638 369912
rect 577590 369900 577596 369912
rect 292632 369872 577596 369900
rect 292632 369860 292638 369872
rect 577590 369860 577596 369872
rect 577648 369860 577654 369912
rect 291562 369792 291568 369844
rect 291620 369832 291626 369844
rect 340874 369832 340880 369844
rect 291620 369804 340880 369832
rect 291620 369792 291626 369804
rect 340874 369792 340880 369804
rect 340932 369792 340938 369844
rect 304718 369724 304724 369776
rect 304776 369764 304782 369776
rect 305086 369764 305092 369776
rect 304776 369736 305092 369764
rect 304776 369724 304782 369736
rect 305086 369724 305092 369736
rect 305144 369724 305150 369776
rect 317598 369724 317604 369776
rect 317656 369764 317662 369776
rect 318058 369764 318064 369776
rect 317656 369736 318064 369764
rect 317656 369724 317662 369736
rect 318058 369724 318064 369736
rect 318116 369724 318122 369776
rect 291930 369588 291936 369640
rect 291988 369628 291994 369640
rect 292206 369628 292212 369640
rect 291988 369600 292212 369628
rect 291988 369588 291994 369600
rect 292206 369588 292212 369600
rect 292264 369628 292270 369640
rect 292264 369600 309134 369628
rect 292264 369588 292270 369600
rect 301406 369560 301412 369572
rect 296180 369532 301412 369560
rect 288986 369424 288992 369436
rect 282886 369396 288992 369424
rect 233970 369112 233976 369164
rect 234028 369152 234034 369164
rect 281442 369152 281448 369164
rect 234028 369124 281448 369152
rect 234028 369112 234034 369124
rect 281442 369112 281448 369124
rect 281500 369112 281506 369164
rect 229830 368636 229836 368688
rect 229888 368676 229894 368688
rect 282886 368676 282914 369396
rect 288986 369384 288992 369396
rect 289044 369384 289050 369436
rect 291470 369424 291476 369436
rect 289786 369396 291476 369424
rect 289786 369356 289814 369396
rect 291470 369384 291476 369396
rect 291528 369384 291534 369436
rect 296180 369356 296208 369532
rect 301406 369520 301412 369532
rect 301464 369520 301470 369572
rect 296346 369452 296352 369504
rect 296404 369492 296410 369504
rect 309106 369492 309134 369600
rect 310606 369588 310612 369640
rect 310664 369628 310670 369640
rect 310974 369628 310980 369640
rect 310664 369600 310980 369628
rect 310664 369588 310670 369600
rect 310974 369588 310980 369600
rect 311032 369588 311038 369640
rect 296404 369464 296576 369492
rect 296404 369452 296410 369464
rect 296548 369424 296576 369464
rect 298066 369464 307156 369492
rect 309106 369464 311894 369492
rect 298066 369424 298094 369464
rect 296548 369396 298094 369424
rect 306926 369384 306932 369436
rect 306984 369384 306990 369436
rect 229888 368648 282914 368676
rect 288544 369328 289814 369356
rect 292546 369328 296208 369356
rect 229888 368636 229894 368648
rect 231118 368568 231124 368620
rect 231176 368608 231182 368620
rect 288544 368608 288572 369328
rect 231176 368580 288572 368608
rect 231176 368568 231182 368580
rect 240134 368500 240140 368552
rect 240192 368540 240198 368552
rect 292546 368540 292574 369328
rect 240192 368512 292574 368540
rect 306944 368540 306972 369384
rect 307128 368676 307156 369464
rect 311866 369152 311894 369464
rect 340874 369180 340880 369232
rect 340932 369220 340938 369232
rect 342162 369220 342168 369232
rect 340932 369192 342168 369220
rect 340932 369180 340938 369192
rect 342162 369180 342168 369192
rect 342220 369220 342226 369232
rect 580626 369220 580632 369232
rect 342220 369192 580632 369220
rect 342220 369180 342226 369192
rect 580626 369180 580632 369192
rect 580684 369180 580690 369232
rect 580350 369152 580356 369164
rect 311866 369124 580356 369152
rect 580350 369112 580356 369124
rect 580408 369112 580414 369164
rect 307128 368648 311894 368676
rect 311866 368608 311894 368648
rect 327902 368608 327908 368620
rect 311866 368580 327908 368608
rect 327902 368568 327908 368580
rect 327960 368568 327966 368620
rect 339310 368540 339316 368552
rect 306944 368512 339316 368540
rect 240192 368500 240198 368512
rect 339310 368500 339316 368512
rect 339368 368500 339374 368552
rect 201494 367752 201500 367804
rect 201552 367792 201558 367804
rect 245654 367792 245660 367804
rect 201552 367764 245660 367792
rect 201552 367752 201558 367764
rect 245654 367752 245660 367764
rect 245712 367752 245718 367804
rect 245654 367004 245660 367056
rect 245712 367044 245718 367056
rect 246298 367044 246304 367056
rect 245712 367016 246304 367044
rect 245712 367004 245718 367016
rect 246298 367004 246304 367016
rect 246356 367044 246362 367056
rect 279878 367044 279884 367056
rect 246356 367016 279884 367044
rect 246356 367004 246362 367016
rect 279878 367004 279884 367016
rect 279936 367004 279942 367056
rect 329742 366324 329748 366376
rect 329800 366364 329806 366376
rect 384022 366364 384028 366376
rect 329800 366336 384028 366364
rect 329800 366324 329806 366336
rect 384022 366324 384028 366336
rect 384080 366324 384086 366376
rect 329650 365644 329656 365696
rect 329708 365684 329714 365696
rect 580166 365684 580172 365696
rect 329708 365656 580172 365684
rect 329708 365644 329714 365656
rect 580166 365644 580172 365656
rect 580224 365644 580230 365696
rect 247034 365032 247040 365084
rect 247092 365072 247098 365084
rect 274542 365072 274548 365084
rect 247092 365044 274548 365072
rect 247092 365032 247098 365044
rect 274542 365032 274548 365044
rect 274600 365032 274606 365084
rect 247678 364964 247684 365016
rect 247736 365004 247742 365016
rect 280154 365004 280160 365016
rect 247736 364976 280160 365004
rect 247736 364964 247742 364976
rect 280154 364964 280160 364976
rect 280212 364964 280218 365016
rect 249150 363604 249156 363656
rect 249208 363644 249214 363656
rect 277302 363644 277308 363656
rect 249208 363616 277308 363644
rect 249208 363604 249214 363616
rect 277302 363604 277308 363616
rect 277360 363604 277366 363656
rect 334986 362176 334992 362228
rect 335044 362216 335050 362228
rect 350810 362216 350816 362228
rect 335044 362188 350816 362216
rect 335044 362176 335050 362188
rect 350810 362176 350816 362188
rect 350868 362176 350874 362228
rect 253382 360816 253388 360868
rect 253440 360856 253446 360868
rect 280614 360856 280620 360868
rect 253440 360828 280620 360856
rect 253440 360816 253446 360828
rect 280614 360816 280620 360828
rect 280672 360816 280678 360868
rect 333514 359524 333520 359576
rect 333572 359564 333578 359576
rect 352098 359564 352104 359576
rect 333572 359536 352104 359564
rect 333572 359524 333578 359536
rect 352098 359524 352104 359536
rect 352156 359524 352162 359576
rect 256786 359456 256792 359508
rect 256844 359496 256850 359508
rect 280706 359496 280712 359508
rect 256844 359468 280712 359496
rect 256844 359456 256850 359468
rect 280706 359456 280712 359468
rect 280764 359456 280770 359508
rect 329650 359456 329656 359508
rect 329708 359496 329714 359508
rect 385402 359496 385408 359508
rect 329708 359468 385408 359496
rect 329708 359456 329714 359468
rect 385402 359456 385408 359468
rect 385460 359456 385466 359508
rect 226978 358776 226984 358828
rect 227036 358816 227042 358828
rect 277670 358816 277676 358828
rect 227036 358788 277676 358816
rect 227036 358776 227042 358788
rect 277670 358776 277676 358788
rect 277728 358816 277734 358828
rect 279418 358816 279424 358828
rect 277728 358788 279424 358816
rect 277728 358776 277734 358788
rect 279418 358776 279424 358788
rect 279476 358776 279482 358828
rect 271046 358708 271052 358760
rect 271104 358748 271110 358760
rect 277854 358748 277860 358760
rect 271104 358720 277860 358748
rect 271104 358708 271110 358720
rect 277854 358708 277860 358720
rect 277912 358708 277918 358760
rect 3142 357416 3148 357468
rect 3200 357456 3206 357468
rect 271046 357456 271052 357468
rect 3200 357428 271052 357456
rect 3200 357416 3206 357428
rect 271046 357416 271052 357428
rect 271104 357416 271110 357468
rect 253290 356668 253296 356720
rect 253348 356708 253354 356720
rect 280706 356708 280712 356720
rect 253348 356680 280712 356708
rect 253348 356668 253354 356680
rect 280706 356668 280712 356680
rect 280764 356668 280770 356720
rect 333790 356668 333796 356720
rect 333848 356708 333854 356720
rect 350718 356708 350724 356720
rect 333848 356680 350724 356708
rect 333848 356668 333854 356680
rect 350718 356668 350724 356680
rect 350776 356668 350782 356720
rect 256050 355308 256056 355360
rect 256108 355348 256114 355360
rect 279234 355348 279240 355360
rect 256108 355320 279240 355348
rect 256108 355308 256114 355320
rect 279234 355308 279240 355320
rect 279292 355308 279298 355360
rect 227070 351160 227076 351212
rect 227128 351200 227134 351212
rect 279326 351200 279332 351212
rect 227128 351172 279332 351200
rect 227128 351160 227134 351172
rect 279326 351160 279332 351172
rect 279384 351160 279390 351212
rect 383838 349052 383844 349104
rect 383896 349092 383902 349104
rect 384390 349092 384396 349104
rect 383896 349064 384396 349092
rect 383896 349052 383902 349064
rect 384390 349052 384396 349064
rect 384448 349052 384454 349104
rect 384390 347760 384396 347812
rect 384448 347800 384454 347812
rect 534074 347800 534080 347812
rect 384448 347772 534080 347800
rect 384448 347760 384454 347772
rect 534074 347760 534080 347772
rect 534132 347760 534138 347812
rect 332042 347012 332048 347064
rect 332100 347052 332106 347064
rect 351546 347052 351552 347064
rect 332100 347024 351552 347052
rect 332100 347012 332106 347024
rect 351546 347012 351552 347024
rect 351604 347012 351610 347064
rect 255406 345652 255412 345704
rect 255464 345692 255470 345704
rect 280706 345692 280712 345704
rect 255464 345664 280712 345692
rect 255464 345652 255470 345664
rect 280706 345652 280712 345664
rect 280764 345652 280770 345704
rect 3326 345040 3332 345092
rect 3384 345080 3390 345092
rect 255406 345080 255412 345092
rect 3384 345052 255412 345080
rect 3384 345040 3390 345052
rect 255406 345040 255412 345052
rect 255464 345040 255470 345092
rect 332226 342864 332232 342916
rect 332284 342904 332290 342916
rect 350258 342904 350264 342916
rect 332284 342876 350264 342904
rect 332284 342864 332290 342876
rect 350258 342864 350264 342876
rect 350316 342864 350322 342916
rect 332502 340144 332508 340196
rect 332560 340184 332566 340196
rect 351638 340184 351644 340196
rect 332560 340156 351644 340184
rect 332560 340144 332566 340156
rect 351638 340144 351644 340156
rect 351696 340144 351702 340196
rect 329006 338716 329012 338768
rect 329064 338756 329070 338768
rect 386966 338756 386972 338768
rect 329064 338728 386972 338756
rect 329064 338716 329070 338728
rect 386966 338716 386972 338728
rect 387024 338716 387030 338768
rect 350258 335996 350264 336048
rect 350316 336036 350322 336048
rect 368750 336036 368756 336048
rect 350316 336008 368756 336036
rect 350316 335996 350322 336008
rect 368750 335996 368756 336008
rect 368808 335996 368814 336048
rect 336458 334568 336464 334620
rect 336516 334608 336522 334620
rect 377030 334608 377036 334620
rect 336516 334580 377036 334608
rect 336516 334568 336522 334580
rect 377030 334568 377036 334580
rect 377088 334568 377094 334620
rect 385218 333956 385224 334008
rect 385276 333996 385282 334008
rect 385678 333996 385684 334008
rect 385276 333968 385684 333996
rect 385276 333956 385282 333968
rect 385678 333956 385684 333968
rect 385736 333996 385742 334008
rect 552014 333996 552020 334008
rect 385736 333968 552020 333996
rect 385736 333956 385742 333968
rect 552014 333956 552020 333968
rect 552072 333956 552078 334008
rect 335170 333208 335176 333260
rect 335228 333248 335234 333260
rect 371786 333248 371792 333260
rect 335228 333220 371792 333248
rect 335228 333208 335234 333220
rect 371786 333208 371792 333220
rect 371844 333208 371850 333260
rect 379698 331236 379704 331288
rect 379756 331276 379762 331288
rect 481634 331276 481640 331288
rect 379756 331248 481640 331276
rect 379756 331236 379762 331248
rect 481634 331236 481640 331248
rect 481692 331236 481698 331288
rect 331122 329060 331128 329112
rect 331180 329100 331186 329112
rect 345566 329100 345572 329112
rect 331180 329072 345572 329100
rect 331180 329060 331186 329072
rect 345566 329060 345572 329072
rect 345624 329060 345630 329112
rect 235350 327700 235356 327752
rect 235408 327740 235414 327752
rect 277946 327740 277952 327752
rect 235408 327712 277952 327740
rect 235408 327700 235414 327712
rect 277946 327700 277952 327712
rect 278004 327700 278010 327752
rect 380894 327088 380900 327140
rect 380952 327128 380958 327140
rect 381354 327128 381360 327140
rect 380952 327100 381360 327128
rect 380952 327088 380958 327100
rect 381354 327088 381360 327100
rect 381412 327128 381418 327140
rect 495434 327128 495440 327140
rect 381412 327100 495440 327128
rect 381412 327088 381418 327100
rect 495434 327088 495440 327100
rect 495492 327088 495498 327140
rect 336918 326340 336924 326392
rect 336976 326380 336982 326392
rect 375650 326380 375656 326392
rect 336976 326352 375656 326380
rect 336976 326340 336982 326352
rect 375650 326340 375656 326352
rect 375708 326340 375714 326392
rect 577590 325456 577596 325508
rect 577648 325496 577654 325508
rect 580718 325496 580724 325508
rect 577648 325468 580724 325496
rect 577648 325456 577654 325468
rect 580718 325456 580724 325468
rect 580776 325456 580782 325508
rect 234062 324912 234068 324964
rect 234120 324952 234126 324964
rect 279510 324952 279516 324964
rect 234120 324924 279516 324952
rect 234120 324912 234126 324924
rect 279510 324912 279516 324924
rect 279568 324912 279574 324964
rect 385770 324300 385776 324352
rect 385828 324340 385834 324352
rect 547966 324340 547972 324352
rect 385828 324312 547972 324340
rect 385828 324300 385834 324312
rect 547966 324300 547972 324312
rect 548024 324300 548030 324352
rect 339310 323620 339316 323672
rect 339368 323660 339374 323672
rect 378410 323660 378416 323672
rect 339368 323632 378416 323660
rect 339368 323620 339374 323632
rect 378410 323620 378416 323632
rect 378468 323620 378474 323672
rect 335078 323552 335084 323604
rect 335136 323592 335142 323604
rect 374362 323592 374368 323604
rect 335136 323564 374368 323592
rect 335136 323552 335142 323564
rect 374362 323552 374368 323564
rect 374420 323552 374426 323604
rect 380894 323008 380900 323060
rect 380952 323048 380958 323060
rect 381262 323048 381268 323060
rect 380952 323020 381268 323048
rect 380952 323008 380958 323020
rect 381262 323008 381268 323020
rect 381320 323048 381326 323060
rect 381320 323020 383654 323048
rect 381320 323008 381326 323020
rect 381538 322940 381544 322992
rect 381596 322980 381602 322992
rect 383378 322980 383384 322992
rect 381596 322952 383384 322980
rect 381596 322940 381602 322952
rect 383378 322940 383384 322952
rect 383436 322940 383442 322992
rect 383626 322980 383654 323020
rect 506474 322980 506480 322992
rect 383626 322952 506480 322980
rect 506474 322940 506480 322952
rect 506532 322940 506538 322992
rect 272242 322260 272248 322312
rect 272300 322300 272306 322312
rect 273162 322300 273168 322312
rect 272300 322272 273168 322300
rect 272300 322260 272306 322272
rect 273162 322260 273168 322272
rect 273220 322260 273226 322312
rect 339954 322260 339960 322312
rect 340012 322300 340018 322312
rect 363690 322300 363696 322312
rect 340012 322272 363696 322300
rect 340012 322260 340018 322272
rect 363690 322260 363696 322272
rect 363748 322260 363754 322312
rect 228450 322192 228456 322244
rect 228508 322232 228514 322244
rect 278038 322232 278044 322244
rect 228508 322204 278044 322232
rect 228508 322192 228514 322204
rect 278038 322192 278044 322204
rect 278096 322192 278102 322244
rect 334066 322192 334072 322244
rect 334124 322232 334130 322244
rect 380894 322232 380900 322244
rect 334124 322204 380900 322232
rect 334124 322192 334130 322204
rect 380894 322192 380900 322204
rect 380952 322192 380958 322244
rect 272518 322124 272524 322176
rect 272576 322164 272582 322176
rect 273162 322164 273168 322176
rect 272576 322136 273168 322164
rect 272576 322124 272582 322136
rect 273162 322124 273168 322136
rect 273220 322124 273226 322176
rect 218698 321716 218704 321768
rect 218756 321756 218762 321768
rect 268562 321756 268568 321768
rect 218756 321728 268568 321756
rect 218756 321716 218762 321728
rect 268562 321716 268568 321728
rect 268620 321716 268626 321768
rect 206738 321648 206744 321700
rect 206796 321688 206802 321700
rect 272518 321688 272524 321700
rect 206796 321660 272524 321688
rect 206796 321648 206802 321660
rect 272518 321648 272524 321660
rect 272576 321648 272582 321700
rect 201402 321580 201408 321632
rect 201460 321620 201466 321632
rect 269850 321620 269856 321632
rect 201460 321592 269856 321620
rect 201460 321580 201466 321592
rect 269850 321580 269856 321592
rect 269908 321620 269914 321632
rect 270310 321620 270316 321632
rect 269908 321592 270316 321620
rect 269908 321580 269914 321592
rect 270310 321580 270316 321592
rect 270368 321580 270374 321632
rect 327902 321376 327908 321428
rect 327960 321416 327966 321428
rect 328178 321416 328184 321428
rect 327960 321388 328184 321416
rect 327960 321376 327966 321388
rect 328178 321376 328184 321388
rect 328236 321376 328242 321428
rect 271322 321104 271328 321156
rect 271380 321144 271386 321156
rect 271598 321144 271604 321156
rect 271380 321116 271604 321144
rect 271380 321104 271386 321116
rect 271598 321104 271604 321116
rect 271656 321104 271662 321156
rect 327810 321104 327816 321156
rect 327868 321144 327874 321156
rect 328086 321144 328092 321156
rect 327868 321116 328092 321144
rect 327868 321104 327874 321116
rect 328086 321104 328092 321116
rect 328144 321104 328150 321156
rect 276750 321076 276756 321088
rect 273226 321048 276756 321076
rect 271598 320968 271604 321020
rect 271656 321008 271662 321020
rect 271782 321008 271788 321020
rect 271656 320980 271788 321008
rect 271656 320968 271662 320980
rect 271782 320968 271788 320980
rect 271840 320968 271846 321020
rect 272978 320900 272984 320952
rect 273036 320940 273042 320952
rect 273226 320940 273254 321048
rect 276750 321036 276756 321048
rect 276808 321076 276814 321088
rect 276808 321048 299934 321076
rect 276808 321036 276814 321048
rect 273036 320912 273254 320940
rect 273036 320900 273042 320912
rect 299906 320748 299934 321048
rect 324286 321048 325694 321076
rect 324286 321008 324314 321048
rect 302206 320980 324314 321008
rect 325666 321008 325694 321048
rect 337010 321036 337016 321088
rect 337068 321076 337074 321088
rect 368658 321076 368664 321088
rect 337068 321048 368664 321076
rect 337068 321036 337074 321048
rect 368658 321036 368664 321048
rect 368716 321036 368722 321088
rect 353386 321008 353392 321020
rect 325666 320980 353392 321008
rect 299888 320696 299894 320748
rect 299946 320696 299952 320748
rect 302206 320668 302234 320980
rect 353386 320968 353392 320980
rect 353444 320968 353450 321020
rect 333146 320900 333152 320952
rect 333204 320940 333210 320952
rect 359550 320940 359556 320952
rect 333204 320912 359556 320940
rect 333204 320900 333210 320912
rect 359550 320900 359556 320912
rect 359608 320900 359614 320952
rect 357434 320872 357440 320884
rect 325666 320844 328454 320872
rect 325666 320804 325694 320844
rect 273226 320640 297036 320668
rect 217870 320492 217876 320544
rect 217928 320532 217934 320544
rect 273226 320532 273254 320640
rect 281626 320560 281632 320612
rect 281684 320600 281690 320612
rect 282270 320600 282276 320612
rect 281684 320572 282276 320600
rect 281684 320560 281690 320572
rect 282270 320560 282276 320572
rect 282328 320560 282334 320612
rect 217928 320504 273254 320532
rect 217928 320492 217934 320504
rect 276842 320424 276848 320476
rect 276900 320464 276906 320476
rect 282178 320464 282184 320476
rect 276900 320436 282184 320464
rect 276900 320424 276906 320436
rect 282178 320424 282184 320436
rect 282236 320424 282242 320476
rect 220538 320220 220544 320272
rect 220596 320260 220602 320272
rect 220596 320232 294138 320260
rect 220596 320220 220602 320232
rect 282178 320152 282184 320204
rect 282236 320192 282242 320204
rect 282236 320164 293908 320192
rect 282236 320152 282242 320164
rect 278498 320084 278504 320136
rect 278556 320124 278562 320136
rect 278556 320096 289906 320124
rect 278556 320084 278562 320096
rect 279970 319948 279976 320000
rect 280028 319988 280034 320000
rect 282178 319988 282184 320000
rect 280028 319960 282184 319988
rect 280028 319948 280034 319960
rect 282178 319948 282184 319960
rect 282236 319948 282242 320000
rect 287302 319960 289814 319988
rect 278038 319880 278044 319932
rect 278096 319920 278102 319932
rect 278096 319892 287146 319920
rect 278096 319880 278102 319892
rect 287118 319796 287146 319892
rect 281902 319744 281908 319796
rect 281960 319784 281966 319796
rect 282362 319784 282368 319796
rect 281960 319756 282368 319784
rect 281960 319744 281966 319756
rect 282362 319744 282368 319756
rect 282420 319744 282426 319796
rect 287118 319756 287152 319796
rect 287146 319744 287152 319756
rect 287204 319744 287210 319796
rect 273898 319716 273904 319728
rect 258046 319688 273904 319716
rect 216306 319540 216312 319592
rect 216364 319580 216370 319592
rect 258046 319580 258074 319688
rect 273898 319676 273904 319688
rect 273956 319716 273962 319728
rect 287302 319716 287330 319960
rect 289032 319880 289038 319932
rect 289090 319880 289096 319932
rect 289050 319852 289078 319880
rect 288912 319824 289078 319852
rect 289786 319852 289814 319960
rect 289878 319920 289906 320096
rect 289878 319892 293816 319920
rect 289786 319824 291700 319852
rect 273956 319688 287330 319716
rect 273956 319676 273962 319688
rect 288802 319676 288808 319728
rect 288860 319716 288866 319728
rect 288912 319716 288940 319824
rect 291672 319784 291700 319824
rect 293494 319784 293500 319796
rect 291672 319756 293500 319784
rect 293494 319744 293500 319756
rect 293552 319744 293558 319796
rect 288860 319688 288940 319716
rect 293788 319716 293816 319892
rect 293880 319784 293908 320164
rect 294110 319852 294138 320232
rect 294506 319880 294512 319932
rect 294564 319920 294570 319932
rect 295012 319920 295018 319932
rect 294564 319892 295018 319920
rect 294564 319880 294570 319892
rect 295012 319880 295018 319892
rect 295070 319880 295076 319932
rect 295748 319920 295754 319932
rect 295306 319892 295754 319920
rect 294782 319852 294788 319864
rect 294110 319824 294788 319852
rect 294782 319812 294788 319824
rect 294840 319812 294846 319864
rect 295306 319784 295334 319892
rect 295748 319880 295754 319892
rect 295806 319880 295812 319932
rect 296852 319880 296858 319932
rect 296910 319880 296916 319932
rect 293880 319756 295334 319784
rect 296870 319716 296898 319880
rect 297008 319784 297036 320640
rect 298388 320640 302234 320668
rect 310486 320776 325694 320804
rect 328426 320804 328454 320844
rect 336108 320844 357440 320872
rect 336108 320804 336136 320844
rect 357434 320832 357440 320844
rect 357492 320832 357498 320884
rect 328426 320776 336136 320804
rect 297082 319812 297088 319864
rect 297140 319852 297146 319864
rect 298388 319852 298416 320640
rect 310486 320532 310514 320776
rect 333146 320736 333152 320748
rect 309244 320504 310514 320532
rect 310578 320708 333152 320736
rect 309244 320396 309272 320504
rect 310578 320464 310606 320708
rect 333146 320696 333152 320708
rect 333204 320696 333210 320748
rect 328454 320668 328460 320680
rect 298802 320368 309272 320396
rect 310072 320436 310606 320464
rect 317386 320640 328460 320668
rect 298802 319932 298830 320368
rect 310072 320260 310100 320436
rect 317386 320396 317414 320640
rect 328454 320628 328460 320640
rect 328512 320628 328518 320680
rect 327626 320492 327632 320544
rect 327684 320532 327690 320544
rect 327684 320504 328454 320532
rect 327684 320492 327690 320504
rect 328426 320396 328454 320504
rect 335538 320396 335544 320408
rect 301470 320232 310100 320260
rect 310164 320368 317414 320396
rect 322308 320368 322934 320396
rect 328426 320368 335544 320396
rect 301470 320124 301498 320232
rect 300182 320096 301498 320124
rect 300182 319932 300210 320096
rect 302160 319960 309134 319988
rect 298784 319920 298790 319932
rect 297140 319824 298416 319852
rect 298480 319892 298790 319920
rect 297140 319812 297146 319824
rect 298480 319784 298508 319892
rect 298784 319880 298790 319892
rect 298842 319880 298848 319932
rect 300164 319880 300170 319932
rect 300222 319880 300228 319932
rect 301544 319880 301550 319932
rect 301602 319880 301608 319932
rect 298554 319812 298560 319864
rect 298612 319852 298618 319864
rect 300182 319852 300210 319880
rect 298612 319824 300210 319852
rect 298612 319812 298618 319824
rect 300532 319812 300538 319864
rect 300590 319852 300596 319864
rect 300762 319852 300768 319864
rect 300590 319824 300768 319852
rect 300590 319812 300596 319824
rect 300762 319812 300768 319824
rect 300820 319812 300826 319864
rect 301314 319784 301320 319796
rect 297008 319756 298508 319784
rect 301148 319756 301320 319784
rect 293788 319688 296898 319716
rect 288860 319676 288866 319688
rect 301148 319660 301176 319756
rect 301314 319744 301320 319756
rect 301372 319744 301378 319796
rect 301562 319784 301590 319880
rect 302160 319864 302188 319960
rect 302372 319880 302378 319932
rect 302430 319880 302436 319932
rect 303016 319880 303022 319932
rect 303074 319880 303080 319932
rect 303200 319880 303206 319932
rect 303258 319880 303264 319932
rect 304028 319880 304034 319932
rect 304086 319880 304092 319932
rect 304304 319880 304310 319932
rect 304362 319880 304368 319932
rect 304396 319880 304402 319932
rect 304454 319880 304460 319932
rect 305316 319880 305322 319932
rect 305374 319880 305380 319932
rect 306788 319920 306794 319932
rect 306346 319892 306794 319920
rect 302142 319812 302148 319864
rect 302200 319812 302206 319864
rect 302234 319784 302240 319796
rect 301562 319756 301820 319784
rect 280062 319608 280068 319660
rect 280120 319648 280126 319660
rect 292482 319648 292488 319660
rect 280120 319620 292488 319648
rect 280120 319608 280126 319620
rect 292482 319608 292488 319620
rect 292540 319608 292546 319660
rect 292666 319608 292672 319660
rect 292724 319648 292730 319660
rect 296898 319648 296904 319660
rect 292724 319620 296904 319648
rect 292724 319608 292730 319620
rect 296898 319608 296904 319620
rect 296956 319608 296962 319660
rect 299750 319608 299756 319660
rect 299808 319648 299814 319660
rect 300854 319648 300860 319660
rect 299808 319620 300860 319648
rect 299808 319608 299814 319620
rect 300854 319608 300860 319620
rect 300912 319608 300918 319660
rect 301130 319608 301136 319660
rect 301188 319608 301194 319660
rect 216364 319552 258074 319580
rect 216364 319540 216370 319552
rect 276566 319540 276572 319592
rect 276624 319580 276630 319592
rect 300946 319580 300952 319592
rect 276624 319552 300952 319580
rect 276624 319540 276630 319552
rect 300946 319540 300952 319552
rect 301004 319540 301010 319592
rect 301498 319540 301504 319592
rect 301556 319580 301562 319592
rect 301792 319580 301820 319756
rect 301556 319552 301820 319580
rect 302160 319756 302240 319784
rect 302160 319580 302188 319756
rect 302234 319744 302240 319756
rect 302292 319744 302298 319796
rect 302234 319608 302240 319660
rect 302292 319648 302298 319660
rect 302390 319648 302418 319880
rect 302464 319812 302470 319864
rect 302522 319812 302528 319864
rect 302292 319620 302418 319648
rect 302482 319648 302510 319812
rect 302482 319620 302648 319648
rect 302292 319608 302298 319620
rect 302620 319592 302648 319620
rect 302326 319580 302332 319592
rect 302160 319552 302332 319580
rect 301556 319540 301562 319552
rect 302326 319540 302332 319552
rect 302384 319540 302390 319592
rect 302602 319540 302608 319592
rect 302660 319540 302666 319592
rect 302786 319540 302792 319592
rect 302844 319580 302850 319592
rect 303034 319580 303062 319880
rect 303218 319592 303246 319880
rect 303660 319812 303666 319864
rect 303718 319812 303724 319864
rect 303678 319728 303706 319812
rect 304046 319728 304074 319880
rect 303614 319676 303620 319728
rect 303672 319688 303706 319728
rect 303672 319676 303678 319688
rect 303982 319676 303988 319728
rect 304040 319688 304074 319728
rect 304040 319676 304046 319688
rect 303338 319608 303344 319660
rect 303396 319648 303402 319660
rect 304322 319648 304350 319880
rect 303396 319620 304350 319648
rect 303396 319608 303402 319620
rect 304414 319592 304442 319880
rect 304488 319812 304494 319864
rect 304546 319812 304552 319864
rect 304856 319812 304862 319864
rect 304914 319812 304920 319864
rect 302844 319552 303062 319580
rect 302844 319540 302850 319552
rect 303154 319540 303160 319592
rect 303212 319552 303246 319592
rect 303212 319540 303218 319552
rect 304350 319540 304356 319592
rect 304408 319552 304442 319592
rect 304408 319540 304414 319552
rect 304506 319524 304534 319812
rect 304874 319660 304902 319812
rect 304810 319608 304816 319660
rect 304868 319620 304902 319660
rect 305334 319648 305362 319880
rect 306236 319812 306242 319864
rect 306294 319812 306300 319864
rect 305454 319676 305460 319728
rect 305512 319716 305518 319728
rect 306254 319716 306282 319812
rect 305512 319688 306282 319716
rect 305512 319676 305518 319688
rect 305822 319648 305828 319660
rect 305334 319620 305828 319648
rect 304868 319608 304874 319620
rect 305822 319608 305828 319620
rect 305880 319608 305886 319660
rect 272886 319512 272892 319524
rect 258046 319484 272892 319512
rect 211062 319404 211068 319456
rect 211120 319444 211126 319456
rect 258046 319444 258074 319484
rect 272886 319472 272892 319484
rect 272944 319512 272950 319524
rect 293126 319512 293132 319524
rect 272944 319484 293132 319512
rect 272944 319472 272950 319484
rect 293126 319472 293132 319484
rect 293184 319472 293190 319524
rect 294598 319472 294604 319524
rect 294656 319512 294662 319524
rect 294966 319512 294972 319524
rect 294656 319484 294972 319512
rect 294656 319472 294662 319484
rect 294966 319472 294972 319484
rect 295024 319472 295030 319524
rect 295886 319472 295892 319524
rect 295944 319512 295950 319524
rect 296162 319512 296168 319524
rect 295944 319484 296168 319512
rect 295944 319472 295950 319484
rect 296162 319472 296168 319484
rect 296220 319472 296226 319524
rect 296898 319472 296904 319524
rect 296956 319512 296962 319524
rect 298094 319512 298100 319524
rect 296956 319484 298100 319512
rect 296956 319472 296962 319484
rect 298094 319472 298100 319484
rect 298152 319472 298158 319524
rect 299446 319484 302556 319512
rect 211120 319416 258074 319444
rect 211120 319404 211126 319416
rect 273806 319404 273812 319456
rect 273864 319444 273870 319456
rect 299446 319444 299474 319484
rect 273864 319416 299474 319444
rect 302528 319444 302556 319484
rect 304442 319472 304448 319524
rect 304500 319484 304534 319524
rect 304500 319472 304506 319484
rect 306346 319444 306374 319892
rect 306788 319880 306794 319892
rect 306846 319880 306852 319932
rect 307432 319880 307438 319932
rect 307490 319880 307496 319932
rect 307524 319880 307530 319932
rect 307582 319880 307588 319932
rect 307450 319784 307478 319880
rect 306576 319756 307478 319784
rect 306576 319728 306604 319756
rect 307542 319728 307570 319880
rect 306558 319676 306564 319728
rect 306616 319676 306622 319728
rect 307478 319676 307484 319728
rect 307536 319688 307570 319728
rect 307536 319676 307542 319688
rect 309106 319512 309134 319960
rect 310164 319864 310192 320368
rect 322308 320328 322336 320368
rect 310532 320300 322336 320328
rect 322906 320328 322934 320368
rect 335538 320356 335544 320368
rect 335596 320356 335602 320408
rect 342346 320328 342352 320340
rect 322906 320300 342352 320328
rect 310238 319880 310244 319932
rect 310296 319880 310302 319932
rect 310146 319812 310152 319864
rect 310204 319812 310210 319864
rect 310256 319580 310284 319880
rect 310532 319660 310560 320300
rect 342346 320288 342352 320300
rect 342404 320288 342410 320340
rect 328454 320220 328460 320272
rect 328512 320260 328518 320272
rect 335446 320260 335452 320272
rect 328512 320232 335452 320260
rect 328512 320220 328518 320232
rect 335446 320220 335452 320232
rect 335504 320220 335510 320272
rect 337010 320192 337016 320204
rect 311912 320164 337016 320192
rect 311204 319920 311210 319932
rect 310624 319892 311210 319920
rect 310624 319660 310652 319892
rect 311204 319880 311210 319892
rect 311262 319880 311268 319932
rect 311912 319660 311940 320164
rect 337010 320152 337016 320164
rect 337068 320152 337074 320204
rect 328270 320124 328276 320136
rect 318766 320096 328276 320124
rect 318766 320056 318794 320096
rect 328270 320084 328276 320096
rect 328328 320084 328334 320136
rect 327626 320056 327632 320068
rect 318444 320028 318794 320056
rect 325114 320028 327632 320056
rect 313384 319960 314102 319988
rect 313136 319920 313142 319932
rect 312004 319892 313142 319920
rect 312004 319864 312032 319892
rect 313136 319880 313142 319892
rect 313194 319880 313200 319932
rect 311986 319812 311992 319864
rect 312044 319812 312050 319864
rect 310514 319608 310520 319660
rect 310572 319608 310578 319660
rect 310606 319608 310612 319660
rect 310664 319608 310670 319660
rect 311894 319608 311900 319660
rect 311952 319608 311958 319660
rect 310330 319580 310336 319592
rect 310256 319552 310336 319580
rect 310330 319540 310336 319552
rect 310388 319540 310394 319592
rect 312262 319540 312268 319592
rect 312320 319580 312326 319592
rect 313182 319580 313188 319592
rect 312320 319552 313188 319580
rect 312320 319540 312326 319552
rect 313182 319540 313188 319552
rect 313240 319540 313246 319592
rect 313384 319580 313412 319960
rect 314074 319932 314102 319960
rect 313780 319880 313786 319932
rect 313838 319880 313844 319932
rect 314056 319880 314062 319932
rect 314114 319880 314120 319932
rect 314608 319880 314614 319932
rect 314666 319880 314672 319932
rect 314700 319880 314706 319932
rect 314758 319880 314764 319932
rect 315344 319880 315350 319932
rect 315402 319880 315408 319932
rect 315528 319880 315534 319932
rect 315586 319920 315592 319932
rect 317276 319920 317282 319932
rect 315586 319880 315620 319920
rect 313798 319852 313826 319880
rect 313798 319824 314378 319852
rect 314350 319592 314378 319824
rect 314626 319660 314654 319880
rect 314562 319608 314568 319660
rect 314620 319620 314654 319660
rect 314620 319608 314626 319620
rect 313550 319580 313556 319592
rect 313384 319552 313556 319580
rect 313550 319540 313556 319552
rect 313608 319540 313614 319592
rect 314350 319552 314384 319592
rect 314378 319540 314384 319552
rect 314436 319540 314442 319592
rect 314718 319580 314746 319880
rect 315114 319608 315120 319660
rect 315172 319648 315178 319660
rect 315362 319648 315390 319880
rect 315592 319660 315620 319880
rect 317248 319880 317282 319920
rect 317334 319880 317340 319932
rect 317828 319920 317834 319932
rect 317800 319880 317834 319920
rect 317886 319880 317892 319932
rect 317248 319796 317276 319880
rect 317800 319796 317828 319880
rect 317920 319812 317926 319864
rect 317978 319812 317984 319864
rect 317138 319744 317144 319796
rect 317196 319744 317202 319796
rect 317230 319744 317236 319796
rect 317288 319744 317294 319796
rect 317782 319744 317788 319796
rect 317840 319744 317846 319796
rect 317156 319660 317184 319744
rect 317938 319728 317966 319812
rect 318242 319744 318248 319796
rect 318300 319784 318306 319796
rect 318444 319784 318472 320028
rect 318300 319756 318472 319784
rect 318766 319960 324130 319988
rect 318300 319744 318306 319756
rect 317874 319676 317880 319728
rect 317932 319688 317966 319728
rect 317932 319676 317938 319688
rect 315172 319620 315390 319648
rect 315172 319608 315178 319620
rect 315574 319608 315580 319660
rect 315632 319608 315638 319660
rect 317138 319608 317144 319660
rect 317196 319608 317202 319660
rect 314838 319580 314844 319592
rect 314718 319552 314844 319580
rect 314838 319540 314844 319552
rect 314896 319540 314902 319592
rect 315482 319540 315488 319592
rect 315540 319580 315546 319592
rect 315666 319580 315672 319592
rect 315540 319552 315672 319580
rect 315540 319540 315546 319552
rect 315666 319540 315672 319552
rect 315724 319540 315730 319592
rect 318766 319580 318794 319960
rect 320864 319880 320870 319932
rect 320922 319880 320928 319932
rect 320956 319880 320962 319932
rect 321014 319880 321020 319932
rect 321416 319920 321422 319932
rect 321342 319892 321422 319920
rect 319576 319812 319582 319864
rect 319634 319812 319640 319864
rect 319852 319812 319858 319864
rect 319910 319812 319916 319864
rect 319594 319660 319622 319812
rect 319870 319660 319898 319812
rect 320726 319744 320732 319796
rect 320784 319784 320790 319796
rect 320882 319784 320910 319880
rect 320784 319756 320910 319784
rect 320784 319744 320790 319756
rect 320974 319728 321002 319880
rect 320910 319676 320916 319728
rect 320968 319688 321002 319728
rect 320968 319676 320974 319688
rect 321342 319660 321370 319892
rect 321416 319880 321422 319892
rect 321474 319880 321480 319932
rect 322152 319880 322158 319932
rect 322210 319880 322216 319932
rect 322796 319880 322802 319932
rect 322854 319880 322860 319932
rect 323992 319880 323998 319932
rect 324050 319880 324056 319932
rect 321692 319852 321698 319864
rect 319594 319620 319628 319660
rect 319622 319608 319628 319620
rect 319680 319608 319686 319660
rect 319870 319620 319904 319660
rect 319898 319608 319904 319620
rect 319956 319608 319962 319660
rect 321278 319608 321284 319660
rect 321336 319620 321370 319660
rect 321572 319824 321698 319852
rect 321336 319608 321342 319620
rect 321572 319592 321600 319824
rect 321692 319812 321698 319824
rect 321750 319812 321756 319864
rect 322014 319784 322020 319796
rect 321756 319756 322020 319784
rect 321756 319660 321784 319756
rect 322014 319744 322020 319756
rect 322072 319744 322078 319796
rect 322170 319716 322198 319880
rect 322704 319812 322710 319864
rect 322762 319812 322768 319864
rect 322722 319784 322750 319812
rect 322032 319688 322198 319716
rect 322584 319756 322750 319784
rect 322032 319660 322060 319688
rect 321738 319608 321744 319660
rect 321796 319608 321802 319660
rect 322014 319608 322020 319660
rect 322072 319608 322078 319660
rect 322198 319608 322204 319660
rect 322256 319648 322262 319660
rect 322474 319648 322480 319660
rect 322256 319620 322480 319648
rect 322256 319608 322262 319620
rect 322474 319608 322480 319620
rect 322532 319608 322538 319660
rect 317432 319552 318794 319580
rect 309106 319484 311894 319512
rect 302528 319416 306374 319444
rect 273864 319404 273870 319416
rect 309778 319404 309784 319456
rect 309836 319444 309842 319456
rect 309962 319444 309968 319456
rect 309836 319416 309968 319444
rect 309836 319404 309842 319416
rect 309962 319404 309968 319416
rect 310020 319404 310026 319456
rect 311866 319444 311894 319484
rect 312814 319472 312820 319524
rect 312872 319512 312878 319524
rect 317432 319512 317460 319552
rect 321554 319540 321560 319592
rect 321612 319540 321618 319592
rect 321646 319540 321652 319592
rect 321704 319580 321710 319592
rect 322584 319580 322612 319756
rect 322814 319728 322842 319880
rect 323486 319812 323492 319864
rect 323544 319812 323550 319864
rect 322750 319676 322756 319728
rect 322808 319688 322842 319728
rect 322808 319676 322814 319688
rect 323394 319676 323400 319728
rect 323452 319716 323458 319728
rect 323504 319716 323532 319812
rect 323452 319688 323532 319716
rect 323452 319676 323458 319688
rect 323854 319676 323860 319728
rect 323912 319716 323918 319728
rect 324010 319716 324038 319880
rect 324102 319852 324130 319960
rect 325114 319932 325142 320028
rect 327626 320016 327632 320028
rect 327684 320016 327690 320068
rect 329926 319988 329932 320000
rect 325206 319960 329932 319988
rect 325096 319880 325102 319932
rect 325154 319880 325160 319932
rect 325206 319852 325234 319960
rect 329926 319948 329932 319960
rect 329984 319948 329990 320000
rect 326660 319880 326666 319932
rect 326718 319880 326724 319932
rect 327120 319880 327126 319932
rect 327178 319920 327184 319932
rect 327626 319920 327632 319932
rect 327178 319892 327632 319920
rect 327178 319880 327184 319892
rect 327626 319880 327632 319892
rect 327684 319880 327690 319932
rect 324102 319824 325234 319852
rect 325280 319812 325286 319864
rect 325338 319812 325344 319864
rect 323912 319688 324038 319716
rect 323912 319676 323918 319688
rect 325050 319676 325056 319728
rect 325108 319716 325114 319728
rect 325298 319716 325326 319812
rect 326430 319744 326436 319796
rect 326488 319744 326494 319796
rect 325108 319688 325326 319716
rect 325108 319676 325114 319688
rect 325694 319676 325700 319728
rect 325752 319716 325758 319728
rect 326448 319716 326476 319744
rect 326678 319728 326706 319880
rect 326752 319812 326758 319864
rect 326810 319812 326816 319864
rect 326770 319784 326798 319812
rect 327074 319784 327080 319796
rect 326770 319756 327080 319784
rect 327074 319744 327080 319756
rect 327132 319744 327138 319796
rect 327166 319744 327172 319796
rect 327224 319784 327230 319796
rect 335354 319784 335360 319796
rect 327224 319756 335360 319784
rect 327224 319744 327230 319756
rect 335354 319744 335360 319756
rect 335412 319744 335418 319796
rect 325752 319688 326476 319716
rect 325752 319676 325758 319688
rect 326614 319676 326620 319728
rect 326672 319688 326706 319728
rect 326672 319676 326678 319688
rect 326798 319676 326804 319728
rect 326856 319716 326862 319728
rect 332318 319716 332324 319728
rect 326856 319688 332324 319716
rect 326856 319676 326862 319688
rect 332318 319676 332324 319688
rect 332376 319676 332382 319728
rect 323486 319608 323492 319660
rect 323544 319648 323550 319660
rect 354858 319648 354864 319660
rect 323544 319620 354864 319648
rect 323544 319608 323550 319620
rect 354858 319608 354864 319620
rect 354916 319608 354922 319660
rect 343358 319580 343364 319592
rect 321704 319552 322612 319580
rect 323964 319552 343364 319580
rect 321704 319540 321710 319552
rect 312872 319484 317460 319512
rect 312872 319472 312878 319484
rect 318058 319472 318064 319524
rect 318116 319512 318122 319524
rect 318242 319512 318248 319524
rect 318116 319484 318248 319512
rect 318116 319472 318122 319484
rect 318242 319472 318248 319484
rect 318300 319472 318306 319524
rect 318334 319472 318340 319524
rect 318392 319512 318398 319524
rect 323964 319512 323992 319552
rect 343358 319540 343364 319552
rect 343416 319540 343422 319592
rect 318392 319484 323992 319512
rect 318392 319472 318398 319484
rect 326338 319472 326344 319524
rect 326396 319512 326402 319524
rect 327166 319512 327172 319524
rect 326396 319484 327172 319512
rect 326396 319472 326402 319484
rect 327166 319472 327172 319484
rect 327224 319472 327230 319524
rect 327350 319472 327356 319524
rect 327408 319512 327414 319524
rect 361758 319512 361764 319524
rect 327408 319484 361764 319512
rect 327408 319472 327414 319484
rect 361758 319472 361764 319484
rect 361816 319472 361822 319524
rect 323486 319444 323492 319456
rect 311866 319416 323492 319444
rect 323486 319404 323492 319416
rect 323544 319404 323550 319456
rect 325050 319404 325056 319456
rect 325108 319444 325114 319456
rect 325326 319444 325332 319456
rect 325108 319416 325332 319444
rect 325108 319404 325114 319416
rect 325326 319404 325332 319416
rect 325384 319404 325390 319456
rect 329926 319404 329932 319456
rect 329984 319444 329990 319456
rect 330110 319444 330116 319456
rect 329984 319416 330116 319444
rect 329984 319404 329990 319416
rect 330110 319404 330116 319416
rect 330168 319444 330174 319456
rect 371694 319444 371700 319456
rect 330168 319416 371700 319444
rect 330168 319404 330174 319416
rect 371694 319404 371700 319416
rect 371752 319404 371758 319456
rect 282914 319336 282920 319388
rect 282972 319376 282978 319388
rect 283098 319376 283104 319388
rect 282972 319348 283104 319376
rect 282972 319336 282978 319348
rect 283098 319336 283104 319348
rect 283156 319336 283162 319388
rect 283374 319336 283380 319388
rect 283432 319376 283438 319388
rect 283558 319376 283564 319388
rect 283432 319348 283564 319376
rect 283432 319336 283438 319348
rect 283558 319336 283564 319348
rect 283616 319336 283622 319388
rect 285214 319336 285220 319388
rect 285272 319376 285278 319388
rect 285674 319376 285680 319388
rect 285272 319348 285680 319376
rect 285272 319336 285278 319348
rect 285674 319336 285680 319348
rect 285732 319336 285738 319388
rect 287514 319336 287520 319388
rect 287572 319376 287578 319388
rect 287974 319376 287980 319388
rect 287572 319348 287980 319376
rect 287572 319336 287578 319348
rect 287974 319336 287980 319348
rect 288032 319336 288038 319388
rect 288894 319336 288900 319388
rect 288952 319376 288958 319388
rect 289814 319376 289820 319388
rect 288952 319348 289820 319376
rect 288952 319336 288958 319348
rect 289814 319336 289820 319348
rect 289872 319336 289878 319388
rect 291286 319336 291292 319388
rect 291344 319376 291350 319388
rect 292022 319376 292028 319388
rect 291344 319348 292028 319376
rect 291344 319336 291350 319348
rect 292022 319336 292028 319348
rect 292080 319336 292086 319388
rect 345934 319376 345940 319388
rect 292546 319348 345940 319376
rect 206646 319268 206652 319320
rect 206704 319308 206710 319320
rect 206704 319280 284432 319308
rect 206704 319268 206710 319280
rect 276474 319200 276480 319252
rect 276532 319240 276538 319252
rect 279970 319240 279976 319252
rect 276532 319212 279976 319240
rect 276532 319200 276538 319212
rect 279970 319200 279976 319212
rect 280028 319200 280034 319252
rect 278314 319132 278320 319184
rect 278372 319172 278378 319184
rect 280062 319172 280068 319184
rect 278372 319144 280068 319172
rect 278372 319132 278378 319144
rect 280062 319132 280068 319144
rect 280120 319132 280126 319184
rect 258258 319104 258264 319116
rect 200086 319076 258264 319104
rect 3418 318792 3424 318844
rect 3476 318832 3482 318844
rect 197354 318832 197360 318844
rect 3476 318804 197360 318832
rect 3476 318792 3482 318804
rect 197354 318792 197360 318804
rect 197412 318832 197418 318844
rect 200086 318832 200114 319076
rect 258258 319064 258264 319076
rect 258316 319104 258322 319116
rect 258810 319104 258816 319116
rect 258316 319076 258816 319104
rect 258316 319064 258322 319076
rect 258810 319064 258816 319076
rect 258868 319064 258874 319116
rect 275922 319064 275928 319116
rect 275980 319104 275986 319116
rect 283098 319104 283104 319116
rect 275980 319076 283104 319104
rect 275980 319064 275986 319076
rect 283098 319064 283104 319076
rect 283156 319064 283162 319116
rect 284404 319104 284432 319280
rect 285030 319268 285036 319320
rect 285088 319308 285094 319320
rect 285582 319308 285588 319320
rect 285088 319280 285588 319308
rect 285088 319268 285094 319280
rect 285582 319268 285588 319280
rect 285640 319268 285646 319320
rect 289998 319268 290004 319320
rect 290056 319308 290062 319320
rect 290366 319308 290372 319320
rect 290056 319280 290372 319308
rect 290056 319268 290062 319280
rect 290366 319268 290372 319280
rect 290424 319308 290430 319320
rect 292546 319308 292574 319348
rect 345934 319336 345940 319348
rect 345992 319336 345998 319388
rect 290424 319280 292574 319308
rect 290424 319268 290430 319280
rect 292758 319268 292764 319320
rect 292816 319308 292822 319320
rect 352926 319308 352932 319320
rect 292816 319280 352932 319308
rect 292816 319268 292822 319280
rect 352926 319268 352932 319280
rect 352984 319268 352990 319320
rect 284478 319200 284484 319252
rect 284536 319240 284542 319252
rect 343910 319240 343916 319252
rect 284536 319212 343916 319240
rect 284536 319200 284542 319212
rect 343910 319200 343916 319212
rect 343968 319200 343974 319252
rect 287146 319132 287152 319184
rect 287204 319172 287210 319184
rect 346486 319172 346492 319184
rect 287204 319144 346492 319172
rect 287204 319132 287210 319144
rect 346486 319132 346492 319144
rect 346544 319132 346550 319184
rect 288986 319104 288992 319116
rect 284404 319076 288992 319104
rect 288986 319064 288992 319076
rect 289044 319104 289050 319116
rect 347958 319104 347964 319116
rect 289044 319076 347964 319104
rect 289044 319064 289050 319076
rect 347958 319064 347964 319076
rect 348016 319064 348022 319116
rect 224310 318996 224316 319048
rect 224368 319036 224374 319048
rect 292758 319036 292764 319048
rect 224368 319008 292764 319036
rect 224368 318996 224374 319008
rect 292758 318996 292764 319008
rect 292816 318996 292822 319048
rect 292942 318996 292948 319048
rect 293000 319036 293006 319048
rect 294414 319036 294420 319048
rect 293000 319008 294420 319036
rect 293000 318996 293006 319008
rect 294414 318996 294420 319008
rect 294472 318996 294478 319048
rect 294782 318996 294788 319048
rect 294840 319036 294846 319048
rect 298554 319036 298560 319048
rect 294840 319008 298560 319036
rect 294840 318996 294846 319008
rect 298554 318996 298560 319008
rect 298612 318996 298618 319048
rect 301130 318996 301136 319048
rect 301188 319036 301194 319048
rect 301682 319036 301688 319048
rect 301188 319008 301688 319036
rect 301188 318996 301194 319008
rect 301682 318996 301688 319008
rect 301740 318996 301746 319048
rect 302510 318996 302516 319048
rect 302568 319036 302574 319048
rect 303154 319036 303160 319048
rect 302568 319008 303160 319036
rect 302568 318996 302574 319008
rect 303154 318996 303160 319008
rect 303212 318996 303218 319048
rect 303706 318996 303712 319048
rect 303764 319036 303770 319048
rect 352466 319036 352472 319048
rect 303764 319008 352472 319036
rect 303764 318996 303770 319008
rect 352466 318996 352472 319008
rect 352524 318996 352530 319048
rect 208210 318928 208216 318980
rect 208268 318968 208274 318980
rect 286962 318968 286968 318980
rect 208268 318940 286968 318968
rect 208268 318928 208274 318940
rect 286962 318928 286968 318940
rect 287020 318968 287026 318980
rect 346578 318968 346584 318980
rect 287020 318940 296484 318968
rect 287020 318928 287026 318940
rect 206554 318860 206560 318912
rect 206612 318900 206618 318912
rect 278038 318900 278044 318912
rect 206612 318872 278044 318900
rect 206612 318860 206618 318872
rect 278038 318860 278044 318872
rect 278096 318860 278102 318912
rect 279510 318860 279516 318912
rect 279568 318900 279574 318912
rect 295978 318900 295984 318912
rect 279568 318872 295984 318900
rect 279568 318860 279574 318872
rect 295978 318860 295984 318872
rect 296036 318860 296042 318912
rect 296456 318900 296484 318940
rect 296640 318940 346584 318968
rect 296640 318900 296668 318940
rect 346578 318928 346584 318940
rect 346636 318928 346642 318980
rect 296456 318872 296668 318900
rect 313458 318860 313464 318912
rect 313516 318900 313522 318912
rect 314562 318900 314568 318912
rect 313516 318872 314568 318900
rect 313516 318860 313522 318872
rect 314562 318860 314568 318872
rect 314620 318860 314626 318912
rect 317966 318860 317972 318912
rect 318024 318900 318030 318912
rect 318334 318900 318340 318912
rect 318024 318872 318340 318900
rect 318024 318860 318030 318872
rect 318334 318860 318340 318872
rect 318392 318860 318398 318912
rect 319530 318860 319536 318912
rect 319588 318900 319594 318912
rect 319714 318900 319720 318912
rect 319588 318872 319720 318900
rect 319588 318860 319594 318872
rect 319714 318860 319720 318872
rect 319772 318860 319778 318912
rect 320082 318860 320088 318912
rect 320140 318900 320146 318912
rect 379054 318900 379060 318912
rect 320140 318872 379060 318900
rect 320140 318860 320146 318872
rect 379054 318860 379060 318872
rect 379112 318860 379118 318912
rect 197412 318804 200114 318832
rect 197412 318792 197418 318804
rect 275554 318792 275560 318844
rect 275612 318832 275618 318844
rect 276842 318832 276848 318844
rect 275612 318804 276848 318832
rect 275612 318792 275618 318804
rect 276842 318792 276848 318804
rect 276900 318792 276906 318844
rect 277670 318792 277676 318844
rect 277728 318832 277734 318844
rect 278498 318832 278504 318844
rect 277728 318804 278504 318832
rect 277728 318792 277734 318804
rect 278498 318792 278504 318804
rect 278556 318792 278562 318844
rect 279786 318792 279792 318844
rect 279844 318832 279850 318844
rect 281442 318832 281448 318844
rect 279844 318804 281448 318832
rect 279844 318792 279850 318804
rect 281442 318792 281448 318804
rect 281500 318832 281506 318844
rect 281902 318832 281908 318844
rect 281500 318804 281908 318832
rect 281500 318792 281506 318804
rect 281902 318792 281908 318804
rect 281960 318792 281966 318844
rect 282178 318792 282184 318844
rect 282236 318832 282242 318844
rect 292942 318832 292948 318844
rect 282236 318804 292948 318832
rect 282236 318792 282242 318804
rect 292942 318792 292948 318804
rect 293000 318792 293006 318844
rect 293586 318792 293592 318844
rect 293644 318832 293650 318844
rect 303706 318832 303712 318844
rect 293644 318804 303712 318832
rect 293644 318792 293650 318804
rect 303706 318792 303712 318804
rect 303764 318792 303770 318844
rect 320174 318792 320180 318844
rect 320232 318832 320238 318844
rect 322934 318832 322940 318844
rect 320232 318804 322940 318832
rect 320232 318792 320238 318804
rect 322934 318792 322940 318804
rect 322992 318792 322998 318844
rect 325418 318792 325424 318844
rect 325476 318832 325482 318844
rect 327350 318832 327356 318844
rect 325476 318804 327356 318832
rect 325476 318792 325482 318804
rect 327350 318792 327356 318804
rect 327408 318792 327414 318844
rect 335354 318792 335360 318844
rect 335412 318832 335418 318844
rect 336458 318832 336464 318844
rect 335412 318804 336464 318832
rect 335412 318792 335418 318804
rect 336458 318792 336464 318804
rect 336516 318792 336522 318844
rect 282086 318724 282092 318776
rect 282144 318764 282150 318776
rect 282454 318764 282460 318776
rect 282144 318736 282460 318764
rect 282144 318724 282150 318736
rect 282454 318724 282460 318736
rect 282512 318764 282518 318776
rect 285306 318764 285312 318776
rect 282512 318736 285312 318764
rect 282512 318724 282518 318736
rect 285306 318724 285312 318736
rect 285364 318724 285370 318776
rect 291654 318724 291660 318776
rect 291712 318764 291718 318776
rect 291930 318764 291936 318776
rect 291712 318736 291936 318764
rect 291712 318724 291718 318736
rect 291930 318724 291936 318736
rect 291988 318724 291994 318776
rect 295978 318724 295984 318776
rect 296036 318764 296042 318776
rect 296438 318764 296444 318776
rect 296036 318736 296444 318764
rect 296036 318724 296042 318736
rect 296438 318724 296444 318736
rect 296496 318724 296502 318776
rect 297266 318724 297272 318776
rect 297324 318764 297330 318776
rect 297450 318764 297456 318776
rect 297324 318736 297456 318764
rect 297324 318724 297330 318736
rect 297450 318724 297456 318736
rect 297508 318724 297514 318776
rect 310974 318724 310980 318776
rect 311032 318764 311038 318776
rect 314562 318764 314568 318776
rect 311032 318736 314568 318764
rect 311032 318724 311038 318736
rect 314562 318724 314568 318736
rect 314620 318724 314626 318776
rect 317782 318724 317788 318776
rect 317840 318764 317846 318776
rect 322474 318764 322480 318776
rect 317840 318736 322480 318764
rect 317840 318724 317846 318736
rect 322474 318724 322480 318736
rect 322532 318724 322538 318776
rect 325878 318724 325884 318776
rect 325936 318764 325942 318776
rect 329650 318764 329656 318776
rect 325936 318736 329656 318764
rect 325936 318724 325942 318736
rect 329650 318724 329656 318736
rect 329708 318724 329714 318776
rect 331766 318724 331772 318776
rect 331824 318764 331830 318776
rect 357066 318764 357072 318776
rect 331824 318736 357072 318764
rect 331824 318724 331830 318736
rect 357066 318724 357072 318736
rect 357124 318724 357130 318776
rect 269298 318656 269304 318708
rect 269356 318696 269362 318708
rect 274082 318696 274088 318708
rect 269356 318668 274088 318696
rect 269356 318656 269362 318668
rect 274082 318656 274088 318668
rect 274140 318696 274146 318708
rect 288158 318696 288164 318708
rect 274140 318668 288164 318696
rect 274140 318656 274146 318668
rect 288158 318656 288164 318668
rect 288216 318656 288222 318708
rect 290458 318656 290464 318708
rect 290516 318696 290522 318708
rect 290516 318668 297404 318696
rect 290516 318656 290522 318668
rect 276934 318588 276940 318640
rect 276992 318628 276998 318640
rect 284202 318628 284208 318640
rect 276992 318600 284208 318628
rect 276992 318588 276998 318600
rect 284202 318588 284208 318600
rect 284260 318588 284266 318640
rect 290642 318588 290648 318640
rect 290700 318628 290706 318640
rect 290700 318600 292436 318628
rect 290700 318588 290706 318600
rect 270218 318520 270224 318572
rect 270276 318560 270282 318572
rect 278038 318560 278044 318572
rect 270276 318532 278044 318560
rect 270276 318520 270282 318532
rect 278038 318520 278044 318532
rect 278096 318520 278102 318572
rect 292298 318560 292304 318572
rect 287670 318532 292304 318560
rect 270034 318452 270040 318504
rect 270092 318492 270098 318504
rect 274450 318492 274456 318504
rect 270092 318464 274456 318492
rect 270092 318452 270098 318464
rect 274450 318452 274456 318464
rect 274508 318492 274514 318504
rect 287670 318492 287698 318532
rect 292298 318520 292304 318532
rect 292356 318520 292362 318572
rect 292408 318560 292436 318600
rect 297376 318560 297404 318668
rect 300854 318656 300860 318708
rect 300912 318696 300918 318708
rect 302418 318696 302424 318708
rect 300912 318668 302424 318696
rect 300912 318656 300918 318668
rect 302418 318656 302424 318668
rect 302476 318656 302482 318708
rect 324774 318656 324780 318708
rect 324832 318696 324838 318708
rect 329558 318696 329564 318708
rect 324832 318668 329564 318696
rect 324832 318656 324838 318668
rect 329558 318656 329564 318668
rect 329616 318656 329622 318708
rect 298094 318588 298100 318640
rect 298152 318628 298158 318640
rect 303982 318628 303988 318640
rect 298152 318600 303988 318628
rect 298152 318588 298158 318600
rect 303982 318588 303988 318600
rect 304040 318588 304046 318640
rect 314746 318588 314752 318640
rect 314804 318628 314810 318640
rect 329466 318628 329472 318640
rect 314804 318600 329472 318628
rect 314804 318588 314810 318600
rect 329466 318588 329472 318600
rect 329524 318588 329530 318640
rect 332226 318560 332232 318572
rect 292408 318532 292574 318560
rect 297376 318532 332232 318560
rect 274508 318464 287698 318492
rect 274508 318452 274514 318464
rect 290366 318452 290372 318504
rect 290424 318492 290430 318504
rect 290642 318492 290648 318504
rect 290424 318464 290648 318492
rect 290424 318452 290430 318464
rect 290642 318452 290648 318464
rect 290700 318452 290706 318504
rect 291746 318452 291752 318504
rect 291804 318492 291810 318504
rect 291930 318492 291936 318504
rect 291804 318464 291936 318492
rect 291804 318452 291810 318464
rect 291930 318452 291936 318464
rect 291988 318452 291994 318504
rect 292546 318492 292574 318532
rect 332226 318520 332232 318532
rect 332284 318520 332290 318572
rect 297726 318492 297732 318504
rect 292546 318464 297732 318492
rect 297726 318452 297732 318464
rect 297784 318452 297790 318504
rect 301498 318452 301504 318504
rect 301556 318492 301562 318504
rect 302694 318492 302700 318504
rect 301556 318464 302700 318492
rect 301556 318452 301562 318464
rect 302694 318452 302700 318464
rect 302752 318452 302758 318504
rect 303982 318452 303988 318504
rect 304040 318492 304046 318504
rect 304626 318492 304632 318504
rect 304040 318464 304632 318492
rect 304040 318452 304046 318464
rect 304626 318452 304632 318464
rect 304684 318452 304690 318504
rect 309502 318452 309508 318504
rect 309560 318492 309566 318504
rect 310238 318492 310244 318504
rect 309560 318464 310244 318492
rect 309560 318452 309566 318464
rect 310238 318452 310244 318464
rect 310296 318452 310302 318504
rect 317690 318452 317696 318504
rect 317748 318492 317754 318504
rect 324774 318492 324780 318504
rect 317748 318464 324780 318492
rect 317748 318452 317754 318464
rect 324774 318452 324780 318464
rect 324832 318452 324838 318504
rect 269390 318384 269396 318436
rect 269448 318424 269454 318436
rect 269942 318424 269948 318436
rect 269448 318396 269948 318424
rect 269448 318384 269454 318396
rect 269942 318384 269948 318396
rect 270000 318384 270006 318436
rect 270310 318384 270316 318436
rect 270368 318424 270374 318436
rect 284754 318424 284760 318436
rect 270368 318396 284760 318424
rect 270368 318384 270374 318396
rect 284754 318384 284760 318396
rect 284812 318384 284818 318436
rect 295886 318424 295892 318436
rect 290016 318396 295892 318424
rect 271690 318316 271696 318368
rect 271748 318356 271754 318368
rect 286134 318356 286140 318368
rect 271748 318328 286140 318356
rect 271748 318316 271754 318328
rect 286134 318316 286140 318328
rect 286192 318316 286198 318368
rect 242526 318248 242532 318300
rect 242584 318288 242590 318300
rect 242584 318260 273254 318288
rect 242584 318248 242590 318260
rect 273226 318220 273254 318260
rect 278038 318248 278044 318300
rect 278096 318288 278102 318300
rect 288066 318288 288072 318300
rect 278096 318260 288072 318288
rect 278096 318248 278102 318260
rect 288066 318248 288072 318260
rect 288124 318248 288130 318300
rect 281534 318220 281540 318232
rect 273226 318192 281540 318220
rect 281534 318180 281540 318192
rect 281592 318220 281598 318232
rect 282730 318220 282736 318232
rect 281592 318192 282736 318220
rect 281592 318180 281598 318192
rect 282730 318180 282736 318192
rect 282788 318180 282794 318232
rect 289906 318220 289912 318232
rect 282886 318192 289912 318220
rect 238754 318112 238760 318164
rect 238812 318152 238818 318164
rect 238812 318124 273254 318152
rect 238812 318112 238818 318124
rect 213822 318044 213828 318096
rect 213880 318084 213886 318096
rect 271322 318084 271328 318096
rect 213880 318056 271328 318084
rect 213880 318044 213886 318056
rect 271322 318044 271328 318056
rect 271380 318084 271386 318096
rect 271690 318084 271696 318096
rect 271380 318056 271696 318084
rect 271380 318044 271386 318056
rect 271690 318044 271696 318056
rect 271748 318044 271754 318096
rect 273226 318084 273254 318124
rect 281626 318112 281632 318164
rect 281684 318152 281690 318164
rect 282886 318152 282914 318192
rect 289906 318180 289912 318192
rect 289964 318180 289970 318232
rect 281684 318124 282914 318152
rect 281684 318112 281690 318124
rect 282270 318084 282276 318096
rect 273226 318056 282276 318084
rect 282270 318044 282276 318056
rect 282328 318044 282334 318096
rect 275830 317976 275836 318028
rect 275888 318016 275894 318028
rect 290016 318016 290044 318396
rect 295886 318384 295892 318396
rect 295944 318384 295950 318436
rect 296438 318384 296444 318436
rect 296496 318424 296502 318436
rect 297174 318424 297180 318436
rect 296496 318396 297180 318424
rect 296496 318384 296502 318396
rect 297174 318384 297180 318396
rect 297232 318384 297238 318436
rect 333514 318424 333520 318436
rect 297376 318396 333520 318424
rect 291286 318316 291292 318368
rect 291344 318356 291350 318368
rect 291746 318356 291752 318368
rect 291344 318328 291752 318356
rect 291344 318316 291350 318328
rect 291746 318316 291752 318328
rect 291804 318356 291810 318368
rect 297376 318356 297404 318396
rect 333514 318384 333520 318396
rect 333572 318384 333578 318436
rect 332042 318356 332048 318368
rect 291804 318328 297404 318356
rect 297468 318328 332048 318356
rect 291804 318316 291810 318328
rect 291470 318248 291476 318300
rect 291528 318288 291534 318300
rect 292482 318288 292488 318300
rect 291528 318260 292488 318288
rect 291528 318248 291534 318260
rect 292482 318248 292488 318260
rect 292540 318288 292546 318300
rect 297468 318288 297496 318328
rect 332042 318316 332048 318328
rect 332100 318316 332106 318368
rect 292540 318260 297496 318288
rect 292540 318248 292546 318260
rect 297726 318248 297732 318300
rect 297784 318288 297790 318300
rect 328086 318288 328092 318300
rect 297784 318260 328092 318288
rect 297784 318248 297790 318260
rect 328086 318248 328092 318260
rect 328144 318248 328150 318300
rect 328730 318248 328736 318300
rect 328788 318288 328794 318300
rect 359458 318288 359464 318300
rect 328788 318260 359464 318288
rect 328788 318248 328794 318260
rect 359458 318248 359464 318260
rect 359516 318248 359522 318300
rect 315022 318180 315028 318232
rect 315080 318220 315086 318232
rect 328178 318220 328184 318232
rect 315080 318192 328184 318220
rect 315080 318180 315086 318192
rect 328178 318180 328184 318192
rect 328236 318180 328242 318232
rect 328822 318180 328828 318232
rect 328880 318220 328886 318232
rect 360930 318220 360936 318232
rect 328880 318192 360936 318220
rect 328880 318180 328886 318192
rect 360930 318180 360936 318192
rect 360988 318180 360994 318232
rect 290550 318112 290556 318164
rect 290608 318152 290614 318164
rect 291102 318152 291108 318164
rect 290608 318124 291108 318152
rect 290608 318112 290614 318124
rect 291102 318112 291108 318124
rect 291160 318152 291166 318164
rect 297266 318152 297272 318164
rect 291160 318124 297272 318152
rect 291160 318112 291166 318124
rect 297266 318112 297272 318124
rect 297324 318112 297330 318164
rect 299290 318112 299296 318164
rect 299348 318152 299354 318164
rect 300486 318152 300492 318164
rect 299348 318124 300492 318152
rect 299348 318112 299354 318124
rect 300486 318112 300492 318124
rect 300544 318112 300550 318164
rect 304626 318112 304632 318164
rect 304684 318152 304690 318164
rect 304902 318152 304908 318164
rect 304684 318124 304908 318152
rect 304684 318112 304690 318124
rect 304902 318112 304908 318124
rect 304960 318112 304966 318164
rect 309870 318112 309876 318164
rect 309928 318152 309934 318164
rect 310146 318152 310152 318164
rect 309928 318124 310152 318152
rect 309928 318112 309934 318124
rect 310146 318112 310152 318124
rect 310204 318112 310210 318164
rect 322290 318112 322296 318164
rect 322348 318152 322354 318164
rect 324038 318152 324044 318164
rect 322348 318124 324044 318152
rect 322348 318112 322354 318124
rect 324038 318112 324044 318124
rect 324096 318112 324102 318164
rect 328638 318112 328644 318164
rect 328696 318152 328702 318164
rect 364518 318152 364524 318164
rect 328696 318124 364524 318152
rect 328696 318112 328702 318124
rect 364518 318112 364524 318124
rect 364576 318112 364582 318164
rect 292114 318044 292120 318096
rect 292172 318084 292178 318096
rect 292574 318084 292580 318096
rect 292172 318056 292580 318084
rect 292172 318044 292178 318056
rect 292574 318044 292580 318056
rect 292632 318084 292638 318096
rect 317506 318084 317512 318096
rect 292632 318056 317512 318084
rect 292632 318044 292638 318056
rect 317506 318044 317512 318056
rect 317564 318044 317570 318096
rect 323118 318044 323124 318096
rect 323176 318084 323182 318096
rect 331398 318084 331404 318096
rect 323176 318056 331404 318084
rect 323176 318044 323182 318056
rect 331398 318044 331404 318056
rect 331456 318084 331462 318096
rect 331766 318084 331772 318096
rect 331456 318056 331772 318084
rect 331456 318044 331462 318056
rect 331766 318044 331772 318056
rect 331824 318044 331830 318096
rect 332318 318044 332324 318096
rect 332376 318084 332382 318096
rect 388254 318084 388260 318096
rect 332376 318056 388260 318084
rect 332376 318044 332382 318056
rect 388254 318044 388260 318056
rect 388312 318044 388318 318096
rect 275888 317988 290044 318016
rect 275888 317976 275894 317988
rect 303154 317976 303160 318028
rect 303212 318016 303218 318028
rect 304994 318016 305000 318028
rect 303212 317988 305000 318016
rect 303212 317976 303218 317988
rect 304994 317976 305000 317988
rect 305052 317976 305058 318028
rect 328454 317976 328460 318028
rect 328512 318016 328518 318028
rect 354214 318016 354220 318028
rect 328512 317988 354220 318016
rect 328512 317976 328518 317988
rect 354214 317976 354220 317988
rect 354272 317976 354278 318028
rect 259178 317908 259184 317960
rect 259236 317948 259242 317960
rect 288526 317948 288532 317960
rect 259236 317920 288532 317948
rect 259236 317908 259242 317920
rect 288526 317908 288532 317920
rect 288584 317908 288590 317960
rect 294506 317908 294512 317960
rect 294564 317948 294570 317960
rect 295058 317948 295064 317960
rect 294564 317920 295064 317948
rect 294564 317908 294570 317920
rect 295058 317908 295064 317920
rect 295116 317908 295122 317960
rect 302602 317908 302608 317960
rect 302660 317948 302666 317960
rect 307386 317948 307392 317960
rect 302660 317920 307392 317948
rect 302660 317908 302666 317920
rect 307386 317908 307392 317920
rect 307444 317908 307450 317960
rect 309870 317908 309876 317960
rect 309928 317948 309934 317960
rect 310422 317948 310428 317960
rect 309928 317920 310428 317948
rect 309928 317908 309934 317920
rect 310422 317908 310428 317920
rect 310480 317908 310486 317960
rect 325694 317908 325700 317960
rect 325752 317948 325758 317960
rect 326982 317948 326988 317960
rect 325752 317920 326988 317948
rect 325752 317908 325758 317920
rect 326982 317908 326988 317920
rect 327040 317908 327046 317960
rect 328546 317908 328552 317960
rect 328604 317948 328610 317960
rect 338574 317948 338580 317960
rect 328604 317920 338580 317948
rect 328604 317908 328610 317920
rect 338574 317908 338580 317920
rect 338632 317908 338638 317960
rect 268562 317840 268568 317892
rect 268620 317880 268626 317892
rect 282914 317880 282920 317892
rect 268620 317852 282920 317880
rect 268620 317840 268626 317852
rect 282914 317840 282920 317852
rect 282972 317840 282978 317892
rect 286042 317840 286048 317892
rect 286100 317880 286106 317892
rect 331122 317880 331128 317892
rect 286100 317852 331128 317880
rect 286100 317840 286106 317852
rect 331122 317840 331128 317852
rect 331180 317840 331186 317892
rect 298094 317812 298100 317824
rect 276676 317784 298100 317812
rect 276676 317756 276704 317784
rect 298094 317772 298100 317784
rect 298152 317772 298158 317824
rect 302602 317772 302608 317824
rect 302660 317812 302666 317824
rect 303430 317812 303436 317824
rect 302660 317784 303436 317812
rect 302660 317772 302666 317784
rect 303430 317772 303436 317784
rect 303488 317772 303494 317824
rect 303706 317772 303712 317824
rect 303764 317812 303770 317824
rect 305362 317812 305368 317824
rect 303764 317784 305368 317812
rect 303764 317772 303770 317784
rect 305362 317772 305368 317784
rect 305420 317772 305426 317824
rect 306834 317772 306840 317824
rect 306892 317812 306898 317824
rect 318058 317812 318064 317824
rect 306892 317784 318064 317812
rect 306892 317772 306898 317784
rect 318058 317772 318064 317784
rect 318116 317772 318122 317824
rect 327166 317772 327172 317824
rect 327224 317812 327230 317824
rect 327442 317812 327448 317824
rect 327224 317784 327448 317812
rect 327224 317772 327230 317784
rect 327442 317772 327448 317784
rect 327500 317772 327506 317824
rect 275462 317704 275468 317756
rect 275520 317744 275526 317756
rect 276658 317744 276664 317756
rect 275520 317716 276664 317744
rect 275520 317704 275526 317716
rect 276658 317704 276664 317716
rect 276716 317704 276722 317756
rect 282914 317704 282920 317756
rect 282972 317744 282978 317756
rect 283098 317744 283104 317756
rect 282972 317716 283104 317744
rect 282972 317704 282978 317716
rect 283098 317704 283104 317716
rect 283156 317704 283162 317756
rect 286042 317744 286048 317756
rect 284036 317716 286048 317744
rect 249794 317636 249800 317688
rect 249852 317676 249858 317688
rect 284036 317676 284064 317716
rect 286042 317704 286048 317716
rect 286100 317704 286106 317756
rect 287330 317704 287336 317756
rect 287388 317744 287394 317756
rect 288250 317744 288256 317756
rect 287388 317716 288256 317744
rect 287388 317704 287394 317716
rect 288250 317704 288256 317716
rect 288308 317704 288314 317756
rect 334986 317744 334992 317756
rect 292546 317716 334992 317744
rect 249852 317648 284064 317676
rect 249852 317636 249858 317648
rect 284110 317636 284116 317688
rect 284168 317676 284174 317688
rect 290182 317676 290188 317688
rect 284168 317648 290188 317676
rect 284168 317636 284174 317648
rect 290182 317636 290188 317648
rect 290240 317636 290246 317688
rect 290274 317636 290280 317688
rect 290332 317676 290338 317688
rect 291102 317676 291108 317688
rect 290332 317648 291108 317676
rect 290332 317636 290338 317648
rect 291102 317636 291108 317648
rect 291160 317636 291166 317688
rect 291194 317636 291200 317688
rect 291252 317676 291258 317688
rect 292298 317676 292304 317688
rect 291252 317648 292304 317676
rect 291252 317636 291258 317648
rect 292298 317636 292304 317648
rect 292356 317676 292362 317688
rect 292546 317676 292574 317716
rect 334986 317704 334992 317716
rect 335044 317704 335050 317756
rect 292356 317648 292574 317676
rect 292356 317636 292362 317648
rect 293494 317636 293500 317688
rect 293552 317676 293558 317688
rect 294230 317676 294236 317688
rect 293552 317648 294236 317676
rect 293552 317636 293558 317648
rect 294230 317636 294236 317648
rect 294288 317636 294294 317688
rect 297266 317636 297272 317688
rect 297324 317676 297330 317688
rect 332502 317676 332508 317688
rect 297324 317648 332508 317676
rect 297324 317636 297330 317648
rect 332502 317636 332508 317648
rect 332560 317636 332566 317688
rect 269390 317568 269396 317620
rect 269448 317608 269454 317620
rect 293678 317608 293684 317620
rect 269448 317580 293684 317608
rect 269448 317568 269454 317580
rect 293678 317568 293684 317580
rect 293736 317568 293742 317620
rect 295058 317568 295064 317620
rect 295116 317608 295122 317620
rect 296622 317608 296628 317620
rect 295116 317580 296628 317608
rect 295116 317568 295122 317580
rect 296622 317568 296628 317580
rect 296680 317568 296686 317620
rect 296714 317568 296720 317620
rect 296772 317608 296778 317620
rect 298278 317608 298284 317620
rect 296772 317580 298284 317608
rect 296772 317568 296778 317580
rect 298278 317568 298284 317580
rect 298336 317568 298342 317620
rect 303430 317568 303436 317620
rect 303488 317608 303494 317620
rect 304810 317608 304816 317620
rect 303488 317580 304816 317608
rect 303488 317568 303494 317580
rect 304810 317568 304816 317580
rect 304868 317568 304874 317620
rect 304902 317568 304908 317620
rect 304960 317608 304966 317620
rect 306466 317608 306472 317620
rect 304960 317580 306472 317608
rect 304960 317568 304966 317580
rect 306466 317568 306472 317580
rect 306524 317568 306530 317620
rect 307386 317568 307392 317620
rect 307444 317608 307450 317620
rect 313642 317608 313648 317620
rect 307444 317580 313648 317608
rect 307444 317568 307450 317580
rect 313642 317568 313648 317580
rect 313700 317568 313706 317620
rect 313936 317580 316356 317608
rect 286318 317500 286324 317552
rect 286376 317540 286382 317552
rect 290826 317540 290832 317552
rect 286376 317512 290832 317540
rect 286376 317500 286382 317512
rect 290826 317500 290832 317512
rect 290884 317500 290890 317552
rect 291194 317500 291200 317552
rect 291252 317540 291258 317552
rect 291930 317540 291936 317552
rect 291252 317512 291936 317540
rect 291252 317500 291258 317512
rect 291930 317500 291936 317512
rect 291988 317540 291994 317552
rect 313936 317540 313964 317580
rect 291988 317512 313964 317540
rect 316328 317540 316356 317580
rect 320634 317568 320640 317620
rect 320692 317608 320698 317620
rect 324774 317608 324780 317620
rect 320692 317580 324780 317608
rect 320692 317568 320698 317580
rect 324774 317568 324780 317580
rect 324832 317568 324838 317620
rect 325326 317568 325332 317620
rect 325384 317608 325390 317620
rect 326982 317608 326988 317620
rect 325384 317580 326988 317608
rect 325384 317568 325390 317580
rect 326982 317568 326988 317580
rect 327040 317568 327046 317620
rect 333790 317540 333796 317552
rect 316328 317512 333796 317540
rect 291988 317500 291994 317512
rect 333790 317500 333796 317512
rect 333848 317500 333854 317552
rect 274542 317432 274548 317484
rect 274600 317472 274606 317484
rect 276934 317472 276940 317484
rect 274600 317444 276940 317472
rect 274600 317432 274606 317444
rect 276934 317432 276940 317444
rect 276992 317432 276998 317484
rect 287146 317432 287152 317484
rect 287204 317472 287210 317484
rect 291010 317472 291016 317484
rect 287204 317444 291016 317472
rect 287204 317432 287210 317444
rect 291010 317432 291016 317444
rect 291068 317432 291074 317484
rect 291102 317432 291108 317484
rect 291160 317472 291166 317484
rect 306834 317472 306840 317484
rect 291160 317444 306840 317472
rect 291160 317432 291166 317444
rect 306834 317432 306840 317444
rect 306892 317432 306898 317484
rect 309318 317432 309324 317484
rect 309376 317472 309382 317484
rect 310514 317472 310520 317484
rect 309376 317444 310520 317472
rect 309376 317432 309382 317444
rect 310514 317432 310520 317444
rect 310572 317432 310578 317484
rect 313642 317432 313648 317484
rect 313700 317472 313706 317484
rect 325418 317472 325424 317484
rect 313700 317444 325424 317472
rect 313700 317432 313706 317444
rect 325418 317432 325424 317444
rect 325476 317432 325482 317484
rect 327534 317432 327540 317484
rect 327592 317472 327598 317484
rect 328178 317472 328184 317484
rect 327592 317444 328184 317472
rect 327592 317432 327598 317444
rect 328178 317432 328184 317444
rect 328236 317432 328242 317484
rect 328362 317432 328368 317484
rect 328420 317472 328426 317484
rect 329558 317472 329564 317484
rect 328420 317444 329564 317472
rect 328420 317432 328426 317444
rect 329558 317432 329564 317444
rect 329616 317432 329622 317484
rect 280154 317364 280160 317416
rect 280212 317404 280218 317416
rect 280982 317404 280988 317416
rect 280212 317376 280988 317404
rect 280212 317364 280218 317376
rect 280982 317364 280988 317376
rect 281040 317404 281046 317416
rect 284938 317404 284944 317416
rect 281040 317376 284944 317404
rect 281040 317364 281046 317376
rect 284938 317364 284944 317376
rect 284996 317364 285002 317416
rect 289722 317364 289728 317416
rect 289780 317404 289786 317416
rect 290090 317404 290096 317416
rect 289780 317376 290096 317404
rect 289780 317364 289786 317376
rect 290090 317364 290096 317376
rect 290148 317364 290154 317416
rect 295334 317364 295340 317416
rect 295392 317404 295398 317416
rect 320358 317404 320364 317416
rect 295392 317376 320364 317404
rect 295392 317364 295398 317376
rect 320358 317364 320364 317376
rect 320416 317404 320422 317416
rect 331030 317404 331036 317416
rect 320416 317376 331036 317404
rect 320416 317364 320422 317376
rect 331030 317364 331036 317376
rect 331088 317364 331094 317416
rect 334986 317364 334992 317416
rect 335044 317404 335050 317416
rect 338666 317404 338672 317416
rect 335044 317376 338672 317404
rect 335044 317364 335050 317376
rect 338666 317364 338672 317376
rect 338724 317364 338730 317416
rect 280798 317296 280804 317348
rect 280856 317336 280862 317348
rect 297266 317336 297272 317348
rect 280856 317308 297272 317336
rect 280856 317296 280862 317308
rect 297266 317296 297272 317308
rect 297324 317296 297330 317348
rect 303246 317296 303252 317348
rect 303304 317336 303310 317348
rect 308214 317336 308220 317348
rect 303304 317308 308220 317336
rect 303304 317296 303310 317308
rect 308214 317296 308220 317308
rect 308272 317296 308278 317348
rect 316678 317296 316684 317348
rect 316736 317336 316742 317348
rect 332134 317336 332140 317348
rect 316736 317308 332140 317336
rect 316736 317296 316742 317308
rect 332134 317296 332140 317308
rect 332192 317296 332198 317348
rect 278682 317228 278688 317280
rect 278740 317268 278746 317280
rect 308398 317268 308404 317280
rect 278740 317240 308404 317268
rect 278740 317228 278746 317240
rect 308398 317228 308404 317240
rect 308456 317228 308462 317280
rect 315942 317228 315948 317280
rect 316000 317268 316006 317280
rect 375558 317268 375564 317280
rect 316000 317240 375564 317268
rect 316000 317228 316006 317240
rect 375558 317228 375564 317240
rect 375616 317268 375622 317280
rect 376662 317268 376668 317280
rect 375616 317240 376668 317268
rect 375616 317228 375622 317240
rect 376662 317228 376668 317240
rect 376720 317228 376726 317280
rect 265894 317160 265900 317212
rect 265952 317200 265958 317212
rect 286410 317200 286416 317212
rect 265952 317172 286416 317200
rect 265952 317160 265958 317172
rect 286410 317160 286416 317172
rect 286468 317160 286474 317212
rect 295610 317160 295616 317212
rect 295668 317200 295674 317212
rect 296346 317200 296352 317212
rect 295668 317172 296352 317200
rect 295668 317160 295674 317172
rect 296346 317160 296352 317172
rect 296404 317160 296410 317212
rect 296990 317160 296996 317212
rect 297048 317200 297054 317212
rect 330754 317200 330760 317212
rect 297048 317172 330760 317200
rect 297048 317160 297054 317172
rect 330754 317160 330760 317172
rect 330812 317160 330818 317212
rect 331674 317160 331680 317212
rect 331732 317200 331738 317212
rect 389634 317200 389640 317212
rect 331732 317172 389640 317200
rect 331732 317160 331738 317172
rect 389634 317160 389640 317172
rect 389692 317160 389698 317212
rect 283834 317132 283840 317144
rect 267706 317104 283840 317132
rect 209590 317024 209596 317076
rect 209648 317064 209654 317076
rect 266354 317064 266360 317076
rect 209648 317036 266360 317064
rect 209648 317024 209654 317036
rect 266354 317024 266360 317036
rect 266412 317024 266418 317076
rect 201310 316956 201316 317008
rect 201368 316996 201374 317008
rect 260650 316996 260656 317008
rect 201368 316968 260656 316996
rect 201368 316956 201374 316968
rect 260650 316956 260656 316968
rect 260708 316996 260714 317008
rect 267706 316996 267734 317104
rect 283834 317092 283840 317104
rect 283892 317092 283898 317144
rect 284294 317092 284300 317144
rect 284352 317132 284358 317144
rect 284478 317132 284484 317144
rect 284352 317104 284484 317132
rect 284352 317092 284358 317104
rect 284478 317092 284484 317104
rect 284536 317092 284542 317144
rect 295518 317092 295524 317144
rect 295576 317132 295582 317144
rect 350074 317132 350080 317144
rect 295576 317104 350080 317132
rect 295576 317092 295582 317104
rect 350074 317092 350080 317104
rect 350132 317092 350138 317144
rect 274450 317024 274456 317076
rect 274508 317064 274514 317076
rect 303798 317064 303804 317076
rect 274508 317036 303804 317064
rect 274508 317024 274514 317036
rect 303798 317024 303804 317036
rect 303856 317064 303862 317076
rect 328454 317064 328460 317076
rect 303856 317036 328460 317064
rect 303856 317024 303862 317036
rect 328454 317024 328460 317036
rect 328512 317024 328518 317076
rect 260708 316968 267734 316996
rect 260708 316956 260714 316968
rect 270954 316956 270960 317008
rect 271012 316996 271018 317008
rect 271012 316968 292574 316996
rect 271012 316956 271018 316968
rect 209038 316888 209044 316940
rect 209096 316928 209102 316940
rect 280154 316928 280160 316940
rect 209096 316900 280160 316928
rect 209096 316888 209102 316900
rect 280154 316888 280160 316900
rect 280212 316888 280218 316940
rect 292546 316928 292574 316968
rect 308214 316956 308220 317008
rect 308272 316996 308278 317008
rect 316678 316996 316684 317008
rect 308272 316968 316684 316996
rect 308272 316956 308278 316968
rect 316678 316956 316684 316968
rect 316736 316956 316742 317008
rect 317046 316956 317052 317008
rect 317104 316996 317110 317008
rect 328546 316996 328552 317008
rect 317104 316968 328552 316996
rect 317104 316956 317110 316968
rect 328546 316956 328552 316968
rect 328604 316956 328610 317008
rect 310698 316928 310704 316940
rect 292546 316900 310704 316928
rect 310698 316888 310704 316900
rect 310756 316928 310762 316940
rect 324038 316928 324044 316940
rect 310756 316900 324044 316928
rect 310756 316888 310762 316900
rect 324038 316888 324044 316900
rect 324096 316888 324102 316940
rect 219066 316820 219072 316872
rect 219124 316860 219130 316872
rect 294414 316860 294420 316872
rect 219124 316832 294420 316860
rect 219124 316820 219130 316832
rect 294414 316820 294420 316832
rect 294472 316820 294478 316872
rect 297266 316820 297272 316872
rect 297324 316860 297330 316872
rect 302234 316860 302240 316872
rect 297324 316832 302240 316860
rect 297324 316820 297330 316832
rect 302234 316820 302240 316832
rect 302292 316860 302298 316872
rect 303338 316860 303344 316872
rect 302292 316832 303344 316860
rect 302292 316820 302298 316832
rect 303338 316820 303344 316832
rect 303396 316820 303402 316872
rect 314562 316820 314568 316872
rect 314620 316860 314626 316872
rect 327258 316860 327264 316872
rect 314620 316832 327264 316860
rect 314620 316820 314626 316832
rect 327258 316820 327264 316832
rect 327316 316860 327322 316872
rect 341334 316860 341340 316872
rect 327316 316832 341340 316860
rect 327316 316820 327322 316832
rect 341334 316820 341340 316832
rect 341392 316820 341398 316872
rect 215110 316752 215116 316804
rect 215168 316792 215174 316804
rect 295518 316792 295524 316804
rect 215168 316764 295524 316792
rect 215168 316752 215174 316764
rect 295518 316752 295524 316764
rect 295576 316752 295582 316804
rect 317874 316752 317880 316804
rect 317932 316792 317938 316804
rect 345934 316792 345940 316804
rect 317932 316764 345940 316792
rect 317932 316752 317938 316764
rect 345934 316752 345940 316764
rect 345992 316792 345998 316804
rect 378042 316792 378048 316804
rect 345992 316764 378048 316792
rect 345992 316752 345998 316764
rect 378042 316752 378048 316764
rect 378100 316752 378106 316804
rect 295978 316684 295984 316736
rect 296036 316724 296042 316736
rect 309870 316724 309876 316736
rect 296036 316696 309876 316724
rect 296036 316684 296042 316696
rect 309870 316684 309876 316696
rect 309928 316724 309934 316736
rect 360194 316724 360200 316736
rect 309928 316696 360200 316724
rect 309928 316684 309934 316696
rect 360194 316684 360200 316696
rect 360252 316684 360258 316736
rect 376662 316684 376668 316736
rect 376720 316724 376726 316736
rect 429838 316724 429844 316736
rect 376720 316696 429844 316724
rect 376720 316684 376726 316696
rect 429838 316684 429844 316696
rect 429896 316684 429902 316736
rect 212258 316616 212264 316668
rect 212316 316656 212322 316668
rect 296990 316656 296996 316668
rect 212316 316628 296996 316656
rect 212316 316616 212322 316628
rect 296990 316616 296996 316628
rect 297048 316616 297054 316668
rect 314746 316616 314752 316668
rect 314804 316656 314810 316668
rect 315390 316656 315396 316668
rect 314804 316628 315396 316656
rect 314804 316616 314810 316628
rect 315390 316616 315396 316628
rect 315448 316616 315454 316668
rect 322658 316616 322664 316668
rect 322716 316656 322722 316668
rect 393498 316656 393504 316668
rect 322716 316628 393504 316656
rect 322716 316616 322722 316628
rect 393498 316616 393504 316628
rect 393556 316616 393562 316668
rect 308398 316548 308404 316600
rect 308456 316588 308462 316600
rect 329282 316588 329288 316600
rect 308456 316560 329288 316588
rect 308456 316548 308462 316560
rect 329282 316548 329288 316560
rect 329340 316548 329346 316600
rect 329374 316548 329380 316600
rect 329432 316588 329438 316600
rect 336550 316588 336556 316600
rect 329432 316560 336556 316588
rect 329432 316548 329438 316560
rect 336550 316548 336556 316560
rect 336608 316548 336614 316600
rect 303338 316480 303344 316532
rect 303396 316520 303402 316532
rect 329098 316520 329104 316532
rect 303396 316492 329104 316520
rect 303396 316480 303402 316492
rect 329098 316480 329104 316492
rect 329156 316480 329162 316532
rect 284662 316412 284668 316464
rect 284720 316452 284726 316464
rect 285306 316452 285312 316464
rect 284720 316424 285312 316452
rect 284720 316412 284726 316424
rect 285306 316412 285312 316424
rect 285364 316412 285370 316464
rect 324590 316412 324596 316464
rect 324648 316452 324654 316464
rect 392302 316452 392308 316464
rect 324648 316424 392308 316452
rect 324648 316412 324654 316424
rect 392302 316412 392308 316424
rect 392360 316412 392366 316464
rect 294322 316344 294328 316396
rect 294380 316384 294386 316396
rect 294874 316384 294880 316396
rect 294380 316356 294880 316384
rect 294380 316344 294386 316356
rect 294874 316344 294880 316356
rect 294932 316344 294938 316396
rect 295610 316344 295616 316396
rect 295668 316384 295674 316396
rect 295794 316384 295800 316396
rect 295668 316356 295800 316384
rect 295668 316344 295674 316356
rect 295794 316344 295800 316356
rect 295852 316344 295858 316396
rect 315390 316344 315396 316396
rect 315448 316384 315454 316396
rect 315942 316384 315948 316396
rect 315448 316356 315948 316384
rect 315448 316344 315454 316356
rect 315942 316344 315948 316356
rect 316000 316344 316006 316396
rect 329190 316344 329196 316396
rect 329248 316384 329254 316396
rect 336642 316384 336648 316396
rect 329248 316356 336648 316384
rect 329248 316344 329254 316356
rect 336642 316344 336648 316356
rect 336700 316344 336706 316396
rect 284662 316276 284668 316328
rect 284720 316316 284726 316328
rect 285122 316316 285128 316328
rect 284720 316288 285128 316316
rect 284720 316276 284726 316288
rect 285122 316276 285128 316288
rect 285180 316276 285186 316328
rect 287054 316276 287060 316328
rect 287112 316316 287118 316328
rect 287514 316316 287520 316328
rect 287112 316288 287520 316316
rect 287112 316276 287118 316288
rect 287514 316276 287520 316288
rect 287572 316276 287578 316328
rect 287790 316276 287796 316328
rect 287848 316316 287854 316328
rect 287974 316316 287980 316328
rect 287848 316288 287980 316316
rect 287848 316276 287854 316288
rect 287974 316276 287980 316288
rect 288032 316276 288038 316328
rect 292758 316276 292764 316328
rect 292816 316316 292822 316328
rect 299198 316316 299204 316328
rect 292816 316288 299204 316316
rect 292816 316276 292822 316288
rect 299198 316276 299204 316288
rect 299256 316276 299262 316328
rect 331674 316276 331680 316328
rect 331732 316316 331738 316328
rect 332042 316316 332048 316328
rect 331732 316288 332048 316316
rect 331732 316276 331738 316288
rect 332042 316276 332048 316288
rect 332100 316276 332106 316328
rect 282270 316208 282276 316260
rect 282328 316248 282334 316260
rect 300854 316248 300860 316260
rect 282328 316220 300860 316248
rect 282328 316208 282334 316220
rect 300854 316208 300860 316220
rect 300912 316208 300918 316260
rect 301682 316208 301688 316260
rect 301740 316248 301746 316260
rect 302142 316248 302148 316260
rect 301740 316220 302148 316248
rect 301740 316208 301746 316220
rect 302142 316208 302148 316220
rect 302200 316208 302206 316260
rect 302418 316208 302424 316260
rect 302476 316248 302482 316260
rect 303522 316248 303528 316260
rect 302476 316220 303528 316248
rect 302476 316208 302482 316220
rect 303522 316208 303528 316220
rect 303580 316208 303586 316260
rect 305270 316208 305276 316260
rect 305328 316248 305334 316260
rect 305546 316248 305552 316260
rect 305328 316220 305552 316248
rect 305328 316208 305334 316220
rect 305546 316208 305552 316220
rect 305604 316208 305610 316260
rect 312078 316208 312084 316260
rect 312136 316248 312142 316260
rect 312814 316248 312820 316260
rect 312136 316220 312820 316248
rect 312136 316208 312142 316220
rect 312814 316208 312820 316220
rect 312872 316208 312878 316260
rect 323026 316208 323032 316260
rect 323084 316248 323090 316260
rect 323486 316248 323492 316260
rect 323084 316220 323492 316248
rect 323084 316208 323090 316220
rect 323486 316208 323492 316220
rect 323544 316208 323550 316260
rect 276750 316140 276756 316192
rect 276808 316180 276814 316192
rect 303154 316180 303160 316192
rect 276808 316152 303160 316180
rect 276808 316140 276814 316152
rect 303154 316140 303160 316152
rect 303212 316180 303218 316192
rect 303338 316180 303344 316192
rect 303212 316152 303344 316180
rect 303212 316140 303218 316152
rect 303338 316140 303344 316152
rect 303396 316140 303402 316192
rect 307846 316140 307852 316192
rect 307904 316180 307910 316192
rect 308030 316180 308036 316192
rect 307904 316152 308036 316180
rect 307904 316140 307910 316152
rect 308030 316140 308036 316152
rect 308088 316140 308094 316192
rect 320910 316140 320916 316192
rect 320968 316180 320974 316192
rect 321278 316180 321284 316192
rect 320968 316152 321284 316180
rect 320968 316140 320974 316152
rect 321278 316140 321284 316152
rect 321336 316140 321342 316192
rect 322934 316140 322940 316192
rect 322992 316180 322998 316192
rect 324130 316180 324136 316192
rect 322992 316152 324136 316180
rect 322992 316140 322998 316152
rect 324130 316140 324136 316152
rect 324188 316140 324194 316192
rect 271322 316072 271328 316124
rect 271380 316112 271386 316124
rect 303706 316112 303712 316124
rect 271380 316084 303712 316112
rect 271380 316072 271386 316084
rect 303706 316072 303712 316084
rect 303764 316072 303770 316124
rect 303798 316072 303804 316124
rect 303856 316112 303862 316124
rect 304350 316112 304356 316124
rect 303856 316084 304356 316112
rect 303856 316072 303862 316084
rect 304350 316072 304356 316084
rect 304408 316072 304414 316124
rect 317690 316072 317696 316124
rect 317748 316112 317754 316124
rect 318334 316112 318340 316124
rect 317748 316084 318340 316112
rect 317748 316072 317754 316084
rect 318334 316072 318340 316084
rect 318392 316072 318398 316124
rect 323302 316072 323308 316124
rect 323360 316112 323366 316124
rect 324222 316112 324228 316124
rect 323360 316084 324228 316112
rect 323360 316072 323366 316084
rect 324222 316072 324228 316084
rect 324280 316072 324286 316124
rect 325050 316072 325056 316124
rect 325108 316112 325114 316124
rect 325418 316112 325424 316124
rect 325108 316084 325424 316112
rect 325108 316072 325114 316084
rect 325418 316072 325424 316084
rect 325476 316072 325482 316124
rect 325878 316072 325884 316124
rect 325936 316112 325942 316124
rect 326246 316112 326252 316124
rect 325936 316084 326252 316112
rect 325936 316072 325942 316084
rect 326246 316072 326252 316084
rect 326304 316072 326310 316124
rect 360194 316072 360200 316124
rect 360252 316112 360258 316124
rect 361390 316112 361396 316124
rect 360252 316084 361396 316112
rect 360252 316072 360258 316084
rect 361390 316072 361396 316084
rect 361448 316072 361454 316124
rect 217686 316004 217692 316056
rect 217744 316044 217750 316056
rect 292758 316044 292764 316056
rect 217744 316016 292764 316044
rect 217744 316004 217750 316016
rect 292758 316004 292764 316016
rect 292816 316004 292822 316056
rect 294322 316004 294328 316056
rect 294380 316044 294386 316056
rect 295150 316044 295156 316056
rect 294380 316016 295156 316044
rect 294380 316004 294386 316016
rect 295150 316004 295156 316016
rect 295208 316004 295214 316056
rect 297266 316004 297272 316056
rect 297324 316044 297330 316056
rect 297634 316044 297640 316056
rect 297324 316016 297640 316044
rect 297324 316004 297330 316016
rect 297634 316004 297640 316016
rect 297692 316004 297698 316056
rect 299842 316004 299848 316056
rect 299900 316044 299906 316056
rect 300578 316044 300584 316056
rect 299900 316016 300584 316044
rect 299900 316004 299906 316016
rect 300578 316004 300584 316016
rect 300636 316004 300642 316056
rect 301038 316004 301044 316056
rect 301096 316044 301102 316056
rect 302050 316044 302056 316056
rect 301096 316016 302056 316044
rect 301096 316004 301102 316016
rect 302050 316004 302056 316016
rect 302108 316004 302114 316056
rect 302234 316004 302240 316056
rect 302292 316044 302298 316056
rect 302970 316044 302976 316056
rect 302292 316016 302976 316044
rect 302292 316004 302298 316016
rect 302970 316004 302976 316016
rect 303028 316004 303034 316056
rect 305454 316004 305460 316056
rect 305512 316044 305518 316056
rect 305914 316044 305920 316056
rect 305512 316016 305920 316044
rect 305512 316004 305518 316016
rect 305914 316004 305920 316016
rect 305972 316004 305978 316056
rect 306742 316004 306748 316056
rect 306800 316044 306806 316056
rect 307294 316044 307300 316056
rect 306800 316016 307300 316044
rect 306800 316004 306806 316016
rect 307294 316004 307300 316016
rect 307352 316004 307358 316056
rect 308030 316004 308036 316056
rect 308088 316044 308094 316056
rect 308490 316044 308496 316056
rect 308088 316016 308496 316044
rect 308088 316004 308094 316016
rect 308490 316004 308496 316016
rect 308548 316004 308554 316056
rect 308582 316004 308588 316056
rect 308640 316044 308646 316056
rect 308950 316044 308956 316056
rect 308640 316016 308956 316044
rect 308640 316004 308646 316016
rect 308950 316004 308956 316016
rect 309008 316004 309014 316056
rect 310882 316004 310888 316056
rect 310940 316044 310946 316056
rect 311710 316044 311716 316056
rect 310940 316016 311716 316044
rect 310940 316004 310946 316016
rect 311710 316004 311716 316016
rect 311768 316004 311774 316056
rect 315022 316004 315028 316056
rect 315080 316044 315086 316056
rect 315482 316044 315488 316056
rect 315080 316016 315488 316044
rect 315080 316004 315086 316016
rect 315482 316004 315488 316016
rect 315540 316004 315546 316056
rect 316126 316004 316132 316056
rect 316184 316044 316190 316056
rect 316494 316044 316500 316056
rect 316184 316016 316500 316044
rect 316184 316004 316190 316016
rect 316494 316004 316500 316016
rect 316552 316004 316558 316056
rect 317506 316004 317512 316056
rect 317564 316044 317570 316056
rect 318242 316044 318248 316056
rect 317564 316016 318248 316044
rect 317564 316004 317570 316016
rect 318242 316004 318248 316016
rect 318300 316004 318306 316056
rect 320450 316004 320456 316056
rect 320508 316044 320514 316056
rect 321278 316044 321284 316056
rect 320508 316016 321284 316044
rect 320508 316004 320514 316016
rect 321278 316004 321284 316016
rect 321336 316004 321342 316056
rect 321554 316004 321560 316056
rect 321612 316044 321618 316056
rect 322842 316044 322848 316056
rect 321612 316016 322848 316044
rect 321612 316004 321618 316016
rect 322842 316004 322848 316016
rect 322900 316004 322906 316056
rect 323026 316004 323032 316056
rect 323084 316044 323090 316056
rect 323670 316044 323676 316056
rect 323084 316016 323676 316044
rect 323084 316004 323090 316016
rect 323670 316004 323676 316016
rect 323728 316004 323734 316056
rect 324406 316004 324412 316056
rect 324464 316044 324470 316056
rect 325602 316044 325608 316056
rect 324464 316016 325608 316044
rect 324464 316004 324470 316016
rect 325602 316004 325608 316016
rect 325660 316004 325666 316056
rect 325970 316004 325976 316056
rect 326028 316044 326034 316056
rect 326430 316044 326436 316056
rect 326028 316016 326436 316044
rect 326028 316004 326034 316016
rect 326430 316004 326436 316016
rect 326488 316004 326494 316056
rect 274358 315936 274364 315988
rect 274416 315976 274422 315988
rect 274416 315948 303338 315976
rect 274416 315936 274422 315948
rect 278774 315868 278780 315920
rect 278832 315908 278838 315920
rect 279142 315908 279148 315920
rect 278832 315880 279148 315908
rect 278832 315868 278838 315880
rect 279142 315868 279148 315880
rect 279200 315908 279206 315920
rect 279200 315880 302234 315908
rect 279200 315868 279206 315880
rect 270402 315800 270408 315852
rect 270460 315840 270466 315852
rect 270460 315812 292574 315840
rect 270460 315800 270466 315812
rect 268654 315772 268660 315784
rect 258046 315744 268660 315772
rect 214834 315460 214840 315512
rect 214892 315500 214898 315512
rect 258046 315500 258074 315744
rect 268654 315732 268660 315744
rect 268712 315772 268718 315784
rect 285766 315772 285772 315784
rect 268712 315744 285772 315772
rect 268712 315732 268718 315744
rect 285766 315732 285772 315744
rect 285824 315732 285830 315784
rect 286134 315732 286140 315784
rect 286192 315772 286198 315784
rect 286686 315772 286692 315784
rect 286192 315744 286692 315772
rect 286192 315732 286198 315744
rect 286686 315732 286692 315744
rect 286744 315732 286750 315784
rect 287330 315732 287336 315784
rect 287388 315772 287394 315784
rect 287698 315772 287704 315784
rect 287388 315744 287704 315772
rect 287388 315732 287394 315744
rect 287698 315732 287704 315744
rect 287756 315732 287762 315784
rect 287790 315732 287796 315784
rect 287848 315772 287854 315784
rect 288342 315772 288348 315784
rect 287848 315744 288348 315772
rect 287848 315732 287854 315744
rect 288342 315732 288348 315744
rect 288400 315732 288406 315784
rect 289262 315732 289268 315784
rect 289320 315772 289326 315784
rect 289722 315772 289728 315784
rect 289320 315744 289728 315772
rect 289320 315732 289326 315744
rect 289722 315732 289728 315744
rect 289780 315732 289786 315784
rect 290274 315732 290280 315784
rect 290332 315772 290338 315784
rect 290642 315772 290648 315784
rect 290332 315744 290648 315772
rect 290332 315732 290338 315744
rect 290642 315732 290648 315744
rect 290700 315732 290706 315784
rect 291286 315732 291292 315784
rect 291344 315772 291350 315784
rect 291562 315772 291568 315784
rect 291344 315744 291568 315772
rect 291344 315732 291350 315744
rect 291562 315732 291568 315744
rect 291620 315732 291626 315784
rect 292546 315772 292574 315812
rect 294230 315800 294236 315852
rect 294288 315840 294294 315852
rect 295242 315840 295248 315852
rect 294288 315812 295248 315840
rect 294288 315800 294294 315812
rect 295242 315800 295248 315812
rect 295300 315800 295306 315852
rect 295702 315800 295708 315852
rect 295760 315840 295766 315852
rect 296530 315840 296536 315852
rect 295760 315812 296536 315840
rect 295760 315800 295766 315812
rect 296530 315800 296536 315812
rect 296588 315800 296594 315852
rect 297358 315800 297364 315852
rect 297416 315840 297422 315852
rect 297910 315840 297916 315852
rect 297416 315812 297916 315840
rect 297416 315800 297422 315812
rect 297910 315800 297916 315812
rect 297968 315800 297974 315852
rect 298186 315800 298192 315852
rect 298244 315840 298250 315852
rect 299106 315840 299112 315852
rect 298244 315812 299112 315840
rect 298244 315800 298250 315812
rect 299106 315800 299112 315812
rect 299164 315800 299170 315852
rect 300026 315800 300032 315852
rect 300084 315840 300090 315852
rect 300394 315840 300400 315852
rect 300084 315812 300400 315840
rect 300084 315800 300090 315812
rect 300394 315800 300400 315812
rect 300452 315800 300458 315852
rect 301130 315800 301136 315852
rect 301188 315840 301194 315852
rect 301774 315840 301780 315852
rect 301188 315812 301780 315840
rect 301188 315800 301194 315812
rect 301774 315800 301780 315812
rect 301832 315800 301838 315852
rect 294414 315772 294420 315784
rect 292546 315744 294420 315772
rect 294414 315732 294420 315744
rect 294472 315732 294478 315784
rect 298278 315732 298284 315784
rect 298336 315772 298342 315784
rect 299382 315772 299388 315784
rect 298336 315744 299388 315772
rect 298336 315732 298342 315744
rect 299382 315732 299388 315744
rect 299440 315732 299446 315784
rect 299934 315732 299940 315784
rect 299992 315772 299998 315784
rect 300210 315772 300216 315784
rect 299992 315744 300216 315772
rect 299992 315732 299998 315744
rect 300210 315732 300216 315744
rect 300268 315732 300274 315784
rect 268746 315664 268752 315716
rect 268804 315704 268810 315716
rect 268804 315676 285996 315704
rect 268804 315664 268810 315676
rect 263318 315596 263324 315648
rect 263376 315636 263382 315648
rect 284846 315636 284852 315648
rect 263376 315608 284852 315636
rect 263376 315596 263382 315608
rect 284846 315596 284852 315608
rect 284904 315596 284910 315648
rect 285968 315568 285996 315676
rect 286042 315664 286048 315716
rect 286100 315704 286106 315716
rect 286778 315704 286784 315716
rect 286100 315676 286784 315704
rect 286100 315664 286106 315676
rect 286778 315664 286784 315676
rect 286836 315664 286842 315716
rect 287238 315664 287244 315716
rect 287296 315704 287302 315716
rect 287882 315704 287888 315716
rect 287296 315676 287888 315704
rect 287296 315664 287302 315676
rect 287882 315664 287888 315676
rect 287940 315664 287946 315716
rect 291470 315664 291476 315716
rect 291528 315704 291534 315716
rect 292390 315704 292396 315716
rect 291528 315676 292396 315704
rect 291528 315664 291534 315676
rect 292390 315664 292396 315676
rect 292448 315664 292454 315716
rect 296806 315664 296812 315716
rect 296864 315704 296870 315716
rect 297910 315704 297916 315716
rect 296864 315676 297916 315704
rect 296864 315664 296870 315676
rect 297910 315664 297916 315676
rect 297968 315664 297974 315716
rect 287422 315596 287428 315648
rect 287480 315636 287486 315648
rect 288066 315636 288072 315648
rect 287480 315608 288072 315636
rect 287480 315596 287486 315608
rect 288066 315596 288072 315608
rect 288124 315596 288130 315648
rect 291562 315596 291568 315648
rect 291620 315636 291626 315648
rect 292206 315636 292212 315648
rect 291620 315608 292212 315636
rect 291620 315596 291626 315608
rect 292206 315596 292212 315608
rect 292264 315596 292270 315648
rect 293218 315596 293224 315648
rect 293276 315636 293282 315648
rect 293770 315636 293776 315648
rect 293276 315608 293776 315636
rect 293276 315596 293282 315608
rect 293770 315596 293776 315608
rect 293828 315596 293834 315648
rect 291194 315568 291200 315580
rect 285968 315540 291200 315568
rect 291194 315528 291200 315540
rect 291252 315528 291258 315580
rect 302206 315568 302234 315880
rect 303310 315772 303338 315948
rect 306834 315936 306840 315988
rect 306892 315976 306898 315988
rect 307018 315976 307024 315988
rect 306892 315948 307024 315976
rect 306892 315936 306898 315948
rect 307018 315936 307024 315948
rect 307076 315936 307082 315988
rect 308214 315936 308220 315988
rect 308272 315976 308278 315988
rect 309042 315976 309048 315988
rect 308272 315948 309048 315976
rect 308272 315936 308278 315948
rect 309042 315936 309048 315948
rect 309100 315936 309106 315988
rect 309778 315936 309784 315988
rect 309836 315976 309842 315988
rect 310238 315976 310244 315988
rect 309836 315948 310244 315976
rect 309836 315936 309842 315948
rect 310238 315936 310244 315948
rect 310296 315936 310302 315988
rect 310698 315936 310704 315988
rect 310756 315976 310762 315988
rect 311434 315976 311440 315988
rect 310756 315948 311440 315976
rect 310756 315936 310762 315948
rect 311434 315936 311440 315948
rect 311492 315936 311498 315988
rect 311526 315936 311532 315988
rect 311584 315976 311590 315988
rect 311802 315976 311808 315988
rect 311584 315948 311808 315976
rect 311584 315936 311590 315948
rect 311802 315936 311808 315948
rect 311860 315936 311866 315988
rect 312170 315936 312176 315988
rect 312228 315976 312234 315988
rect 312630 315976 312636 315988
rect 312228 315948 312636 315976
rect 312228 315936 312234 315948
rect 312630 315936 312636 315948
rect 312688 315936 312694 315988
rect 314930 315936 314936 315988
rect 314988 315976 314994 315988
rect 315666 315976 315672 315988
rect 314988 315948 315672 315976
rect 314988 315936 314994 315948
rect 315666 315936 315672 315948
rect 315724 315936 315730 315988
rect 316218 315936 316224 315988
rect 316276 315976 316282 315988
rect 316954 315976 316960 315988
rect 316276 315948 316960 315976
rect 316276 315936 316282 315948
rect 316954 315936 316960 315948
rect 317012 315936 317018 315988
rect 317874 315936 317880 315988
rect 317932 315976 317938 315988
rect 318518 315976 318524 315988
rect 317932 315948 318524 315976
rect 317932 315936 317938 315948
rect 318518 315936 318524 315948
rect 318576 315936 318582 315988
rect 318628 315948 319208 315976
rect 304166 315868 304172 315920
rect 304224 315908 304230 315920
rect 304718 315908 304724 315920
rect 304224 315880 304724 315908
rect 304224 315868 304230 315880
rect 304718 315868 304724 315880
rect 304776 315868 304782 315920
rect 306650 315868 306656 315920
rect 306708 315908 306714 315920
rect 307662 315908 307668 315920
rect 306708 315880 307668 315908
rect 306708 315868 306714 315880
rect 307662 315868 307668 315880
rect 307720 315868 307726 315920
rect 308122 315868 308128 315920
rect 308180 315908 308186 315920
rect 308674 315908 308680 315920
rect 308180 315880 308680 315908
rect 308180 315868 308186 315880
rect 308674 315868 308680 315880
rect 308732 315868 308738 315920
rect 315206 315868 315212 315920
rect 315264 315908 315270 315920
rect 315942 315908 315948 315920
rect 315264 315880 315948 315908
rect 315264 315868 315270 315880
rect 315942 315868 315948 315880
rect 316000 315908 316006 315920
rect 318628 315908 318656 315948
rect 316000 315880 318656 315908
rect 316000 315868 316006 315880
rect 305178 315800 305184 315852
rect 305236 315840 305242 315852
rect 305730 315840 305736 315852
rect 305236 315812 305736 315840
rect 305236 315800 305242 315812
rect 305730 315800 305736 315812
rect 305788 315800 305794 315852
rect 307018 315800 307024 315852
rect 307076 315840 307082 315852
rect 307570 315840 307576 315852
rect 307076 315812 307576 315840
rect 307076 315800 307082 315812
rect 307570 315800 307576 315812
rect 307628 315800 307634 315852
rect 309686 315800 309692 315852
rect 309744 315840 309750 315852
rect 310238 315840 310244 315852
rect 309744 315812 310244 315840
rect 309744 315800 309750 315812
rect 310238 315800 310244 315812
rect 310296 315800 310302 315852
rect 314930 315800 314936 315852
rect 314988 315840 314994 315852
rect 315850 315840 315856 315852
rect 314988 315812 315856 315840
rect 314988 315800 314994 315812
rect 315850 315800 315856 315812
rect 315908 315800 315914 315852
rect 306466 315772 306472 315784
rect 303310 315744 306472 315772
rect 306466 315732 306472 315744
rect 306524 315772 306530 315784
rect 307754 315772 307760 315784
rect 306524 315744 307760 315772
rect 306524 315732 306530 315744
rect 307754 315732 307760 315744
rect 307812 315732 307818 315784
rect 313090 315732 313096 315784
rect 313148 315772 313154 315784
rect 313148 315744 317552 315772
rect 313148 315732 313154 315744
rect 313918 315664 313924 315716
rect 313976 315704 313982 315716
rect 314378 315704 314384 315716
rect 313976 315676 314384 315704
rect 313976 315664 313982 315676
rect 314378 315664 314384 315676
rect 314436 315664 314442 315716
rect 317524 315704 317552 315744
rect 317598 315732 317604 315784
rect 317656 315772 317662 315784
rect 318610 315772 318616 315784
rect 317656 315744 318616 315772
rect 317656 315732 317662 315744
rect 318610 315732 318616 315744
rect 318668 315732 318674 315784
rect 319180 315772 319208 315948
rect 320174 315936 320180 315988
rect 320232 315976 320238 315988
rect 320726 315976 320732 315988
rect 320232 315948 320732 315976
rect 320232 315936 320238 315948
rect 320726 315936 320732 315948
rect 320784 315976 320790 315988
rect 341426 315976 341432 315988
rect 320784 315948 341432 315976
rect 320784 315936 320790 315948
rect 341426 315936 341432 315948
rect 341484 315936 341490 315988
rect 361390 315936 361396 315988
rect 361448 315976 361454 315988
rect 366542 315976 366548 315988
rect 361448 315948 366548 315976
rect 361448 315936 361454 315948
rect 366542 315936 366548 315948
rect 366600 315936 366606 315988
rect 320450 315868 320456 315920
rect 320508 315908 320514 315920
rect 372890 315908 372896 315920
rect 320508 315880 372896 315908
rect 320508 315868 320514 315880
rect 372890 315868 372896 315880
rect 372948 315868 372954 315920
rect 319254 315800 319260 315852
rect 319312 315840 319318 315852
rect 372798 315840 372804 315852
rect 319312 315812 372804 315840
rect 319312 315800 319318 315812
rect 372798 315800 372804 315812
rect 372856 315800 372862 315852
rect 374178 315772 374184 315784
rect 319180 315744 374184 315772
rect 374178 315732 374184 315744
rect 374236 315732 374242 315784
rect 320450 315704 320456 315716
rect 317524 315676 320456 315704
rect 320450 315664 320456 315676
rect 320508 315664 320514 315716
rect 320542 315664 320548 315716
rect 320600 315704 320606 315716
rect 321094 315704 321100 315716
rect 320600 315676 321100 315704
rect 320600 315664 320606 315676
rect 321094 315664 321100 315676
rect 321152 315664 321158 315716
rect 321738 315664 321744 315716
rect 321796 315704 321802 315716
rect 322566 315704 322572 315716
rect 321796 315676 322572 315704
rect 321796 315664 321802 315676
rect 322566 315664 322572 315676
rect 322624 315664 322630 315716
rect 324038 315664 324044 315716
rect 324096 315704 324102 315716
rect 344922 315704 344928 315716
rect 324096 315676 344928 315704
rect 324096 315664 324102 315676
rect 344922 315664 344928 315676
rect 344980 315664 344986 315716
rect 303338 315596 303344 315648
rect 303396 315636 303402 315648
rect 328638 315636 328644 315648
rect 303396 315608 328644 315636
rect 303396 315596 303402 315608
rect 328638 315596 328644 315608
rect 328696 315596 328702 315648
rect 310974 315568 310980 315580
rect 302206 315540 310980 315568
rect 310974 315528 310980 315540
rect 311032 315528 311038 315580
rect 316770 315528 316776 315580
rect 316828 315568 316834 315580
rect 338298 315568 338304 315580
rect 316828 315540 338304 315568
rect 316828 315528 316834 315540
rect 338298 315528 338304 315540
rect 338356 315568 338362 315580
rect 354122 315568 354128 315580
rect 338356 315540 354128 315568
rect 338356 315528 338362 315540
rect 354122 315528 354128 315540
rect 354180 315528 354186 315580
rect 214892 315472 258074 315500
rect 214892 315460 214898 315472
rect 276658 315460 276664 315512
rect 276716 315500 276722 315512
rect 293678 315500 293684 315512
rect 276716 315472 293684 315500
rect 276716 315460 276722 315472
rect 293678 315460 293684 315472
rect 293736 315460 293742 315512
rect 293770 315460 293776 315512
rect 293828 315500 293834 315512
rect 306374 315500 306380 315512
rect 293828 315472 306380 315500
rect 293828 315460 293834 315472
rect 306374 315460 306380 315472
rect 306432 315460 306438 315512
rect 314654 315460 314660 315512
rect 314712 315500 314718 315512
rect 348878 315500 348884 315512
rect 314712 315472 348884 315500
rect 314712 315460 314718 315472
rect 348878 315460 348884 315472
rect 348936 315500 348942 315512
rect 374270 315500 374276 315512
rect 348936 315472 374276 315500
rect 348936 315460 348942 315472
rect 374270 315460 374276 315472
rect 374328 315460 374334 315512
rect 214926 315392 214932 315444
rect 214984 315432 214990 315444
rect 270402 315432 270408 315444
rect 214984 315404 270408 315432
rect 214984 315392 214990 315404
rect 270402 315392 270408 315404
rect 270460 315392 270466 315444
rect 273990 315392 273996 315444
rect 274048 315432 274054 315444
rect 294138 315432 294144 315444
rect 274048 315404 294144 315432
rect 274048 315392 274054 315404
rect 294138 315392 294144 315404
rect 294196 315392 294202 315444
rect 295150 315392 295156 315444
rect 295208 315432 295214 315444
rect 309594 315432 309600 315444
rect 295208 315404 309600 315432
rect 295208 315392 295214 315404
rect 309594 315392 309600 315404
rect 309652 315392 309658 315444
rect 316402 315392 316408 315444
rect 316460 315432 316466 315444
rect 351454 315432 351460 315444
rect 316460 315404 351460 315432
rect 316460 315392 316466 315404
rect 351454 315392 351460 315404
rect 351512 315432 351518 315444
rect 383470 315432 383476 315444
rect 351512 315404 383476 315432
rect 351512 315392 351518 315404
rect 383470 315392 383476 315404
rect 383528 315392 383534 315444
rect 209682 315324 209688 315376
rect 209740 315364 209746 315376
rect 268746 315364 268752 315376
rect 209740 315336 268752 315364
rect 209740 315324 209746 315336
rect 268746 315324 268752 315336
rect 268804 315324 268810 315376
rect 285766 315324 285772 315376
rect 285824 315364 285830 315376
rect 292022 315364 292028 315376
rect 285824 315336 292028 315364
rect 285824 315324 285830 315336
rect 292022 315324 292028 315336
rect 292080 315324 292086 315376
rect 293126 315324 293132 315376
rect 293184 315364 293190 315376
rect 293954 315364 293960 315376
rect 293184 315336 293960 315364
rect 293184 315324 293190 315336
rect 293954 315324 293960 315336
rect 294012 315324 294018 315376
rect 312446 315324 312452 315376
rect 312504 315364 312510 315376
rect 347590 315364 347596 315376
rect 312504 315336 347596 315364
rect 312504 315324 312510 315336
rect 347590 315324 347596 315336
rect 347648 315364 347654 315376
rect 384574 315364 384580 315376
rect 347648 315336 384580 315364
rect 347648 315324 347654 315336
rect 384574 315324 384580 315336
rect 384632 315324 384638 315376
rect 216398 315256 216404 315308
rect 216456 315296 216462 315308
rect 278774 315296 278780 315308
rect 216456 315268 278780 315296
rect 216456 315256 216462 315268
rect 278774 315256 278780 315268
rect 278832 315256 278838 315308
rect 292758 315256 292764 315308
rect 292816 315296 292822 315308
rect 293310 315296 293316 315308
rect 292816 315268 293316 315296
rect 292816 315256 292822 315268
rect 293310 315256 293316 315268
rect 293368 315256 293374 315308
rect 313734 315256 313740 315308
rect 313792 315296 313798 315308
rect 328638 315296 328644 315308
rect 313792 315268 328644 315296
rect 313792 315256 313798 315268
rect 328638 315256 328644 315268
rect 328696 315296 328702 315308
rect 382826 315296 382832 315308
rect 328696 315268 382832 315296
rect 328696 315256 328702 315268
rect 382826 315256 382832 315268
rect 382884 315296 382890 315308
rect 398926 315296 398932 315308
rect 382884 315268 398932 315296
rect 382884 315256 382890 315268
rect 398926 315256 398932 315268
rect 398984 315256 398990 315308
rect 278498 315188 278504 315240
rect 278556 315228 278562 315240
rect 320082 315228 320088 315240
rect 278556 315200 320088 315228
rect 278556 315188 278562 315200
rect 320082 315188 320088 315200
rect 320140 315188 320146 315240
rect 325510 315188 325516 315240
rect 325568 315228 325574 315240
rect 333882 315228 333888 315240
rect 325568 315200 333888 315228
rect 325568 315188 325574 315200
rect 333882 315188 333888 315200
rect 333940 315188 333946 315240
rect 312446 315120 312452 315172
rect 312504 315160 312510 315172
rect 312998 315160 313004 315172
rect 312504 315132 313004 315160
rect 312504 315120 312510 315132
rect 312998 315120 313004 315132
rect 313056 315120 313062 315172
rect 313918 315120 313924 315172
rect 313976 315160 313982 315172
rect 379974 315160 379980 315172
rect 313976 315132 379980 315160
rect 313976 315120 313982 315132
rect 379974 315120 379980 315132
rect 380032 315120 380038 315172
rect 280890 315052 280896 315104
rect 280948 315092 280954 315104
rect 319806 315092 319812 315104
rect 280948 315064 319812 315092
rect 280948 315052 280954 315064
rect 319806 315052 319812 315064
rect 319864 315052 319870 315104
rect 324866 315052 324872 315104
rect 324924 315092 324930 315104
rect 325602 315092 325608 315104
rect 324924 315064 325608 315092
rect 324924 315052 324930 315064
rect 325602 315052 325608 315064
rect 325660 315052 325666 315104
rect 300854 314984 300860 315036
rect 300912 315024 300918 315036
rect 328730 315024 328736 315036
rect 300912 314996 328736 315024
rect 300912 314984 300918 314996
rect 328730 314984 328736 314996
rect 328788 314984 328794 315036
rect 312998 314916 313004 314968
rect 313056 314956 313062 314968
rect 319254 314956 319260 314968
rect 313056 314928 319260 314956
rect 313056 314916 313062 314928
rect 319254 314916 319260 314928
rect 319312 314916 319318 314968
rect 324590 314916 324596 314968
rect 324648 314956 324654 314968
rect 325510 314956 325516 314968
rect 324648 314928 325516 314956
rect 324648 314916 324654 314928
rect 325510 314916 325516 314928
rect 325568 314916 325574 314968
rect 208302 314644 208308 314696
rect 208360 314684 208366 314696
rect 267366 314684 267372 314696
rect 208360 314656 267372 314684
rect 208360 314644 208366 314656
rect 267366 314644 267372 314656
rect 267424 314644 267430 314696
rect 271506 314576 271512 314628
rect 271564 314616 271570 314628
rect 271564 314588 273254 314616
rect 271564 314576 271570 314588
rect 273226 314548 273254 314588
rect 278406 314576 278412 314628
rect 278464 314616 278470 314628
rect 284754 314616 284760 314628
rect 278464 314588 284760 314616
rect 278464 314576 278470 314588
rect 284754 314576 284760 314588
rect 284812 314616 284818 314628
rect 285582 314616 285588 314628
rect 284812 314588 285588 314616
rect 284812 314576 284818 314588
rect 285582 314576 285588 314588
rect 285640 314576 285646 314628
rect 304902 314576 304908 314628
rect 304960 314616 304966 314628
rect 340598 314616 340604 314628
rect 304960 314588 340604 314616
rect 304960 314576 304966 314588
rect 340598 314576 340604 314588
rect 340656 314576 340662 314628
rect 284478 314548 284484 314560
rect 273226 314520 284484 314548
rect 284478 314508 284484 314520
rect 284536 314548 284542 314560
rect 285214 314548 285220 314560
rect 284536 314520 285220 314548
rect 284536 314508 284542 314520
rect 285214 314508 285220 314520
rect 285272 314508 285278 314560
rect 299198 314508 299204 314560
rect 299256 314548 299262 314560
rect 337746 314548 337752 314560
rect 299256 314520 337752 314548
rect 299256 314508 299262 314520
rect 337746 314508 337752 314520
rect 337804 314508 337810 314560
rect 277118 314440 277124 314492
rect 277176 314480 277182 314492
rect 280154 314480 280160 314492
rect 277176 314452 280160 314480
rect 277176 314440 277182 314452
rect 280154 314440 280160 314452
rect 280212 314440 280218 314492
rect 318150 314440 318156 314492
rect 318208 314480 318214 314492
rect 318610 314480 318616 314492
rect 318208 314452 318616 314480
rect 318208 314440 318214 314452
rect 318610 314440 318616 314452
rect 318668 314480 318674 314492
rect 384666 314480 384672 314492
rect 318668 314452 384672 314480
rect 318668 314440 318674 314452
rect 384666 314440 384672 314452
rect 384724 314440 384730 314492
rect 319070 314372 319076 314424
rect 319128 314412 319134 314424
rect 320082 314412 320088 314424
rect 319128 314384 320088 314412
rect 319128 314372 319134 314384
rect 320082 314372 320088 314384
rect 320140 314412 320146 314424
rect 380066 314412 380072 314424
rect 320140 314384 380072 314412
rect 320140 314372 320146 314384
rect 380066 314372 380072 314384
rect 380124 314372 380130 314424
rect 285950 314304 285956 314356
rect 286008 314344 286014 314356
rect 286502 314344 286508 314356
rect 286008 314316 286508 314344
rect 286008 314304 286014 314316
rect 286502 314304 286508 314316
rect 286560 314304 286566 314356
rect 316862 314304 316868 314356
rect 316920 314344 316926 314356
rect 376846 314344 376852 314356
rect 316920 314316 376852 314344
rect 316920 314304 316926 314316
rect 376846 314304 376852 314316
rect 376904 314304 376910 314356
rect 288710 314236 288716 314288
rect 288768 314276 288774 314288
rect 289078 314276 289084 314288
rect 288768 314248 289084 314276
rect 288768 314236 288774 314248
rect 289078 314236 289084 314248
rect 289136 314236 289142 314288
rect 318702 314236 318708 314288
rect 318760 314276 318766 314288
rect 378318 314276 378324 314288
rect 318760 314248 378324 314276
rect 318760 314236 318766 314248
rect 378318 314236 378324 314248
rect 378376 314236 378382 314288
rect 280154 314168 280160 314220
rect 280212 314208 280218 314220
rect 293494 314208 293500 314220
rect 280212 314180 293500 314208
rect 280212 314168 280218 314180
rect 293494 314168 293500 314180
rect 293552 314168 293558 314220
rect 296438 314168 296444 314220
rect 296496 314208 296502 314220
rect 356606 314208 356612 314220
rect 296496 314180 356612 314208
rect 296496 314168 296502 314180
rect 356606 314168 356612 314180
rect 356664 314168 356670 314220
rect 282178 314100 282184 314152
rect 282236 314140 282242 314152
rect 304074 314140 304080 314152
rect 282236 314112 304080 314140
rect 282236 314100 282242 314112
rect 304074 314100 304080 314112
rect 304132 314140 304138 314152
rect 363874 314140 363880 314152
rect 304132 314112 363880 314140
rect 304132 314100 304138 314112
rect 363874 314100 363880 314112
rect 363932 314100 363938 314152
rect 271414 314032 271420 314084
rect 271472 314072 271478 314084
rect 295978 314072 295984 314084
rect 271472 314044 295984 314072
rect 271472 314032 271478 314044
rect 295978 314032 295984 314044
rect 296036 314032 296042 314084
rect 311894 314032 311900 314084
rect 311952 314072 311958 314084
rect 312078 314072 312084 314084
rect 311952 314044 312084 314072
rect 311952 314032 311958 314044
rect 312078 314032 312084 314044
rect 312136 314032 312142 314084
rect 319162 314032 319168 314084
rect 319220 314072 319226 314084
rect 319990 314072 319996 314084
rect 319220 314044 319996 314072
rect 319220 314032 319226 314044
rect 319990 314032 319996 314044
rect 320048 314072 320054 314084
rect 379238 314072 379244 314084
rect 320048 314044 379244 314072
rect 320048 314032 320054 314044
rect 379238 314032 379244 314044
rect 379296 314032 379302 314084
rect 216214 313964 216220 314016
rect 216272 314004 216278 314016
rect 292574 314004 292580 314016
rect 216272 313976 292580 314004
rect 216272 313964 216278 313976
rect 292574 313964 292580 313976
rect 292632 313964 292638 314016
rect 300946 313964 300952 314016
rect 301004 314004 301010 314016
rect 301314 314004 301320 314016
rect 301004 313976 301320 314004
rect 301004 313964 301010 313976
rect 301314 313964 301320 313976
rect 301372 314004 301378 314016
rect 351362 314004 351368 314016
rect 301372 313976 351368 314004
rect 301372 313964 301378 313976
rect 351362 313964 351368 313976
rect 351420 313964 351426 314016
rect 220446 313896 220452 313948
rect 220504 313936 220510 313948
rect 314194 313936 314200 313948
rect 220504 313908 314200 313936
rect 220504 313896 220510 313908
rect 314194 313896 314200 313908
rect 314252 313896 314258 313948
rect 322382 313896 322388 313948
rect 322440 313936 322446 313948
rect 322750 313936 322756 313948
rect 322440 313908 322756 313936
rect 322440 313896 322446 313908
rect 322750 313896 322756 313908
rect 322808 313896 322814 313948
rect 324774 313896 324780 313948
rect 324832 313936 324838 313948
rect 330018 313936 330024 313948
rect 324832 313908 330024 313936
rect 324832 313896 324838 313908
rect 330018 313896 330024 313908
rect 330076 313936 330082 313948
rect 337654 313936 337660 313948
rect 330076 313908 337660 313936
rect 330076 313896 330082 313908
rect 337654 313896 337660 313908
rect 337712 313896 337718 313948
rect 378318 313896 378324 313948
rect 378376 313936 378382 313948
rect 466454 313936 466460 313948
rect 378376 313908 466460 313936
rect 378376 313896 378382 313908
rect 466454 313896 466460 313908
rect 466512 313896 466518 313948
rect 300946 313828 300952 313880
rect 301004 313868 301010 313880
rect 301590 313868 301596 313880
rect 301004 313840 301596 313868
rect 301004 313828 301010 313840
rect 301590 313828 301596 313840
rect 301648 313828 301654 313880
rect 310974 313828 310980 313880
rect 311032 313868 311038 313880
rect 329926 313868 329932 313880
rect 311032 313840 329932 313868
rect 311032 313828 311038 313840
rect 329926 313828 329932 313840
rect 329984 313828 329990 313880
rect 312078 313760 312084 313812
rect 312136 313800 312142 313812
rect 312722 313800 312728 313812
rect 312136 313772 312728 313800
rect 312136 313760 312142 313772
rect 312722 313760 312728 313772
rect 312780 313760 312786 313812
rect 318150 313760 318156 313812
rect 318208 313800 318214 313812
rect 318702 313800 318708 313812
rect 318208 313772 318708 313800
rect 318208 313760 318214 313772
rect 318702 313760 318708 313772
rect 318760 313760 318766 313812
rect 386046 313800 386052 313812
rect 321526 313772 386052 313800
rect 317322 313692 317328 313744
rect 317380 313732 317386 313744
rect 321526 313732 321554 313772
rect 386046 313760 386052 313772
rect 386104 313760 386110 313812
rect 317380 313704 321554 313732
rect 317380 313692 317386 313704
rect 322750 313692 322756 313744
rect 322808 313732 322814 313744
rect 389542 313732 389548 313744
rect 322808 313704 389548 313732
rect 322808 313692 322814 313704
rect 389542 313692 389548 313704
rect 389600 313692 389606 313744
rect 329926 313624 329932 313676
rect 329984 313664 329990 313676
rect 330110 313664 330116 313676
rect 329984 313636 330116 313664
rect 329984 313624 329990 313636
rect 330110 313624 330116 313636
rect 330168 313624 330174 313676
rect 293678 313488 293684 313540
rect 293736 313528 293742 313540
rect 300854 313528 300860 313540
rect 293736 313500 300860 313528
rect 293736 313488 293742 313500
rect 300854 313488 300860 313500
rect 300912 313488 300918 313540
rect 275830 313420 275836 313472
rect 275888 313460 275894 313472
rect 293862 313460 293868 313472
rect 275888 313432 293868 313460
rect 275888 313420 275894 313432
rect 293862 313420 293868 313432
rect 293920 313420 293926 313472
rect 327442 313420 327448 313472
rect 327500 313460 327506 313472
rect 328270 313460 328276 313472
rect 327500 313432 328276 313460
rect 327500 313420 327506 313432
rect 328270 313420 328276 313432
rect 328328 313420 328334 313472
rect 215202 313352 215208 313404
rect 215260 313392 215266 313404
rect 298094 313392 298100 313404
rect 215260 313364 298100 313392
rect 215260 313352 215266 313364
rect 298094 313352 298100 313364
rect 298152 313352 298158 313404
rect 212442 313284 212448 313336
rect 212500 313324 212506 313336
rect 293678 313324 293684 313336
rect 212500 313296 293684 313324
rect 212500 313284 212506 313296
rect 293678 313284 293684 313296
rect 293736 313284 293742 313336
rect 293862 313284 293868 313336
rect 293920 313324 293926 313336
rect 299842 313324 299848 313336
rect 293920 313296 299848 313324
rect 293920 313284 293926 313296
rect 299842 313284 299848 313296
rect 299900 313284 299906 313336
rect 311894 313284 311900 313336
rect 311952 313324 311958 313336
rect 319622 313324 319628 313336
rect 311952 313296 319628 313324
rect 311952 313284 311958 313296
rect 319622 313284 319628 313296
rect 319680 313284 319686 313336
rect 263226 313216 263232 313268
rect 263284 313256 263290 313268
rect 287054 313256 287060 313268
rect 263284 313228 287060 313256
rect 263284 313216 263290 313228
rect 287054 313216 287060 313228
rect 287112 313216 287118 313268
rect 308306 313216 308312 313268
rect 308364 313256 308370 313268
rect 309042 313256 309048 313268
rect 308364 313228 309048 313256
rect 308364 313216 308370 313228
rect 309042 313216 309048 313228
rect 309100 313216 309106 313268
rect 309870 313216 309876 313268
rect 309928 313256 309934 313268
rect 310054 313256 310060 313268
rect 309928 313228 310060 313256
rect 309928 313216 309934 313228
rect 310054 313216 310060 313228
rect 310112 313216 310118 313268
rect 327074 313256 327080 313268
rect 310164 313228 327080 313256
rect 277026 313148 277032 313200
rect 277084 313188 277090 313200
rect 278866 313188 278872 313200
rect 277084 313160 278872 313188
rect 277084 313148 277090 313160
rect 278866 313148 278872 313160
rect 278924 313148 278930 313200
rect 307754 313148 307760 313200
rect 307812 313188 307818 313200
rect 310164 313188 310192 313228
rect 327074 313216 327080 313228
rect 327132 313216 327138 313268
rect 327810 313216 327816 313268
rect 327868 313256 327874 313268
rect 330202 313256 330208 313268
rect 327868 313228 330208 313256
rect 327868 313216 327874 313228
rect 330202 313216 330208 313228
rect 330260 313216 330266 313268
rect 333514 313216 333520 313268
rect 333572 313256 333578 313268
rect 333882 313256 333888 313268
rect 333572 313228 333888 313256
rect 333572 313216 333578 313228
rect 333882 313216 333888 313228
rect 333940 313256 333946 313268
rect 340414 313256 340420 313268
rect 333940 313228 340420 313256
rect 333940 313216 333946 313228
rect 340414 313216 340420 313228
rect 340472 313216 340478 313268
rect 534718 313216 534724 313268
rect 534776 313256 534782 313268
rect 579614 313256 579620 313268
rect 534776 313228 579620 313256
rect 534776 313216 534782 313228
rect 579614 313216 579620 313228
rect 579672 313216 579678 313268
rect 329006 313188 329012 313200
rect 307812 313160 310192 313188
rect 310256 313160 329012 313188
rect 307812 313148 307818 313160
rect 309042 313080 309048 313132
rect 309100 313120 309106 313132
rect 310256 313120 310284 313160
rect 329006 313148 329012 313160
rect 329064 313148 329070 313200
rect 309100 313092 310284 313120
rect 309100 313080 309106 313092
rect 311618 313080 311624 313132
rect 311676 313120 311682 313132
rect 371602 313120 371608 313132
rect 311676 313092 371608 313120
rect 311676 313080 311682 313092
rect 371602 313080 371608 313092
rect 371660 313080 371666 313132
rect 317138 313012 317144 313064
rect 317196 313052 317202 313064
rect 377674 313052 377680 313064
rect 317196 313024 377680 313052
rect 317196 313012 317202 313024
rect 377674 313012 377680 313024
rect 377732 313012 377738 313064
rect 303706 312944 303712 312996
rect 303764 312984 303770 312996
rect 365162 312984 365168 312996
rect 303764 312956 365168 312984
rect 303764 312944 303770 312956
rect 365162 312944 365168 312956
rect 365220 312944 365226 312996
rect 310330 312876 310336 312928
rect 310388 312916 310394 312928
rect 370314 312916 370320 312928
rect 310388 312888 370320 312916
rect 310388 312876 310394 312888
rect 370314 312876 370320 312888
rect 370372 312876 370378 312928
rect 298094 312808 298100 312860
rect 298152 312848 298158 312860
rect 298646 312848 298652 312860
rect 298152 312820 298652 312848
rect 298152 312808 298158 312820
rect 298646 312808 298652 312820
rect 298704 312848 298710 312860
rect 358722 312848 358728 312860
rect 298704 312820 358728 312848
rect 298704 312808 298710 312820
rect 358722 312808 358728 312820
rect 358780 312808 358786 312860
rect 209498 312740 209504 312792
rect 209556 312780 209562 312792
rect 263226 312780 263232 312792
rect 209556 312752 263232 312780
rect 209556 312740 209562 312752
rect 263226 312740 263232 312752
rect 263284 312740 263290 312792
rect 294598 312780 294604 312792
rect 292546 312752 294604 312780
rect 210878 312672 210884 312724
rect 210936 312712 210942 312724
rect 265894 312712 265900 312724
rect 210936 312684 265900 312712
rect 210936 312672 210942 312684
rect 265894 312672 265900 312684
rect 265952 312672 265958 312724
rect 277946 312672 277952 312724
rect 278004 312712 278010 312724
rect 292546 312712 292574 312752
rect 294598 312740 294604 312752
rect 294656 312780 294662 312792
rect 342070 312780 342076 312792
rect 294656 312752 342076 312780
rect 294656 312740 294662 312752
rect 342070 312740 342076 312752
rect 342128 312740 342134 312792
rect 278004 312684 292574 312712
rect 278004 312672 278010 312684
rect 303614 312672 303620 312724
rect 303672 312712 303678 312724
rect 350166 312712 350172 312724
rect 303672 312684 350172 312712
rect 303672 312672 303678 312684
rect 350166 312672 350172 312684
rect 350224 312672 350230 312724
rect 205450 312604 205456 312656
rect 205508 312644 205514 312656
rect 288250 312644 288256 312656
rect 205508 312616 288256 312644
rect 205508 312604 205514 312616
rect 288250 312604 288256 312616
rect 288308 312604 288314 312656
rect 309870 312604 309876 312656
rect 309928 312644 309934 312656
rect 328822 312644 328828 312656
rect 309928 312616 328828 312644
rect 309928 312604 309934 312616
rect 328822 312604 328828 312616
rect 328880 312604 328886 312656
rect 334250 312604 334256 312656
rect 334308 312644 334314 312656
rect 390646 312644 390652 312656
rect 334308 312616 390652 312644
rect 334308 312604 334314 312616
rect 390646 312604 390652 312616
rect 390704 312604 390710 312656
rect 219158 312536 219164 312588
rect 219216 312576 219222 312588
rect 310974 312576 310980 312588
rect 219216 312548 310980 312576
rect 219216 312536 219222 312548
rect 310974 312536 310980 312548
rect 311032 312536 311038 312588
rect 320634 312536 320640 312588
rect 320692 312576 320698 312588
rect 321186 312576 321192 312588
rect 320692 312548 321192 312576
rect 320692 312536 320698 312548
rect 321186 312536 321192 312548
rect 321244 312536 321250 312588
rect 323946 312536 323952 312588
rect 324004 312576 324010 312588
rect 330110 312576 330116 312588
rect 324004 312548 330116 312576
rect 324004 312536 324010 312548
rect 330110 312536 330116 312548
rect 330168 312576 330174 312588
rect 389450 312576 389456 312588
rect 330168 312548 389456 312576
rect 330168 312536 330174 312548
rect 389450 312536 389456 312548
rect 389508 312536 389514 312588
rect 498194 312576 498200 312588
rect 393286 312548 498200 312576
rect 300118 312468 300124 312520
rect 300176 312508 300182 312520
rect 343542 312508 343548 312520
rect 300176 312480 343548 312508
rect 300176 312468 300182 312480
rect 343542 312468 343548 312480
rect 343600 312468 343606 312520
rect 319806 312400 319812 312452
rect 319864 312440 319870 312452
rect 320726 312440 320732 312452
rect 319864 312412 320732 312440
rect 319864 312400 319870 312412
rect 320726 312400 320732 312412
rect 320784 312400 320790 312452
rect 320818 312332 320824 312384
rect 320876 312372 320882 312384
rect 321370 312372 321376 312384
rect 320876 312344 321376 312372
rect 320876 312332 320882 312344
rect 321370 312332 321376 312344
rect 321428 312372 321434 312384
rect 392210 312372 392216 312384
rect 321428 312344 392216 312372
rect 321428 312332 321434 312344
rect 392210 312332 392216 312344
rect 392268 312372 392274 312384
rect 393286 312372 393314 312548
rect 498194 312536 498200 312548
rect 498252 312536 498258 312588
rect 392268 312344 393314 312372
rect 392268 312332 392274 312344
rect 322106 312264 322112 312316
rect 322164 312304 322170 312316
rect 388070 312304 388076 312316
rect 322164 312276 388076 312304
rect 322164 312264 322170 312276
rect 388070 312264 388076 312276
rect 388128 312264 388134 312316
rect 313182 312196 313188 312248
rect 313240 312236 313246 312248
rect 323118 312236 323124 312248
rect 313240 312208 323124 312236
rect 313240 312196 313246 312208
rect 323118 312196 323124 312208
rect 323176 312196 323182 312248
rect 278866 311992 278872 312044
rect 278924 312032 278930 312044
rect 309134 312032 309140 312044
rect 278924 312004 309140 312032
rect 278924 311992 278930 312004
rect 309134 311992 309140 312004
rect 309192 311992 309198 312044
rect 282730 311924 282736 311976
rect 282788 311964 282794 311976
rect 319806 311964 319812 311976
rect 282788 311936 319812 311964
rect 282788 311924 282794 311936
rect 319806 311924 319812 311936
rect 319864 311924 319870 311976
rect 278590 311856 278596 311908
rect 278648 311896 278654 311908
rect 320634 311896 320640 311908
rect 278648 311868 320640 311896
rect 278648 311856 278654 311868
rect 320634 311856 320640 311868
rect 320692 311856 320698 311908
rect 259270 311828 259276 311840
rect 258046 311800 259276 311828
rect 202598 311448 202604 311500
rect 202656 311488 202662 311500
rect 258046 311488 258074 311800
rect 259270 311788 259276 311800
rect 259328 311828 259334 311840
rect 288526 311828 288532 311840
rect 259328 311800 288532 311828
rect 259328 311788 259334 311800
rect 288526 311788 288532 311800
rect 288584 311788 288590 311840
rect 312446 311788 312452 311840
rect 312504 311828 312510 311840
rect 313182 311828 313188 311840
rect 312504 311800 313188 311828
rect 312504 311788 312510 311800
rect 313182 311788 313188 311800
rect 313240 311788 313246 311840
rect 313550 311788 313556 311840
rect 313608 311828 313614 311840
rect 314562 311828 314568 311840
rect 313608 311800 314568 311828
rect 313608 311788 313614 311800
rect 314562 311788 314568 311800
rect 314620 311828 314626 311840
rect 375282 311828 375288 311840
rect 314620 311800 375288 311828
rect 314620 311788 314626 311800
rect 375282 311788 375288 311800
rect 375340 311788 375346 311840
rect 263042 311720 263048 311772
rect 263100 311760 263106 311772
rect 263410 311760 263416 311772
rect 263100 311732 263416 311760
rect 263100 311720 263106 311732
rect 263410 311720 263416 311732
rect 263468 311760 263474 311772
rect 288618 311760 288624 311772
rect 263468 311732 288624 311760
rect 263468 311720 263474 311732
rect 288618 311720 288624 311732
rect 288676 311720 288682 311772
rect 310974 311720 310980 311772
rect 311032 311760 311038 311772
rect 311802 311760 311808 311772
rect 311032 311732 311808 311760
rect 311032 311720 311038 311732
rect 311802 311720 311808 311732
rect 311860 311760 311866 311772
rect 371418 311760 371424 311772
rect 311860 311732 371424 311760
rect 311860 311720 311866 311732
rect 371418 311720 371424 311732
rect 371476 311720 371482 311772
rect 297266 311652 297272 311704
rect 297324 311692 297330 311704
rect 356974 311692 356980 311704
rect 297324 311664 356980 311692
rect 297324 311652 297330 311664
rect 356974 311652 356980 311664
rect 357032 311652 357038 311704
rect 294690 311584 294696 311636
rect 294748 311624 294754 311636
rect 300210 311624 300216 311636
rect 294748 311596 300216 311624
rect 294748 311584 294754 311596
rect 300210 311584 300216 311596
rect 300268 311584 300274 311636
rect 313274 311584 313280 311636
rect 313332 311624 313338 311636
rect 313642 311624 313648 311636
rect 313332 311596 313648 311624
rect 313332 311584 313338 311596
rect 313642 311584 313648 311596
rect 313700 311624 313706 311636
rect 373350 311624 373356 311636
rect 313700 311596 373356 311624
rect 313700 311584 313706 311596
rect 373350 311584 373356 311596
rect 373408 311584 373414 311636
rect 298922 311516 298928 311568
rect 298980 311556 298986 311568
rect 358170 311556 358176 311568
rect 298980 311528 358176 311556
rect 298980 311516 298986 311528
rect 358170 311516 358176 311528
rect 358228 311516 358234 311568
rect 202656 311460 258074 311488
rect 202656 311448 202662 311460
rect 289262 311448 289268 311500
rect 289320 311488 289326 311500
rect 302878 311488 302884 311500
rect 289320 311460 302884 311488
rect 289320 311448 289326 311460
rect 302878 311448 302884 311460
rect 302936 311488 302942 311500
rect 361666 311488 361672 311500
rect 302936 311460 361672 311488
rect 302936 311448 302942 311460
rect 361666 311448 361672 311460
rect 361724 311448 361730 311500
rect 208118 311380 208124 311432
rect 208176 311420 208182 311432
rect 270126 311420 270132 311432
rect 208176 311392 270132 311420
rect 208176 311380 208182 311392
rect 270126 311380 270132 311392
rect 270184 311380 270190 311432
rect 297358 311380 297364 311432
rect 297416 311420 297422 311432
rect 355502 311420 355508 311432
rect 297416 311392 355508 311420
rect 297416 311380 297422 311392
rect 355502 311380 355508 311392
rect 355560 311380 355566 311432
rect 200022 311312 200028 311364
rect 200080 311352 200086 311364
rect 263042 311352 263048 311364
rect 200080 311324 263048 311352
rect 200080 311312 200086 311324
rect 263042 311312 263048 311324
rect 263100 311312 263106 311364
rect 267642 311312 267648 311364
rect 267700 311352 267706 311364
rect 271874 311352 271880 311364
rect 267700 311324 271880 311352
rect 267700 311312 267706 311324
rect 271874 311312 271880 311324
rect 271932 311352 271938 311364
rect 286318 311352 286324 311364
rect 271932 311324 286324 311352
rect 271932 311312 271938 311324
rect 286318 311312 286324 311324
rect 286376 311312 286382 311364
rect 286410 311312 286416 311364
rect 286468 311352 286474 311364
rect 309962 311352 309968 311364
rect 286468 311324 309968 311352
rect 286468 311312 286474 311324
rect 309962 311312 309968 311324
rect 310020 311352 310026 311364
rect 362218 311352 362224 311364
rect 310020 311324 362224 311352
rect 310020 311312 310026 311324
rect 362218 311312 362224 311324
rect 362276 311312 362282 311364
rect 214742 311244 214748 311296
rect 214800 311284 214806 311296
rect 281626 311284 281632 311296
rect 214800 311256 281632 311284
rect 214800 311244 214806 311256
rect 281626 311244 281632 311256
rect 281684 311244 281690 311296
rect 283742 311244 283748 311296
rect 283800 311284 283806 311296
rect 313274 311284 313280 311296
rect 283800 311256 313280 311284
rect 283800 311244 283806 311256
rect 313274 311244 313280 311256
rect 313332 311244 313338 311296
rect 323118 311244 323124 311296
rect 323176 311284 323182 311296
rect 371510 311284 371516 311296
rect 323176 311256 371516 311284
rect 323176 311244 323182 311256
rect 371510 311244 371516 311256
rect 371568 311244 371574 311296
rect 211982 311176 211988 311228
rect 212040 311216 212046 311228
rect 284846 311216 284852 311228
rect 212040 311188 284852 311216
rect 212040 311176 212046 311188
rect 284846 311176 284852 311188
rect 284904 311176 284910 311228
rect 295702 311176 295708 311228
rect 295760 311216 295766 311228
rect 295978 311216 295984 311228
rect 295760 311188 295984 311216
rect 295760 311176 295766 311188
rect 295978 311176 295984 311188
rect 296036 311216 296042 311228
rect 339126 311216 339132 311228
rect 296036 311188 339132 311216
rect 296036 311176 296042 311188
rect 339126 311176 339132 311188
rect 339184 311176 339190 311228
rect 204162 311108 204168 311160
rect 204220 311148 204226 311160
rect 284386 311148 284392 311160
rect 204220 311120 284392 311148
rect 204220 311108 204226 311120
rect 284386 311108 284392 311120
rect 284444 311108 284450 311160
rect 293218 311108 293224 311160
rect 293276 311148 293282 311160
rect 333330 311148 333336 311160
rect 293276 311120 333336 311148
rect 293276 311108 293282 311120
rect 333330 311108 333336 311120
rect 333388 311108 333394 311160
rect 342254 311148 342260 311160
rect 335326 311120 342260 311148
rect 308214 311040 308220 311092
rect 308272 311080 308278 311092
rect 335326 311080 335354 311120
rect 342254 311108 342260 311120
rect 342312 311148 342318 311160
rect 343450 311148 343456 311160
rect 342312 311120 343456 311148
rect 342312 311108 342318 311120
rect 343450 311108 343456 311120
rect 343508 311108 343514 311160
rect 308272 311052 335354 311080
rect 308272 311040 308278 311052
rect 296714 310972 296720 311024
rect 296772 311012 296778 311024
rect 297450 311012 297456 311024
rect 296772 310984 297456 311012
rect 296772 310972 296778 310984
rect 297450 310972 297456 310984
rect 297508 311012 297514 311024
rect 331950 311012 331956 311024
rect 297508 310984 331956 311012
rect 297508 310972 297514 310984
rect 331950 310972 331956 310984
rect 332008 310972 332014 311024
rect 310790 310904 310796 310956
rect 310848 310944 310854 310956
rect 311158 310944 311164 310956
rect 310848 310916 311164 310944
rect 310848 310904 310854 310916
rect 311158 310904 311164 310916
rect 311216 310944 311222 310956
rect 340322 310944 340328 310956
rect 311216 310916 340328 310944
rect 311216 310904 311222 310916
rect 340322 310904 340328 310916
rect 340380 310904 340386 310956
rect 212166 310428 212172 310480
rect 212224 310468 212230 310480
rect 212224 310440 277394 310468
rect 212224 310428 212230 310440
rect 277366 310332 277394 310440
rect 298554 310428 298560 310480
rect 298612 310468 298618 310480
rect 299106 310468 299112 310480
rect 298612 310440 299112 310468
rect 298612 310428 298618 310440
rect 299106 310428 299112 310440
rect 299164 310428 299170 310480
rect 313458 310428 313464 310480
rect 313516 310468 313522 310480
rect 314194 310468 314200 310480
rect 313516 310440 314200 310468
rect 313516 310428 313522 310440
rect 314194 310428 314200 310440
rect 314252 310468 314258 310480
rect 374914 310468 374920 310480
rect 314252 310440 374920 310468
rect 314252 310428 314258 310440
rect 374914 310428 374920 310440
rect 374972 310468 374978 310480
rect 375282 310468 375288 310480
rect 374972 310440 375288 310468
rect 374972 310428 374978 310440
rect 375282 310428 375288 310440
rect 375340 310428 375346 310480
rect 287882 310360 287888 310412
rect 287940 310400 287946 310412
rect 303614 310400 303620 310412
rect 287940 310372 303620 310400
rect 287940 310360 287946 310372
rect 303614 310360 303620 310372
rect 303672 310360 303678 310412
rect 312262 310360 312268 310412
rect 312320 310400 312326 310412
rect 312906 310400 312912 310412
rect 312320 310372 312912 310400
rect 312320 310360 312326 310372
rect 312906 310360 312912 310372
rect 312964 310400 312970 310412
rect 373626 310400 373632 310412
rect 312964 310372 373632 310400
rect 312964 310360 312970 310372
rect 373626 310360 373632 310372
rect 373684 310360 373690 310412
rect 296714 310332 296720 310344
rect 277366 310304 296720 310332
rect 296714 310292 296720 310304
rect 296772 310292 296778 310344
rect 355410 310332 355416 310344
rect 298940 310304 355416 310332
rect 282362 310224 282368 310276
rect 282420 310264 282426 310276
rect 298830 310264 298836 310276
rect 282420 310236 298836 310264
rect 282420 310224 282426 310236
rect 298830 310224 298836 310236
rect 298888 310224 298894 310276
rect 282822 310156 282828 310208
rect 282880 310196 282886 310208
rect 291838 310196 291844 310208
rect 282880 310168 291844 310196
rect 282880 310156 282886 310168
rect 291838 310156 291844 310168
rect 291896 310156 291902 310208
rect 296070 310196 296076 310208
rect 293236 310168 296076 310196
rect 287054 310128 287060 310140
rect 277366 310100 287060 310128
rect 265986 310020 265992 310072
rect 266044 310060 266050 310072
rect 273346 310060 273352 310072
rect 266044 310032 273352 310060
rect 266044 310020 266050 310032
rect 273346 310020 273352 310032
rect 273404 310060 273410 310072
rect 277366 310060 277394 310100
rect 287054 310088 287060 310100
rect 287112 310088 287118 310140
rect 273404 310032 277394 310060
rect 273404 310020 273410 310032
rect 279970 310020 279976 310072
rect 280028 310060 280034 310072
rect 293236 310060 293264 310168
rect 296070 310156 296076 310168
rect 296128 310196 296134 310208
rect 298940 310196 298968 310304
rect 355410 310292 355416 310304
rect 355468 310292 355474 310344
rect 317506 310224 317512 310276
rect 317564 310264 317570 310276
rect 318610 310264 318616 310276
rect 317564 310236 318616 310264
rect 317564 310224 317570 310236
rect 318610 310224 318616 310236
rect 318668 310264 318674 310276
rect 376294 310264 376300 310276
rect 318668 310236 376300 310264
rect 318668 310224 318674 310236
rect 376294 310224 376300 310236
rect 376352 310224 376358 310276
rect 296128 310168 298968 310196
rect 296128 310156 296134 310168
rect 299106 310156 299112 310208
rect 299164 310196 299170 310208
rect 356882 310196 356888 310208
rect 299164 310168 356888 310196
rect 299164 310156 299170 310168
rect 356882 310156 356888 310168
rect 356940 310156 356946 310208
rect 294322 310088 294328 310140
rect 294380 310128 294386 310140
rect 294966 310128 294972 310140
rect 294380 310100 294972 310128
rect 294380 310088 294386 310100
rect 294966 310088 294972 310100
rect 295024 310128 295030 310140
rect 344738 310128 344744 310140
rect 295024 310100 344744 310128
rect 295024 310088 295030 310100
rect 344738 310088 344744 310100
rect 344796 310088 344802 310140
rect 280028 310032 293264 310060
rect 280028 310020 280034 310032
rect 298830 310020 298836 310072
rect 298888 310060 298894 310072
rect 301314 310060 301320 310072
rect 298888 310032 301320 310060
rect 298888 310020 298894 310032
rect 301314 310020 301320 310032
rect 301372 310020 301378 310072
rect 347406 310060 347412 310072
rect 306346 310032 347412 310060
rect 222194 309952 222200 310004
rect 222252 309992 222258 310004
rect 282638 309992 282644 310004
rect 222252 309964 282644 309992
rect 222252 309952 222258 309964
rect 282638 309952 282644 309964
rect 282696 309952 282702 310004
rect 283650 309952 283656 310004
rect 283708 309992 283714 310004
rect 302142 309992 302148 310004
rect 283708 309964 302148 309992
rect 283708 309952 283714 309964
rect 302142 309952 302148 309964
rect 302200 309992 302206 310004
rect 306346 309992 306374 310032
rect 347406 310020 347412 310032
rect 347464 310020 347470 310072
rect 302200 309964 306374 309992
rect 302200 309952 302206 309964
rect 308122 309952 308128 310004
rect 308180 309992 308186 310004
rect 354030 309992 354036 310004
rect 308180 309964 354036 309992
rect 308180 309952 308186 309964
rect 354030 309952 354036 309964
rect 354088 309952 354094 310004
rect 265710 309884 265716 309936
rect 265768 309924 265774 309936
rect 332778 309924 332784 309936
rect 265768 309896 332784 309924
rect 265768 309884 265774 309896
rect 332778 309884 332784 309896
rect 332836 309884 332842 309936
rect 260190 309816 260196 309868
rect 260248 309856 260254 309868
rect 332594 309856 332600 309868
rect 260248 309828 332600 309856
rect 260248 309816 260254 309828
rect 332594 309816 332600 309828
rect 332652 309816 332658 309868
rect 291838 309748 291844 309800
rect 291896 309788 291902 309800
rect 298002 309788 298008 309800
rect 291896 309760 298008 309788
rect 291896 309748 291902 309760
rect 298002 309748 298008 309760
rect 298060 309788 298066 309800
rect 341978 309788 341984 309800
rect 298060 309760 341984 309788
rect 298060 309748 298066 309760
rect 341978 309748 341984 309760
rect 342036 309748 342042 309800
rect 375282 309748 375288 309800
rect 375340 309788 375346 309800
rect 414014 309788 414020 309800
rect 375340 309760 414020 309788
rect 375340 309748 375346 309760
rect 414014 309748 414020 309760
rect 414072 309748 414078 309800
rect 304994 309680 305000 309732
rect 305052 309720 305058 309732
rect 305638 309720 305644 309732
rect 305052 309692 305644 309720
rect 305052 309680 305058 309692
rect 305638 309680 305644 309692
rect 305696 309720 305702 309732
rect 347498 309720 347504 309732
rect 305696 309692 347504 309720
rect 305696 309680 305702 309692
rect 347498 309680 347504 309692
rect 347556 309680 347562 309732
rect 298738 309612 298744 309664
rect 298796 309652 298802 309664
rect 300486 309652 300492 309664
rect 298796 309624 300492 309652
rect 298796 309612 298802 309624
rect 300486 309612 300492 309624
rect 300544 309652 300550 309664
rect 333422 309652 333428 309664
rect 300544 309624 333428 309652
rect 300544 309612 300550 309624
rect 333422 309612 333428 309624
rect 333480 309612 333486 309664
rect 321278 309544 321284 309596
rect 321336 309584 321342 309596
rect 346026 309584 346032 309596
rect 321336 309556 346032 309584
rect 321336 309544 321342 309556
rect 346026 309544 346032 309556
rect 346084 309544 346090 309596
rect 328454 309476 328460 309528
rect 328512 309516 328518 309528
rect 328638 309516 328644 309528
rect 328512 309488 328644 309516
rect 328512 309476 328518 309488
rect 328638 309476 328644 309488
rect 328696 309476 328702 309528
rect 296070 309136 296076 309188
rect 296128 309176 296134 309188
rect 307018 309176 307024 309188
rect 296128 309148 307024 309176
rect 296128 309136 296134 309148
rect 307018 309136 307024 309148
rect 307076 309176 307082 309188
rect 307478 309176 307484 309188
rect 307076 309148 307484 309176
rect 307076 309136 307082 309148
rect 307478 309136 307484 309148
rect 307536 309136 307542 309188
rect 270402 309068 270408 309120
rect 270460 309108 270466 309120
rect 292758 309108 292764 309120
rect 270460 309080 292764 309108
rect 270460 309068 270466 309080
rect 292758 309068 292764 309080
rect 292816 309068 292822 309120
rect 302510 309068 302516 309120
rect 302568 309108 302574 309120
rect 303062 309108 303068 309120
rect 302568 309080 303068 309108
rect 302568 309068 302574 309080
rect 303062 309068 303068 309080
rect 303120 309068 303126 309120
rect 334894 309108 334900 309120
rect 306346 309080 334900 309108
rect 303982 309040 303988 309052
rect 296686 309012 303988 309040
rect 277118 308796 277124 308848
rect 277176 308836 277182 308848
rect 296686 308836 296714 309012
rect 303982 309000 303988 309012
rect 304040 309040 304046 309052
rect 306346 309040 306374 309080
rect 334894 309068 334900 309080
rect 334952 309068 334958 309120
rect 304040 309012 306374 309040
rect 304040 309000 304046 309012
rect 306834 309000 306840 309052
rect 306892 309040 306898 309052
rect 307202 309040 307208 309052
rect 306892 309012 307208 309040
rect 306892 309000 306898 309012
rect 307202 309000 307208 309012
rect 307260 309000 307266 309052
rect 309778 309000 309784 309052
rect 309836 309040 309842 309052
rect 337562 309040 337568 309052
rect 309836 309012 337568 309040
rect 309836 309000 309842 309012
rect 337562 309000 337568 309012
rect 337620 309000 337626 309052
rect 307478 308932 307484 308984
rect 307536 308972 307542 308984
rect 368290 308972 368296 308984
rect 307536 308944 368296 308972
rect 307536 308932 307542 308944
rect 368290 308932 368296 308944
rect 368348 308932 368354 308984
rect 307202 308864 307208 308916
rect 307260 308904 307266 308916
rect 366450 308904 366456 308916
rect 307260 308876 366456 308904
rect 307260 308864 307266 308876
rect 366450 308864 366456 308876
rect 366508 308864 366514 308916
rect 277176 308808 296714 308836
rect 277176 308796 277182 308808
rect 305454 308796 305460 308848
rect 305512 308836 305518 308848
rect 306098 308836 306104 308848
rect 305512 308808 306104 308836
rect 305512 308796 305518 308808
rect 306098 308796 306104 308808
rect 306156 308836 306162 308848
rect 363598 308836 363604 308848
rect 306156 308808 363604 308836
rect 306156 308796 306162 308808
rect 363598 308796 363604 308808
rect 363656 308796 363662 308848
rect 293402 308728 293408 308780
rect 293460 308768 293466 308780
rect 310514 308768 310520 308780
rect 293460 308740 310520 308768
rect 293460 308728 293466 308740
rect 310514 308728 310520 308740
rect 310572 308768 310578 308780
rect 365806 308768 365812 308780
rect 310572 308740 365812 308768
rect 310572 308728 310578 308740
rect 365806 308728 365812 308740
rect 365864 308728 365870 308780
rect 300394 308660 300400 308712
rect 300452 308700 300458 308712
rect 305546 308700 305552 308712
rect 300452 308672 305552 308700
rect 300452 308660 300458 308672
rect 305546 308660 305552 308672
rect 305604 308700 305610 308712
rect 360838 308700 360844 308712
rect 305604 308672 360844 308700
rect 305604 308660 305610 308672
rect 360838 308660 360844 308672
rect 360896 308660 360902 308712
rect 303062 308592 303068 308644
rect 303120 308632 303126 308644
rect 352834 308632 352840 308644
rect 303120 308604 352840 308632
rect 303120 308592 303126 308604
rect 352834 308592 352840 308604
rect 352892 308592 352898 308644
rect 296990 308524 296996 308576
rect 297048 308564 297054 308576
rect 339034 308564 339040 308576
rect 297048 308536 339040 308564
rect 297048 308524 297054 308536
rect 339034 308524 339040 308536
rect 339092 308524 339098 308576
rect 213546 308456 213552 308508
rect 213604 308496 213610 308508
rect 269574 308496 269580 308508
rect 213604 308468 269580 308496
rect 213604 308456 213610 308468
rect 269574 308456 269580 308468
rect 269632 308496 269638 308508
rect 270402 308496 270408 308508
rect 269632 308468 270408 308496
rect 269632 308456 269638 308468
rect 270402 308456 270408 308468
rect 270460 308456 270466 308508
rect 302602 308456 302608 308508
rect 302660 308496 302666 308508
rect 343174 308496 343180 308508
rect 302660 308468 343180 308496
rect 302660 308456 302666 308468
rect 343174 308456 343180 308468
rect 343232 308456 343238 308508
rect 221918 308388 221924 308440
rect 221976 308428 221982 308440
rect 301406 308428 301412 308440
rect 221976 308400 301412 308428
rect 221976 308388 221982 308400
rect 301406 308388 301412 308400
rect 301464 308388 301470 308440
rect 303614 308388 303620 308440
rect 303672 308428 303678 308440
rect 364886 308428 364892 308440
rect 303672 308400 364892 308428
rect 303672 308388 303678 308400
rect 364886 308388 364892 308400
rect 364944 308388 364950 308440
rect 286778 308320 286784 308372
rect 286836 308360 286842 308372
rect 327534 308360 327540 308372
rect 286836 308332 327540 308360
rect 286836 308320 286842 308332
rect 327534 308320 327540 308332
rect 327592 308320 327598 308372
rect 296990 308252 296996 308304
rect 297048 308292 297054 308304
rect 297450 308292 297456 308304
rect 297048 308264 297456 308292
rect 297048 308252 297054 308264
rect 297450 308252 297456 308264
rect 297508 308252 297514 308304
rect 307478 308252 307484 308304
rect 307536 308292 307542 308304
rect 367922 308292 367928 308304
rect 307536 308264 367928 308292
rect 307536 308252 307542 308264
rect 367922 308252 367928 308264
rect 367980 308252 367986 308304
rect 315114 308184 315120 308236
rect 315172 308224 315178 308236
rect 315482 308224 315488 308236
rect 315172 308196 315488 308224
rect 315172 308184 315178 308196
rect 315482 308184 315488 308196
rect 315540 308224 315546 308236
rect 389358 308224 389364 308236
rect 315540 308196 389364 308224
rect 315540 308184 315546 308196
rect 389358 308184 389364 308196
rect 389416 308184 389422 308236
rect 284018 307844 284024 307896
rect 284076 307884 284082 307896
rect 308582 307884 308588 307896
rect 284076 307856 308588 307884
rect 284076 307844 284082 307856
rect 308582 307844 308588 307856
rect 308640 307884 308646 307896
rect 308950 307884 308956 307896
rect 308640 307856 308956 307884
rect 308640 307844 308646 307856
rect 308950 307844 308956 307856
rect 309008 307844 309014 307896
rect 210602 307776 210608 307828
rect 210660 307816 210666 307828
rect 296162 307816 296168 307828
rect 210660 307788 296168 307816
rect 210660 307776 210666 307788
rect 296162 307776 296168 307788
rect 296220 307776 296226 307828
rect 304442 307776 304448 307828
rect 304500 307816 304506 307828
rect 306742 307816 306748 307828
rect 304500 307788 306748 307816
rect 304500 307776 304506 307788
rect 306742 307776 306748 307788
rect 306800 307816 306806 307828
rect 307478 307816 307484 307828
rect 306800 307788 307484 307816
rect 306800 307776 306806 307788
rect 307478 307776 307484 307788
rect 307536 307776 307542 307828
rect 261938 307708 261944 307760
rect 261996 307748 262002 307760
rect 287790 307748 287796 307760
rect 261996 307720 287796 307748
rect 261996 307708 262002 307720
rect 287790 307708 287796 307720
rect 287848 307708 287854 307760
rect 298370 307708 298376 307760
rect 298428 307748 298434 307760
rect 299198 307748 299204 307760
rect 298428 307720 299204 307748
rect 298428 307708 298434 307720
rect 299198 307708 299204 307720
rect 299256 307708 299262 307760
rect 299566 307708 299572 307760
rect 299624 307748 299630 307760
rect 300486 307748 300492 307760
rect 299624 307720 300492 307748
rect 299624 307708 299630 307720
rect 300486 307708 300492 307720
rect 300544 307708 300550 307760
rect 301038 307708 301044 307760
rect 301096 307748 301102 307760
rect 301590 307748 301596 307760
rect 301096 307720 301596 307748
rect 301096 307708 301102 307720
rect 301590 307708 301596 307720
rect 301648 307708 301654 307760
rect 304258 307708 304264 307760
rect 304316 307748 304322 307760
rect 305822 307748 305828 307760
rect 304316 307720 305828 307748
rect 304316 307708 304322 307720
rect 305822 307708 305828 307720
rect 305880 307708 305886 307760
rect 314286 307708 314292 307760
rect 314344 307748 314350 307760
rect 394970 307748 394976 307760
rect 314344 307720 394976 307748
rect 314344 307708 314350 307720
rect 394970 307708 394976 307720
rect 395028 307748 395034 307760
rect 395982 307748 395988 307760
rect 395028 307720 395988 307748
rect 395028 307708 395034 307720
rect 395982 307708 395988 307720
rect 396040 307708 396046 307760
rect 280982 307640 280988 307692
rect 281040 307680 281046 307692
rect 301774 307680 301780 307692
rect 281040 307652 301780 307680
rect 281040 307640 281046 307652
rect 301774 307640 301780 307652
rect 301832 307680 301838 307692
rect 360654 307680 360660 307692
rect 301832 307652 360660 307680
rect 301832 307640 301838 307652
rect 360654 307640 360660 307652
rect 360712 307640 360718 307692
rect 260742 307572 260748 307624
rect 260800 307612 260806 307624
rect 283190 307612 283196 307624
rect 260800 307584 283196 307612
rect 260800 307572 260806 307584
rect 283190 307572 283196 307584
rect 283248 307572 283254 307624
rect 303522 307572 303528 307624
rect 303580 307612 303586 307624
rect 304534 307612 304540 307624
rect 303580 307584 304540 307612
rect 303580 307572 303586 307584
rect 304534 307572 304540 307584
rect 304592 307572 304598 307624
rect 363782 307612 363788 307624
rect 306346 307584 363788 307612
rect 301498 307504 301504 307556
rect 301556 307544 301562 307556
rect 302418 307544 302424 307556
rect 301556 307516 302424 307544
rect 301556 307504 301562 307516
rect 302418 307504 302424 307516
rect 302476 307544 302482 307556
rect 306346 307544 306374 307584
rect 363782 307572 363788 307584
rect 363840 307572 363846 307624
rect 302476 307516 306374 307544
rect 302476 307504 302482 307516
rect 320634 307504 320640 307556
rect 320692 307544 320698 307556
rect 381722 307544 381728 307556
rect 320692 307516 381728 307544
rect 320692 307504 320698 307516
rect 381722 307504 381728 307516
rect 381780 307504 381786 307556
rect 299198 307436 299204 307488
rect 299256 307476 299262 307488
rect 356790 307476 356796 307488
rect 299256 307448 356796 307476
rect 299256 307436 299262 307448
rect 356790 307436 356796 307448
rect 356848 307436 356854 307488
rect 274358 307368 274364 307420
rect 274416 307408 274422 307420
rect 302234 307408 302240 307420
rect 274416 307380 302240 307408
rect 274416 307368 274422 307380
rect 302234 307368 302240 307380
rect 302292 307368 302298 307420
rect 312170 307368 312176 307420
rect 312228 307408 312234 307420
rect 370590 307408 370596 307420
rect 312228 307380 370596 307408
rect 312228 307368 312234 307380
rect 370590 307368 370596 307380
rect 370648 307368 370654 307420
rect 275922 307300 275928 307352
rect 275980 307340 275986 307352
rect 303890 307340 303896 307352
rect 275980 307312 303896 307340
rect 275980 307300 275986 307312
rect 303890 307300 303896 307312
rect 303948 307340 303954 307352
rect 358078 307340 358084 307352
rect 303948 307312 358084 307340
rect 303948 307300 303954 307312
rect 358078 307300 358084 307312
rect 358136 307300 358142 307352
rect 300302 307232 300308 307284
rect 300360 307272 300366 307284
rect 301130 307272 301136 307284
rect 300360 307244 301136 307272
rect 300360 307232 300366 307244
rect 301130 307232 301136 307244
rect 301188 307232 301194 307284
rect 301590 307232 301596 307284
rect 301648 307272 301654 307284
rect 344554 307272 344560 307284
rect 301648 307244 344560 307272
rect 301648 307232 301654 307244
rect 344554 307232 344560 307244
rect 344612 307232 344618 307284
rect 202506 307164 202512 307216
rect 202564 307204 202570 307216
rect 261938 307204 261944 307216
rect 202564 307176 261944 307204
rect 202564 307164 202570 307176
rect 261938 307164 261944 307176
rect 261996 307164 262002 307216
rect 300486 307164 300492 307216
rect 300544 307204 300550 307216
rect 341886 307204 341892 307216
rect 300544 307176 341892 307204
rect 300544 307164 300550 307176
rect 341886 307164 341892 307176
rect 341944 307164 341950 307216
rect 217594 307096 217600 307148
rect 217652 307136 217658 307148
rect 300026 307136 300032 307148
rect 217652 307108 300032 307136
rect 217652 307096 217658 307108
rect 300026 307096 300032 307108
rect 300084 307136 300090 307148
rect 300084 307108 301084 307136
rect 300084 307096 300090 307108
rect 209406 307028 209412 307080
rect 209464 307068 209470 307080
rect 297726 307068 297732 307080
rect 209464 307040 297732 307068
rect 209464 307028 209470 307040
rect 297726 307028 297732 307040
rect 297784 307028 297790 307080
rect 301056 306864 301084 307108
rect 305362 307096 305368 307148
rect 305420 307136 305426 307148
rect 345750 307136 345756 307148
rect 305420 307108 345756 307136
rect 305420 307096 305426 307108
rect 345750 307096 345756 307108
rect 345808 307096 345814 307148
rect 301130 307028 301136 307080
rect 301188 307068 301194 307080
rect 336182 307068 336188 307080
rect 301188 307040 336188 307068
rect 301188 307028 301194 307040
rect 336182 307028 336188 307040
rect 336240 307028 336246 307080
rect 395982 307028 395988 307080
rect 396040 307068 396046 307080
rect 409874 307068 409880 307080
rect 396040 307040 409880 307068
rect 396040 307028 396046 307040
rect 409874 307028 409880 307040
rect 409932 307028 409938 307080
rect 329374 306960 329380 307012
rect 329432 307000 329438 307012
rect 332778 307000 332784 307012
rect 329432 306972 332784 307000
rect 329432 306960 329438 306972
rect 332778 306960 332784 306972
rect 332836 306960 332842 307012
rect 302234 306892 302240 306944
rect 302292 306932 302298 306944
rect 338942 306932 338948 306944
rect 302292 306904 338948 306932
rect 302292 306892 302298 306904
rect 338942 306892 338948 306904
rect 339000 306892 339006 306944
rect 336274 306864 336280 306876
rect 301056 306836 336280 306864
rect 336274 306824 336280 306836
rect 336332 306824 336338 306876
rect 280062 306348 280068 306400
rect 280120 306388 280126 306400
rect 303522 306388 303528 306400
rect 280120 306360 303528 306388
rect 280120 306348 280126 306360
rect 303522 306348 303528 306360
rect 303580 306348 303586 306400
rect 266078 306280 266084 306332
rect 266136 306320 266142 306332
rect 285950 306320 285956 306332
rect 266136 306292 285956 306320
rect 266136 306280 266142 306292
rect 285950 306280 285956 306292
rect 286008 306280 286014 306332
rect 297818 306280 297824 306332
rect 297876 306320 297882 306332
rect 359182 306320 359188 306332
rect 297876 306292 359188 306320
rect 297876 306280 297882 306292
rect 359182 306280 359188 306292
rect 359240 306280 359246 306332
rect 291562 306212 291568 306264
rect 291620 306252 291626 306264
rect 351178 306252 351184 306264
rect 291620 306224 351184 306252
rect 291620 306212 291626 306224
rect 351178 306212 351184 306224
rect 351236 306212 351242 306264
rect 295610 306144 295616 306196
rect 295668 306184 295674 306196
rect 355778 306184 355784 306196
rect 295668 306156 355784 306184
rect 295668 306144 295674 306156
rect 355778 306144 355784 306156
rect 355836 306144 355842 306196
rect 294782 306076 294788 306128
rect 294840 306116 294846 306128
rect 352742 306116 352748 306128
rect 294840 306088 352748 306116
rect 294840 306076 294846 306088
rect 352742 306076 352748 306088
rect 352800 306076 352806 306128
rect 295058 306008 295064 306060
rect 295116 306048 295122 306060
rect 348418 306048 348424 306060
rect 295116 306020 348424 306048
rect 295116 306008 295122 306020
rect 348418 306008 348424 306020
rect 348476 306008 348482 306060
rect 294414 305940 294420 305992
rect 294472 305980 294478 305992
rect 347314 305980 347320 305992
rect 294472 305952 347320 305980
rect 294472 305940 294478 305952
rect 347314 305940 347320 305952
rect 347372 305940 347378 305992
rect 210326 305872 210332 305924
rect 210384 305912 210390 305924
rect 266078 305912 266084 305924
rect 210384 305884 266084 305912
rect 210384 305872 210390 305884
rect 266078 305872 266084 305884
rect 266136 305872 266142 305924
rect 295058 305912 295064 305924
rect 291764 305884 295064 305912
rect 217410 305804 217416 305856
rect 217468 305844 217474 305856
rect 291562 305844 291568 305856
rect 217468 305816 291568 305844
rect 217468 305804 217474 305816
rect 291562 305804 291568 305816
rect 291620 305804 291626 305856
rect 217502 305736 217508 305788
rect 217560 305776 217566 305788
rect 291764 305776 291792 305884
rect 295058 305872 295064 305884
rect 295116 305872 295122 305924
rect 296898 305912 296904 305924
rect 296686 305884 296904 305912
rect 296686 305844 296714 305884
rect 296898 305872 296904 305884
rect 296956 305912 296962 305924
rect 349798 305912 349804 305924
rect 296956 305884 349804 305912
rect 296956 305872 296962 305884
rect 349798 305872 349804 305884
rect 349856 305872 349862 305924
rect 217560 305748 291792 305776
rect 294892 305816 296714 305844
rect 217560 305736 217566 305748
rect 214466 305668 214472 305720
rect 214524 305708 214530 305720
rect 294782 305708 294788 305720
rect 214524 305680 294788 305708
rect 214524 305668 214530 305680
rect 294782 305668 294788 305680
rect 294840 305668 294846 305720
rect 214650 305600 214656 305652
rect 214708 305640 214714 305652
rect 294892 305640 294920 305816
rect 304350 305804 304356 305856
rect 304408 305844 304414 305856
rect 316218 305844 316224 305856
rect 304408 305816 316224 305844
rect 304408 305804 304414 305816
rect 316218 305804 316224 305816
rect 316276 305844 316282 305856
rect 316954 305844 316960 305856
rect 316276 305816 316960 305844
rect 316276 305804 316282 305816
rect 316954 305804 316960 305816
rect 317012 305804 317018 305856
rect 319622 305804 319628 305856
rect 319680 305844 319686 305856
rect 372154 305844 372160 305856
rect 319680 305816 372160 305844
rect 319680 305804 319686 305816
rect 372154 305804 372160 305816
rect 372212 305804 372218 305856
rect 296162 305736 296168 305788
rect 296220 305776 296226 305788
rect 336366 305776 336372 305788
rect 296220 305748 336372 305776
rect 296220 305736 296226 305748
rect 336366 305736 336372 305748
rect 336424 305736 336430 305788
rect 214708 305612 294920 305640
rect 214708 305600 214714 305612
rect 300854 305600 300860 305652
rect 300912 305640 300918 305652
rect 340230 305640 340236 305652
rect 300912 305612 340236 305640
rect 300912 305600 300918 305612
rect 340230 305600 340236 305612
rect 340288 305600 340294 305652
rect 285030 305532 285036 305584
rect 285088 305572 285094 305584
rect 327718 305572 327724 305584
rect 285088 305544 327724 305572
rect 285088 305532 285094 305544
rect 327718 305532 327724 305544
rect 327776 305532 327782 305584
rect 287514 305464 287520 305516
rect 287572 305504 287578 305516
rect 330478 305504 330484 305516
rect 287572 305476 330484 305504
rect 287572 305464 287578 305476
rect 330478 305464 330484 305476
rect 330536 305464 330542 305516
rect 316954 305396 316960 305448
rect 317012 305436 317018 305448
rect 353938 305436 353944 305448
rect 317012 305408 353944 305436
rect 317012 305396 317018 305408
rect 353938 305396 353944 305408
rect 353996 305396 354002 305448
rect 330570 305368 330576 305380
rect 296686 305340 330576 305368
rect 263870 305260 263876 305312
rect 263928 305300 263934 305312
rect 264698 305300 264704 305312
rect 263928 305272 264704 305300
rect 263928 305260 263934 305272
rect 264698 305260 264704 305272
rect 264756 305260 264762 305312
rect 291470 305260 291476 305312
rect 291528 305300 291534 305312
rect 292022 305300 292028 305312
rect 291528 305272 292028 305300
rect 291528 305260 291534 305272
rect 292022 305260 292028 305272
rect 292080 305300 292086 305312
rect 296686 305300 296714 305340
rect 330570 305328 330576 305340
rect 330628 305328 330634 305380
rect 292080 305272 296714 305300
rect 292080 305260 292086 305272
rect 209222 305124 209228 305176
rect 209280 305164 209286 305176
rect 266998 305164 267004 305176
rect 209280 305136 267004 305164
rect 209280 305124 209286 305136
rect 266998 305124 267004 305136
rect 267056 305164 267062 305176
rect 267056 305136 267734 305164
rect 267056 305124 267062 305136
rect 205542 305056 205548 305108
rect 205600 305096 205606 305108
rect 265710 305096 265716 305108
rect 205600 305068 265716 305096
rect 205600 305056 205606 305068
rect 265710 305056 265716 305068
rect 265768 305056 265774 305108
rect 204070 304988 204076 305040
rect 204128 305028 204134 305040
rect 263870 305028 263876 305040
rect 204128 305000 263876 305028
rect 204128 304988 204134 305000
rect 263870 304988 263876 305000
rect 263928 304988 263934 305040
rect 267706 304960 267734 305136
rect 287514 304988 287520 305040
rect 287572 305028 287578 305040
rect 287790 305028 287796 305040
rect 287572 305000 287796 305028
rect 287572 304988 287578 305000
rect 287790 304988 287796 305000
rect 287848 304988 287854 305040
rect 291930 304988 291936 305040
rect 291988 305028 291994 305040
rect 295610 305028 295616 305040
rect 291988 305000 295616 305028
rect 291988 304988 291994 305000
rect 295610 304988 295616 305000
rect 295668 304988 295674 305040
rect 297358 304988 297364 305040
rect 297416 305028 297422 305040
rect 297818 305028 297824 305040
rect 297416 305000 297824 305028
rect 297416 304988 297422 305000
rect 297818 304988 297824 305000
rect 297876 304988 297882 305040
rect 299934 304988 299940 305040
rect 299992 305028 299998 305040
rect 300854 305028 300860 305040
rect 299992 305000 300860 305028
rect 299992 304988 299998 305000
rect 300854 304988 300860 305000
rect 300912 304988 300918 305040
rect 285858 304960 285864 304972
rect 267706 304932 285864 304960
rect 285858 304920 285864 304932
rect 285916 304920 285922 304972
rect 317598 304920 317604 304972
rect 317656 304960 317662 304972
rect 330662 304960 330668 304972
rect 317656 304932 330668 304960
rect 317656 304920 317662 304932
rect 330662 304920 330668 304932
rect 330720 304920 330726 304972
rect 281074 304852 281080 304904
rect 281132 304892 281138 304904
rect 294046 304892 294052 304904
rect 281132 304864 294052 304892
rect 281132 304852 281138 304864
rect 294046 304852 294052 304864
rect 294104 304892 294110 304904
rect 354398 304892 354404 304904
rect 294104 304864 354404 304892
rect 294104 304852 294110 304864
rect 354398 304852 354404 304864
rect 354456 304852 354462 304904
rect 303154 304784 303160 304836
rect 303212 304824 303218 304836
rect 314654 304824 314660 304836
rect 303212 304796 314660 304824
rect 303212 304784 303218 304796
rect 314654 304784 314660 304796
rect 314712 304824 314718 304836
rect 315022 304824 315028 304836
rect 314712 304796 315028 304824
rect 314712 304784 314718 304796
rect 315022 304784 315028 304796
rect 315080 304784 315086 304836
rect 319806 304784 319812 304836
rect 319864 304824 319870 304836
rect 381814 304824 381820 304836
rect 319864 304796 381820 304824
rect 319864 304784 319870 304796
rect 381814 304784 381820 304796
rect 381872 304784 381878 304836
rect 311986 304716 311992 304768
rect 312044 304756 312050 304768
rect 373442 304756 373448 304768
rect 312044 304728 373448 304756
rect 312044 304716 312050 304728
rect 373442 304716 373448 304728
rect 373500 304716 373506 304768
rect 301774 304648 301780 304700
rect 301832 304688 301838 304700
rect 310606 304688 310612 304700
rect 301832 304660 310612 304688
rect 301832 304648 301838 304660
rect 310606 304648 310612 304660
rect 310664 304688 310670 304700
rect 370498 304688 370504 304700
rect 310664 304660 370504 304688
rect 310664 304648 310670 304660
rect 370498 304648 370504 304660
rect 370556 304648 370562 304700
rect 295334 304580 295340 304632
rect 295392 304620 295398 304632
rect 295518 304620 295524 304632
rect 295392 304592 295524 304620
rect 295392 304580 295398 304592
rect 295518 304580 295524 304592
rect 295576 304620 295582 304632
rect 355134 304620 355140 304632
rect 295576 304592 355140 304620
rect 295576 304580 295582 304592
rect 355134 304580 355140 304592
rect 355192 304580 355198 304632
rect 341610 304552 341616 304564
rect 296686 304524 341616 304552
rect 282638 304444 282644 304496
rect 282696 304484 282702 304496
rect 294874 304484 294880 304496
rect 282696 304456 294880 304484
rect 282696 304444 282702 304456
rect 294874 304444 294880 304456
rect 294932 304484 294938 304496
rect 296686 304484 296714 304524
rect 341610 304512 341616 304524
rect 341668 304512 341674 304564
rect 334802 304484 334808 304496
rect 294932 304456 296714 304484
rect 306346 304456 334808 304484
rect 294932 304444 294938 304456
rect 288158 304376 288164 304428
rect 288216 304416 288222 304428
rect 296438 304416 296444 304428
rect 288216 304388 296444 304416
rect 288216 304376 288222 304388
rect 296438 304376 296444 304388
rect 296496 304416 296502 304428
rect 306346 304416 306374 304456
rect 334802 304444 334808 304456
rect 334860 304444 334866 304496
rect 296496 304388 306374 304416
rect 296496 304376 296502 304388
rect 309502 304376 309508 304428
rect 309560 304416 309566 304428
rect 343082 304416 343088 304428
rect 309560 304388 343088 304416
rect 309560 304376 309566 304388
rect 343082 304376 343088 304388
rect 343140 304376 343146 304428
rect 294782 304308 294788 304360
rect 294840 304348 294846 304360
rect 311986 304348 311992 304360
rect 294840 304320 311992 304348
rect 294840 304308 294846 304320
rect 311986 304308 311992 304320
rect 312044 304308 312050 304360
rect 314930 304308 314936 304360
rect 314988 304348 314994 304360
rect 315298 304348 315304 304360
rect 314988 304320 315304 304348
rect 314988 304308 314994 304320
rect 315298 304308 315304 304320
rect 315356 304348 315362 304360
rect 347130 304348 347136 304360
rect 315356 304320 347136 304348
rect 315356 304308 315362 304320
rect 347130 304308 347136 304320
rect 347188 304308 347194 304360
rect 286686 304240 286692 304292
rect 286744 304280 286750 304292
rect 317598 304280 317604 304292
rect 286744 304252 317604 304280
rect 286744 304240 286750 304252
rect 317598 304240 317604 304252
rect 317656 304240 317662 304292
rect 320726 304240 320732 304292
rect 320784 304280 320790 304292
rect 321278 304280 321284 304292
rect 320784 304252 321284 304280
rect 320784 304240 320790 304252
rect 321278 304240 321284 304252
rect 321336 304240 321342 304292
rect 314654 304172 314660 304224
rect 314712 304212 314718 304224
rect 387794 304212 387800 304224
rect 314712 304184 387800 304212
rect 314712 304172 314718 304184
rect 387794 304172 387800 304184
rect 387852 304172 387858 304224
rect 309502 303764 309508 303816
rect 309560 303804 309566 303816
rect 309962 303804 309968 303816
rect 309560 303776 309968 303804
rect 309560 303764 309566 303776
rect 309962 303764 309968 303776
rect 310020 303764 310026 303816
rect 270310 303628 270316 303680
rect 270368 303668 270374 303680
rect 313274 303668 313280 303680
rect 270368 303640 313280 303668
rect 270368 303628 270374 303640
rect 313274 303628 313280 303640
rect 313332 303628 313338 303680
rect 269022 303560 269028 303612
rect 269080 303600 269086 303612
rect 287422 303600 287428 303612
rect 269080 303572 287428 303600
rect 269080 303560 269086 303572
rect 287422 303560 287428 303572
rect 287480 303560 287486 303612
rect 303430 303560 303436 303612
rect 303488 303600 303494 303612
rect 369026 303600 369032 303612
rect 303488 303572 369032 303600
rect 303488 303560 303494 303572
rect 369026 303560 369032 303572
rect 369084 303560 369090 303612
rect 365714 303532 365720 303544
rect 301976 303504 365720 303532
rect 301976 303476 302004 303504
rect 365714 303492 365720 303504
rect 365772 303492 365778 303544
rect 286318 303424 286324 303476
rect 286376 303464 286382 303476
rect 301958 303464 301964 303476
rect 286376 303436 301964 303464
rect 286376 303424 286382 303436
rect 301958 303424 301964 303436
rect 302016 303424 302022 303476
rect 302786 303424 302792 303476
rect 302844 303464 302850 303476
rect 364702 303464 364708 303476
rect 302844 303436 364708 303464
rect 302844 303424 302850 303436
rect 364702 303424 364708 303436
rect 364760 303424 364766 303476
rect 299382 303356 299388 303408
rect 299440 303396 299446 303408
rect 359366 303396 359372 303408
rect 299440 303368 359372 303396
rect 299440 303356 299446 303368
rect 359366 303356 359372 303368
rect 359424 303356 359430 303408
rect 288066 303288 288072 303340
rect 288124 303328 288130 303340
rect 300946 303328 300952 303340
rect 288124 303300 300952 303328
rect 288124 303288 288130 303300
rect 300946 303288 300952 303300
rect 301004 303288 301010 303340
rect 307662 303288 307668 303340
rect 307720 303328 307726 303340
rect 331858 303328 331864 303340
rect 307720 303300 331864 303328
rect 307720 303288 307726 303300
rect 331858 303288 331864 303300
rect 331916 303288 331922 303340
rect 288342 303220 288348 303272
rect 288400 303260 288406 303272
rect 300762 303260 300768 303272
rect 288400 303232 300768 303260
rect 288400 303220 288406 303232
rect 300762 303220 300768 303232
rect 300820 303260 300826 303272
rect 360378 303260 360384 303272
rect 300820 303232 360384 303260
rect 300820 303220 300826 303232
rect 360378 303220 360384 303232
rect 360436 303220 360442 303272
rect 298278 303152 298284 303204
rect 298336 303192 298342 303204
rect 356698 303192 356704 303204
rect 298336 303164 356704 303192
rect 298336 303152 298342 303164
rect 356698 303152 356704 303164
rect 356756 303152 356762 303204
rect 279326 303084 279332 303136
rect 279384 303124 279390 303136
rect 299842 303124 299848 303136
rect 279384 303096 299848 303124
rect 279384 303084 279390 303096
rect 299842 303084 299848 303096
rect 299900 303124 299906 303136
rect 334710 303124 334716 303136
rect 299900 303096 334716 303124
rect 299900 303084 299906 303096
rect 334710 303084 334716 303096
rect 334768 303084 334774 303136
rect 299658 303016 299664 303068
rect 299716 303056 299722 303068
rect 352650 303056 352656 303068
rect 299716 303028 352656 303056
rect 299716 303016 299722 303028
rect 352650 303016 352656 303028
rect 352708 303016 352714 303068
rect 205358 302948 205364 303000
rect 205416 302988 205422 303000
rect 269022 302988 269028 303000
rect 205416 302960 269028 302988
rect 205416 302948 205422 302960
rect 269022 302948 269028 302960
rect 269080 302948 269086 303000
rect 301130 302948 301136 303000
rect 301188 302988 301194 303000
rect 349890 302988 349896 303000
rect 301188 302960 349896 302988
rect 301188 302948 301194 302960
rect 349890 302948 349896 302960
rect 349948 302948 349954 303000
rect 220262 302880 220268 302932
rect 220320 302920 220326 302932
rect 298186 302920 298192 302932
rect 220320 302892 298192 302920
rect 220320 302880 220326 302892
rect 298186 302880 298192 302892
rect 298244 302920 298250 302932
rect 299382 302920 299388 302932
rect 298244 302892 299388 302920
rect 298244 302880 298250 302892
rect 299382 302880 299388 302892
rect 299440 302880 299446 302932
rect 300946 302880 300952 302932
rect 301004 302920 301010 302932
rect 348602 302920 348608 302932
rect 301004 302892 348608 302920
rect 301004 302880 301010 302892
rect 348602 302880 348608 302892
rect 348660 302880 348666 302932
rect 395982 302880 395988 302932
rect 396040 302920 396046 302932
rect 565814 302920 565820 302932
rect 396040 302892 565820 302920
rect 396040 302880 396046 302892
rect 565814 302880 565820 302892
rect 565872 302880 565878 302932
rect 299750 302812 299756 302864
rect 299808 302852 299814 302864
rect 341702 302852 341708 302864
rect 299808 302824 341708 302852
rect 299808 302812 299814 302824
rect 341702 302812 341708 302824
rect 341760 302812 341766 302864
rect 303798 302744 303804 302796
rect 303856 302784 303862 302796
rect 304534 302784 304540 302796
rect 303856 302756 304540 302784
rect 303856 302744 303862 302756
rect 304534 302744 304540 302756
rect 304592 302784 304598 302796
rect 337470 302784 337476 302796
rect 304592 302756 337476 302784
rect 304592 302744 304598 302756
rect 337470 302744 337476 302756
rect 337528 302744 337534 302796
rect 321646 302676 321652 302728
rect 321704 302716 321710 302728
rect 322474 302716 322480 302728
rect 321704 302688 322480 302716
rect 321704 302676 321710 302688
rect 322474 302676 322480 302688
rect 322532 302716 322538 302728
rect 383286 302716 383292 302728
rect 322532 302688 383292 302716
rect 322532 302676 322538 302688
rect 383286 302676 383292 302688
rect 383344 302676 383350 302728
rect 213270 302268 213276 302320
rect 213328 302308 213334 302320
rect 259546 302308 259552 302320
rect 213328 302280 259552 302308
rect 213328 302268 213334 302280
rect 259546 302268 259552 302280
rect 259604 302308 259610 302320
rect 260190 302308 260196 302320
rect 259604 302280 260196 302308
rect 259604 302268 259610 302280
rect 260190 302268 260196 302280
rect 260248 302268 260254 302320
rect 202690 302200 202696 302252
rect 202748 302240 202754 302252
rect 262490 302240 262496 302252
rect 202748 302212 262496 302240
rect 202748 302200 202754 302212
rect 262490 302200 262496 302212
rect 262548 302240 262554 302252
rect 262950 302240 262956 302252
rect 262548 302212 262956 302240
rect 262548 302200 262554 302212
rect 262950 302200 262956 302212
rect 263008 302200 263014 302252
rect 299658 302200 299664 302252
rect 299716 302240 299722 302252
rect 300210 302240 300216 302252
rect 299716 302212 300216 302240
rect 299716 302200 299722 302212
rect 300210 302200 300216 302212
rect 300268 302200 300274 302252
rect 302786 302200 302792 302252
rect 302844 302240 302850 302252
rect 303246 302240 303252 302252
rect 302844 302212 303252 302240
rect 302844 302200 302850 302212
rect 303246 302200 303252 302212
rect 303304 302200 303310 302252
rect 264974 302132 264980 302184
rect 265032 302172 265038 302184
rect 266262 302172 266268 302184
rect 265032 302144 266268 302172
rect 265032 302132 265038 302144
rect 266262 302132 266268 302144
rect 266320 302172 266326 302184
rect 287330 302172 287336 302184
rect 266320 302144 287336 302172
rect 266320 302132 266326 302144
rect 287330 302132 287336 302144
rect 287388 302132 287394 302184
rect 321646 302132 321652 302184
rect 321704 302172 321710 302184
rect 394786 302172 394792 302184
rect 321704 302144 394792 302172
rect 321704 302132 321710 302144
rect 394786 302132 394792 302144
rect 394844 302132 394850 302184
rect 296162 302064 296168 302116
rect 296220 302104 296226 302116
rect 296622 302104 296628 302116
rect 296220 302076 296628 302104
rect 296220 302064 296226 302076
rect 296622 302064 296628 302076
rect 296680 302104 296686 302116
rect 358446 302104 358452 302116
rect 296680 302076 358452 302104
rect 296680 302064 296686 302076
rect 358446 302064 358452 302076
rect 358504 302064 358510 302116
rect 300670 301996 300676 302048
rect 300728 302036 300734 302048
rect 360746 302036 360752 302048
rect 300728 302008 360752 302036
rect 300728 301996 300734 302008
rect 360746 301996 360752 302008
rect 360804 301996 360810 302048
rect 300578 301928 300584 301980
rect 300636 301968 300642 301980
rect 359274 301968 359280 301980
rect 300636 301940 359280 301968
rect 300636 301928 300642 301940
rect 359274 301928 359280 301940
rect 359332 301928 359338 301980
rect 312814 301860 312820 301912
rect 312872 301900 312878 301912
rect 312998 301900 313004 301912
rect 312872 301872 313004 301900
rect 312872 301860 312878 301872
rect 312998 301860 313004 301872
rect 313056 301900 313062 301912
rect 372062 301900 372068 301912
rect 313056 301872 372068 301900
rect 313056 301860 313062 301872
rect 372062 301860 372068 301872
rect 372120 301860 372126 301912
rect 293954 301792 293960 301844
rect 294012 301832 294018 301844
rect 294506 301832 294512 301844
rect 294012 301804 294512 301832
rect 294012 301792 294018 301804
rect 294506 301792 294512 301804
rect 294564 301832 294570 301844
rect 351270 301832 351276 301844
rect 294564 301804 351276 301832
rect 294564 301792 294570 301804
rect 351270 301792 351276 301804
rect 351328 301792 351334 301844
rect 295334 301724 295340 301776
rect 295392 301764 295398 301776
rect 295886 301764 295892 301776
rect 295392 301736 295892 301764
rect 295392 301724 295398 301736
rect 295886 301724 295892 301736
rect 295944 301764 295950 301776
rect 352558 301764 352564 301776
rect 295944 301736 352564 301764
rect 295944 301724 295950 301736
rect 352558 301724 352564 301736
rect 352616 301724 352622 301776
rect 344370 301696 344376 301708
rect 296686 301668 344376 301696
rect 286594 301628 286600 301640
rect 277366 301600 286600 301628
rect 262122 301520 262128 301572
rect 262180 301560 262186 301572
rect 275002 301560 275008 301572
rect 262180 301532 275008 301560
rect 262180 301520 262186 301532
rect 275002 301520 275008 301532
rect 275060 301560 275066 301572
rect 277366 301560 277394 301600
rect 286594 301588 286600 301600
rect 286652 301588 286658 301640
rect 288802 301588 288808 301640
rect 288860 301628 288866 301640
rect 289630 301628 289636 301640
rect 288860 301600 289636 301628
rect 288860 301588 288866 301600
rect 289630 301588 289636 301600
rect 289688 301628 289694 301640
rect 296686 301628 296714 301668
rect 344370 301656 344376 301668
rect 344428 301656 344434 301708
rect 289688 301600 296714 301628
rect 289688 301588 289694 301600
rect 297910 301588 297916 301640
rect 297968 301628 297974 301640
rect 348694 301628 348700 301640
rect 297968 301600 348700 301628
rect 297968 301588 297974 301600
rect 348694 301588 348700 301600
rect 348752 301588 348758 301640
rect 275060 301532 277394 301560
rect 275060 301520 275066 301532
rect 283926 301520 283932 301572
rect 283984 301560 283990 301572
rect 293126 301560 293132 301572
rect 283984 301532 293132 301560
rect 283984 301520 283990 301532
rect 293126 301520 293132 301532
rect 293184 301560 293190 301572
rect 293184 301532 296714 301560
rect 293184 301520 293190 301532
rect 207842 301452 207848 301504
rect 207900 301492 207906 301504
rect 264974 301492 264980 301504
rect 207900 301464 264980 301492
rect 207900 301452 207906 301464
rect 264974 301452 264980 301464
rect 265032 301452 265038 301504
rect 296686 301424 296714 301532
rect 299474 301520 299480 301572
rect 299532 301560 299538 301572
rect 300578 301560 300584 301572
rect 299532 301532 300584 301560
rect 299532 301520 299538 301532
rect 300578 301520 300584 301532
rect 300636 301560 300642 301572
rect 348786 301560 348792 301572
rect 300636 301532 348792 301560
rect 300636 301520 300642 301532
rect 348786 301520 348792 301532
rect 348844 301520 348850 301572
rect 321554 301452 321560 301504
rect 321612 301492 321618 301504
rect 322658 301492 322664 301504
rect 321612 301464 322664 301492
rect 321612 301452 321618 301464
rect 322658 301452 322664 301464
rect 322716 301492 322722 301504
rect 381538 301492 381544 301504
rect 322716 301464 381544 301492
rect 322716 301452 322722 301464
rect 381538 301452 381544 301464
rect 381596 301452 381602 301504
rect 336090 301424 336096 301436
rect 296686 301396 336096 301424
rect 336090 301384 336096 301396
rect 336148 301384 336154 301436
rect 255406 301316 255412 301368
rect 255464 301356 255470 301368
rect 256142 301356 256148 301368
rect 255464 301328 256148 301356
rect 255464 301316 255470 301328
rect 256142 301316 256148 301328
rect 256200 301316 256206 301368
rect 263686 301316 263692 301368
rect 263744 301356 263750 301368
rect 264330 301356 264336 301368
rect 263744 301328 264336 301356
rect 263744 301316 263750 301328
rect 264330 301316 264336 301328
rect 264388 301316 264394 301368
rect 197446 300976 197452 301028
rect 197504 301016 197510 301028
rect 255406 301016 255412 301028
rect 197504 300988 255412 301016
rect 197504 300976 197510 300988
rect 255406 300976 255412 300988
rect 255464 300976 255470 301028
rect 202138 300908 202144 300960
rect 202196 300948 202202 300960
rect 261478 300948 261484 300960
rect 202196 300920 261484 300948
rect 202196 300908 202202 300920
rect 261478 300908 261484 300920
rect 261536 300908 261542 300960
rect 204438 300840 204444 300892
rect 204496 300880 204502 300892
rect 263686 300880 263692 300892
rect 204496 300852 263692 300880
rect 204496 300840 204502 300852
rect 263686 300840 263692 300852
rect 263744 300840 263750 300892
rect 255406 300772 255412 300824
rect 255464 300812 255470 300824
rect 255958 300812 255964 300824
rect 255464 300784 255964 300812
rect 255464 300772 255470 300784
rect 255958 300772 255964 300784
rect 256016 300772 256022 300824
rect 262122 300772 262128 300824
rect 262180 300812 262186 300824
rect 286134 300812 286140 300824
rect 262180 300784 286140 300812
rect 262180 300772 262186 300784
rect 286134 300772 286140 300784
rect 286192 300772 286198 300824
rect 291102 300772 291108 300824
rect 291160 300812 291166 300824
rect 367554 300812 367560 300824
rect 291160 300784 367560 300812
rect 291160 300772 291166 300784
rect 367554 300772 367560 300784
rect 367612 300772 367618 300824
rect 265066 300704 265072 300756
rect 265124 300744 265130 300756
rect 265618 300744 265624 300756
rect 265124 300716 265624 300744
rect 265124 300704 265130 300716
rect 265618 300704 265624 300716
rect 265676 300704 265682 300756
rect 306558 300704 306564 300756
rect 306616 300744 306622 300756
rect 307018 300744 307024 300756
rect 306616 300716 307024 300744
rect 306616 300704 306622 300716
rect 307018 300704 307024 300716
rect 307076 300704 307082 300756
rect 335998 300744 336004 300756
rect 311176 300716 336004 300744
rect 305638 300636 305644 300688
rect 305696 300676 305702 300688
rect 307662 300676 307668 300688
rect 305696 300648 307668 300676
rect 305696 300636 305702 300648
rect 307662 300636 307668 300648
rect 307720 300636 307726 300688
rect 303706 300568 303712 300620
rect 303764 300608 303770 300620
rect 304626 300608 304632 300620
rect 303764 300580 304632 300608
rect 303764 300568 303770 300580
rect 304626 300568 304632 300580
rect 304684 300608 304690 300620
rect 311176 300608 311204 300716
rect 335998 300704 336004 300716
rect 336056 300704 336062 300756
rect 369946 300676 369952 300688
rect 304684 300580 311204 300608
rect 311268 300648 369952 300676
rect 304684 300568 304690 300580
rect 307110 300500 307116 300552
rect 307168 300540 307174 300552
rect 307662 300540 307668 300552
rect 307168 300512 307668 300540
rect 307168 300500 307174 300512
rect 307662 300500 307668 300512
rect 307720 300540 307726 300552
rect 311268 300540 311296 300648
rect 369946 300636 369952 300648
rect 370004 300636 370010 300688
rect 314746 300568 314752 300620
rect 314804 300608 314810 300620
rect 315850 300608 315856 300620
rect 314804 300580 315856 300608
rect 314804 300568 314810 300580
rect 315850 300568 315856 300580
rect 315908 300608 315914 300620
rect 376570 300608 376576 300620
rect 315908 300580 376576 300608
rect 315908 300568 315914 300580
rect 376570 300568 376576 300580
rect 376628 300568 376634 300620
rect 307720 300512 311296 300540
rect 307720 300500 307726 300512
rect 311342 300500 311348 300552
rect 311400 300540 311406 300552
rect 367646 300540 367652 300552
rect 311400 300512 367652 300540
rect 311400 300500 311406 300512
rect 367646 300500 367652 300512
rect 367704 300500 367710 300552
rect 283098 300432 283104 300484
rect 283156 300472 283162 300484
rect 341794 300472 341800 300484
rect 283156 300444 341800 300472
rect 283156 300432 283162 300444
rect 341794 300432 341800 300444
rect 341852 300432 341858 300484
rect 302234 300364 302240 300416
rect 302292 300404 302298 300416
rect 362034 300404 362040 300416
rect 302292 300376 362040 300404
rect 302292 300364 302298 300376
rect 362034 300364 362040 300376
rect 362092 300364 362098 300416
rect 305270 300296 305276 300348
rect 305328 300336 305334 300348
rect 305546 300336 305552 300348
rect 305328 300308 305552 300336
rect 305328 300296 305334 300308
rect 305546 300296 305552 300308
rect 305604 300336 305610 300348
rect 345658 300336 345664 300348
rect 305604 300308 345664 300336
rect 305604 300296 305610 300308
rect 345658 300296 345664 300308
rect 345716 300296 345722 300348
rect 304258 300228 304264 300280
rect 304316 300268 304322 300280
rect 343266 300268 343272 300280
rect 304316 300240 343272 300268
rect 304316 300228 304322 300240
rect 343266 300228 343272 300240
rect 343324 300228 343330 300280
rect 205266 300160 205272 300212
rect 205324 300200 205330 300212
rect 262122 300200 262128 300212
rect 205324 300172 262128 300200
rect 205324 300160 205330 300172
rect 262122 300160 262128 300172
rect 262180 300160 262186 300212
rect 307754 300160 307760 300212
rect 307812 300200 307818 300212
rect 344646 300200 344652 300212
rect 307812 300172 344652 300200
rect 307812 300160 307818 300172
rect 344646 300160 344652 300172
rect 344704 300160 344710 300212
rect 193214 300092 193220 300144
rect 193272 300132 193278 300144
rect 254026 300132 254032 300144
rect 193272 300104 254032 300132
rect 193272 300092 193278 300104
rect 254026 300092 254032 300104
rect 254084 300092 254090 300144
rect 286962 300092 286968 300144
rect 287020 300132 287026 300144
rect 303706 300132 303712 300144
rect 287020 300104 303712 300132
rect 287020 300092 287026 300104
rect 303706 300092 303712 300104
rect 303764 300092 303770 300144
rect 305178 300092 305184 300144
rect 305236 300132 305242 300144
rect 306190 300132 306196 300144
rect 305236 300104 306196 300132
rect 305236 300092 305242 300104
rect 306190 300092 306196 300104
rect 306248 300132 306254 300144
rect 338758 300132 338764 300144
rect 306248 300104 338764 300132
rect 306248 300092 306254 300104
rect 338758 300092 338764 300104
rect 338816 300092 338822 300144
rect 308030 300024 308036 300076
rect 308088 300064 308094 300076
rect 336182 300064 336188 300076
rect 308088 300036 336188 300064
rect 308088 300024 308094 300036
rect 336182 300024 336188 300036
rect 336240 300024 336246 300076
rect 307018 299956 307024 300008
rect 307076 299996 307082 300008
rect 311342 299996 311348 300008
rect 307076 299968 311348 299996
rect 307076 299956 307082 299968
rect 311342 299956 311348 299968
rect 311400 299956 311406 300008
rect 333238 299996 333244 300008
rect 311452 299968 333244 299996
rect 306926 299888 306932 299940
rect 306984 299928 306990 299940
rect 311452 299928 311480 299968
rect 333238 299956 333244 299968
rect 333296 299956 333302 300008
rect 374638 299928 374644 299940
rect 306984 299900 311480 299928
rect 315868 299900 374644 299928
rect 306984 299888 306990 299900
rect 309410 299820 309416 299872
rect 309468 299860 309474 299872
rect 315868 299860 315896 299900
rect 374638 299888 374644 299900
rect 374696 299888 374702 299940
rect 309468 299832 315896 299860
rect 309468 299820 309474 299832
rect 216030 299616 216036 299668
rect 216088 299656 216094 299668
rect 259822 299656 259828 299668
rect 216088 299628 259828 299656
rect 216088 299616 216094 299628
rect 259822 299616 259828 299628
rect 259880 299656 259886 299668
rect 260098 299656 260104 299668
rect 259880 299628 260104 299656
rect 259880 299616 259886 299628
rect 260098 299616 260104 299628
rect 260156 299616 260162 299668
rect 204346 299548 204352 299600
rect 204404 299588 204410 299600
rect 265066 299588 265072 299600
rect 204404 299560 265072 299588
rect 204404 299548 204410 299560
rect 265066 299548 265072 299560
rect 265124 299548 265130 299600
rect 194594 299480 194600 299532
rect 194652 299520 194658 299532
rect 255406 299520 255412 299532
rect 194652 299492 255412 299520
rect 194652 299480 194658 299492
rect 255406 299480 255412 299492
rect 255464 299480 255470 299532
rect 4154 299412 4160 299464
rect 4212 299452 4218 299464
rect 221734 299452 221740 299464
rect 4212 299424 221740 299452
rect 4212 299412 4218 299424
rect 221734 299412 221740 299424
rect 221792 299452 221798 299464
rect 256694 299452 256700 299464
rect 221792 299424 256700 299452
rect 221792 299412 221798 299424
rect 256694 299412 256700 299424
rect 256752 299452 256758 299464
rect 257338 299452 257344 299464
rect 256752 299424 257344 299452
rect 256752 299412 256758 299424
rect 257338 299412 257344 299424
rect 257396 299412 257402 299464
rect 288710 299412 288716 299464
rect 288768 299452 288774 299464
rect 289354 299452 289360 299464
rect 288768 299424 289360 299452
rect 288768 299412 288774 299424
rect 289354 299412 289360 299424
rect 289412 299412 289418 299464
rect 316126 299412 316132 299464
rect 316184 299452 316190 299464
rect 316770 299452 316776 299464
rect 316184 299424 316776 299452
rect 316184 299412 316190 299424
rect 316770 299412 316776 299424
rect 316828 299452 316834 299464
rect 378594 299452 378600 299464
rect 316828 299424 378600 299452
rect 316828 299412 316834 299424
rect 378594 299412 378600 299424
rect 378652 299412 378658 299464
rect 288250 299344 288256 299396
rect 288308 299384 288314 299396
rect 348326 299384 348332 299396
rect 288308 299356 348332 299384
rect 288308 299344 288314 299356
rect 348326 299344 348332 299356
rect 348384 299344 348390 299396
rect 316034 299276 316040 299328
rect 316092 299316 316098 299328
rect 316862 299316 316868 299328
rect 316092 299288 316868 299316
rect 316092 299276 316098 299288
rect 316862 299276 316868 299288
rect 316920 299316 316926 299328
rect 376478 299316 376484 299328
rect 316920 299288 376484 299316
rect 316920 299276 316926 299288
rect 376478 299276 376484 299288
rect 376536 299276 376542 299328
rect 289446 299208 289452 299260
rect 289504 299248 289510 299260
rect 348970 299248 348976 299260
rect 289504 299220 348976 299248
rect 289504 299208 289510 299220
rect 348970 299208 348976 299220
rect 349028 299208 349034 299260
rect 289354 299140 289360 299192
rect 289412 299180 289418 299192
rect 347222 299180 347228 299192
rect 289412 299152 347228 299180
rect 289412 299140 289418 299152
rect 347222 299140 347228 299152
rect 347280 299140 347286 299192
rect 287698 299072 287704 299124
rect 287756 299112 287762 299124
rect 290918 299112 290924 299124
rect 287756 299084 290924 299112
rect 287756 299072 287762 299084
rect 290918 299072 290924 299084
rect 290976 299112 290982 299124
rect 345842 299112 345848 299124
rect 290976 299084 345848 299112
rect 290976 299072 290982 299084
rect 345842 299072 345848 299084
rect 345900 299072 345906 299124
rect 284110 299004 284116 299056
rect 284168 299044 284174 299056
rect 290090 299044 290096 299056
rect 284168 299016 290096 299044
rect 284168 299004 284174 299016
rect 290090 299004 290096 299016
rect 290148 299044 290154 299056
rect 344462 299044 344468 299056
rect 290148 299016 344468 299044
rect 290148 299004 290154 299016
rect 344462 299004 344468 299016
rect 344520 299004 344526 299056
rect 338850 298976 338856 298988
rect 296686 298948 338856 298976
rect 207750 298800 207756 298852
rect 207808 298840 207814 298852
rect 290826 298840 290832 298852
rect 207808 298812 290832 298840
rect 207808 298800 207814 298812
rect 290826 298800 290832 298812
rect 290884 298840 290890 298852
rect 296686 298840 296714 298948
rect 338850 298936 338856 298948
rect 338908 298936 338914 298988
rect 311526 298868 311532 298920
rect 311584 298908 311590 298920
rect 349982 298908 349988 298920
rect 311584 298880 349988 298908
rect 311584 298868 311590 298880
rect 349982 298868 349988 298880
rect 350040 298868 350046 298920
rect 290884 298812 296714 298840
rect 290884 298800 290890 298812
rect 336182 298800 336188 298852
rect 336240 298840 336246 298852
rect 369118 298840 369124 298852
rect 336240 298812 369124 298840
rect 336240 298800 336246 298812
rect 369118 298800 369124 298812
rect 369176 298800 369182 298852
rect 233142 298732 233148 298784
rect 233200 298772 233206 298784
rect 580166 298772 580172 298784
rect 233200 298744 580172 298772
rect 233200 298732 233206 298744
rect 580166 298732 580172 298744
rect 580224 298732 580230 298784
rect 218790 298256 218796 298308
rect 218848 298296 218854 298308
rect 264422 298296 264428 298308
rect 218848 298268 264428 298296
rect 218848 298256 218854 298268
rect 264422 298256 264428 298268
rect 264480 298256 264486 298308
rect 193398 298188 193404 298240
rect 193456 298228 193462 298240
rect 253198 298228 253204 298240
rect 193456 298200 253204 298228
rect 193456 298188 193462 298200
rect 253198 298188 253204 298200
rect 253256 298188 253262 298240
rect 193306 298120 193312 298172
rect 193364 298160 193370 298172
rect 253382 298160 253388 298172
rect 193364 298132 253388 298160
rect 193364 298120 193370 298132
rect 253382 298120 253388 298132
rect 253440 298120 253446 298172
rect 244550 298052 244556 298104
rect 244608 298092 244614 298104
rect 245194 298092 245200 298104
rect 244608 298064 245200 298092
rect 244608 298052 244614 298064
rect 245194 298052 245200 298064
rect 245252 298052 245258 298104
rect 250070 298052 250076 298104
rect 250128 298092 250134 298104
rect 250530 298092 250536 298104
rect 250128 298064 250536 298092
rect 250128 298052 250134 298064
rect 250530 298052 250536 298064
rect 250588 298052 250594 298104
rect 283834 298052 283840 298104
rect 283892 298092 283898 298104
rect 284202 298092 284208 298104
rect 283892 298064 284208 298092
rect 283892 298052 283898 298064
rect 284202 298052 284208 298064
rect 284260 298052 284266 298104
rect 288618 298052 288624 298104
rect 288676 298092 288682 298104
rect 289722 298092 289728 298104
rect 288676 298064 289728 298092
rect 288676 298052 288682 298064
rect 289722 298052 289728 298064
rect 289780 298052 289786 298104
rect 291286 298052 291292 298104
rect 291344 298092 291350 298104
rect 292298 298092 292304 298104
rect 291344 298064 292304 298092
rect 291344 298052 291350 298064
rect 292298 298052 292304 298064
rect 292356 298052 292362 298104
rect 293770 298052 293776 298104
rect 293828 298092 293834 298104
rect 366082 298092 366088 298104
rect 293828 298064 366088 298092
rect 293828 298052 293834 298064
rect 366082 298052 366088 298064
rect 366140 298052 366146 298104
rect 305086 297984 305092 298036
rect 305144 298024 305150 298036
rect 305454 298024 305460 298036
rect 305144 297996 305460 298024
rect 305144 297984 305150 297996
rect 305454 297984 305460 297996
rect 305512 298024 305518 298036
rect 368934 298024 368940 298036
rect 305512 297996 368940 298024
rect 305512 297984 305518 297996
rect 368934 297984 368940 297996
rect 368992 297984 368998 298036
rect 309318 297916 309324 297968
rect 309376 297956 309382 297968
rect 310054 297956 310060 297968
rect 309376 297928 310060 297956
rect 309376 297916 309382 297928
rect 310054 297916 310060 297928
rect 310112 297956 310118 297968
rect 310112 297928 316034 297956
rect 310112 297916 310118 297928
rect 316006 297888 316034 297928
rect 319346 297916 319352 297968
rect 319404 297956 319410 297968
rect 319622 297956 319628 297968
rect 319404 297928 319628 297956
rect 319404 297916 319410 297928
rect 319622 297916 319628 297928
rect 319680 297956 319686 297968
rect 382642 297956 382648 297968
rect 319680 297928 382648 297956
rect 319680 297916 319686 297928
rect 382642 297916 382648 297928
rect 382700 297916 382706 297968
rect 373166 297888 373172 297900
rect 316006 297860 373172 297888
rect 373166 297848 373172 297860
rect 373224 297848 373230 297900
rect 308674 297780 308680 297832
rect 308732 297820 308738 297832
rect 369302 297820 369308 297832
rect 308732 297792 369308 297820
rect 308732 297780 308738 297792
rect 369302 297780 369308 297792
rect 369360 297780 369366 297832
rect 307570 297712 307576 297764
rect 307628 297752 307634 297764
rect 367462 297752 367468 297764
rect 307628 297724 367468 297752
rect 307628 297712 307634 297724
rect 367462 297712 367468 297724
rect 367520 297712 367526 297764
rect 289538 297644 289544 297696
rect 289596 297684 289602 297696
rect 306282 297684 306288 297696
rect 289596 297656 306288 297684
rect 289596 297644 289602 297656
rect 306282 297644 306288 297656
rect 306340 297684 306346 297696
rect 364978 297684 364984 297696
rect 306340 297656 364984 297684
rect 306340 297644 306346 297656
rect 364978 297644 364984 297656
rect 365036 297644 365042 297696
rect 263502 297576 263508 297628
rect 263560 297616 263566 297628
rect 264054 297616 264060 297628
rect 263560 297588 264060 297616
rect 263560 297576 263566 297588
rect 264054 297576 264060 297588
rect 264112 297576 264118 297628
rect 303522 297576 303528 297628
rect 303580 297616 303586 297628
rect 363414 297616 363420 297628
rect 303580 297588 363420 297616
rect 303580 297576 303586 297588
rect 363414 297576 363420 297588
rect 363472 297576 363478 297628
rect 283834 297508 283840 297560
rect 283892 297548 283898 297560
rect 337378 297548 337384 297560
rect 283892 297520 337384 297548
rect 283892 297508 283898 297520
rect 337378 297508 337384 297520
rect 337436 297508 337442 297560
rect 230474 297440 230480 297492
rect 230532 297480 230538 297492
rect 242250 297480 242256 297492
rect 230532 297452 242256 297480
rect 230532 297440 230538 297452
rect 242250 297440 242256 297452
rect 242308 297440 242314 297492
rect 292298 297440 292304 297492
rect 292356 297480 292362 297492
rect 342990 297480 342996 297492
rect 292356 297452 342996 297480
rect 292356 297440 292362 297452
rect 342990 297440 342996 297452
rect 343048 297440 343054 297492
rect 203058 297372 203064 297424
rect 203116 297412 203122 297424
rect 263502 297412 263508 297424
rect 203116 297384 263508 297412
rect 203116 297372 203122 297384
rect 263502 297372 263508 297384
rect 263560 297372 263566 297424
rect 271690 297372 271696 297424
rect 271748 297412 271754 297424
rect 315666 297412 315672 297424
rect 271748 297384 315672 297412
rect 271748 297372 271754 297384
rect 315666 297372 315672 297384
rect 315724 297412 315730 297424
rect 335078 297412 335084 297424
rect 315724 297384 335084 297412
rect 315724 297372 315730 297384
rect 335078 297372 335084 297384
rect 335136 297372 335142 297424
rect 307938 297304 307944 297356
rect 307996 297344 308002 297356
rect 348510 297344 348516 297356
rect 307996 297316 348516 297344
rect 307996 297304 308002 297316
rect 348510 297304 348516 297316
rect 348568 297304 348574 297356
rect 178678 297236 178684 297288
rect 178736 297276 178742 297288
rect 234062 297276 234068 297288
rect 178736 297248 234068 297276
rect 178736 297236 178742 297248
rect 234062 297236 234068 297248
rect 234120 297236 234126 297288
rect 187694 297168 187700 297220
rect 187752 297208 187758 297220
rect 245010 297208 245016 297220
rect 187752 297180 245016 297208
rect 187752 297168 187758 297180
rect 245010 297168 245016 297180
rect 245068 297168 245074 297220
rect 202966 297100 202972 297152
rect 203024 297140 203030 297152
rect 262858 297140 262864 297152
rect 203024 297112 262864 297140
rect 203024 297100 203030 297112
rect 262858 297100 262864 297112
rect 262916 297100 262922 297152
rect 176654 297032 176660 297084
rect 176712 297072 176718 297084
rect 236638 297072 236644 297084
rect 176712 297044 236644 297072
rect 176712 297032 176718 297044
rect 236638 297032 236644 297044
rect 236696 297032 236702 297084
rect 293310 297032 293316 297084
rect 293368 297072 293374 297084
rect 293770 297072 293776 297084
rect 293368 297044 293776 297072
rect 293368 297032 293374 297044
rect 293770 297032 293776 297044
rect 293828 297032 293834 297084
rect 195974 296964 195980 297016
rect 196032 297004 196038 297016
rect 256878 297004 256884 297016
rect 196032 296976 256884 297004
rect 196032 296964 196038 296976
rect 256878 296964 256884 296976
rect 256936 296964 256942 297016
rect 173894 296896 173900 296948
rect 173952 296936 173958 296948
rect 235350 296936 235356 296948
rect 173952 296908 235356 296936
rect 173952 296896 173958 296908
rect 235350 296896 235356 296908
rect 235408 296896 235414 296948
rect 189074 296828 189080 296880
rect 189132 296868 189138 296880
rect 250070 296868 250076 296880
rect 189132 296840 250076 296868
rect 189132 296828 189138 296840
rect 250070 296828 250076 296840
rect 250128 296828 250134 296880
rect 183554 296760 183560 296812
rect 183612 296800 183618 296812
rect 244550 296800 244556 296812
rect 183612 296772 244556 296800
rect 183612 296760 183618 296772
rect 244550 296760 244556 296772
rect 244608 296760 244614 296812
rect 203978 296692 203984 296744
rect 204036 296732 204042 296744
rect 288618 296732 288624 296744
rect 204036 296704 288624 296732
rect 204036 296692 204042 296704
rect 288618 296692 288624 296704
rect 288676 296692 288682 296744
rect 305914 296692 305920 296744
rect 305972 296732 305978 296744
rect 306926 296732 306932 296744
rect 305972 296704 306932 296732
rect 305972 296692 305978 296704
rect 306926 296692 306932 296704
rect 306984 296692 306990 296744
rect 287974 296624 287980 296676
rect 288032 296664 288038 296676
rect 346946 296664 346952 296676
rect 288032 296636 346952 296664
rect 288032 296624 288038 296636
rect 346946 296624 346952 296636
rect 347004 296624 347010 296676
rect 236822 296080 236828 296132
rect 236880 296120 236886 296132
rect 245102 296120 245108 296132
rect 236880 296092 245108 296120
rect 236880 296080 236886 296092
rect 245102 296080 245108 296092
rect 245160 296080 245166 296132
rect 169754 296012 169760 296064
rect 169812 296052 169818 296064
rect 230474 296052 230480 296064
rect 169812 296024 230480 296052
rect 169812 296012 169818 296024
rect 230474 296012 230480 296024
rect 230532 296012 230538 296064
rect 240134 296052 240140 296064
rect 238726 296024 240140 296052
rect 210510 295944 210516 295996
rect 210568 295984 210574 295996
rect 235166 295984 235172 295996
rect 210568 295956 235172 295984
rect 210568 295944 210574 295956
rect 235166 295944 235172 295956
rect 235224 295944 235230 295996
rect 212902 295876 212908 295928
rect 212960 295916 212966 295928
rect 238726 295916 238754 296024
rect 240134 296012 240140 296024
rect 240192 296052 240198 296064
rect 264514 296052 264520 296064
rect 240192 296024 264520 296052
rect 240192 296012 240198 296024
rect 264514 296012 264520 296024
rect 264572 296012 264578 296064
rect 272334 295984 272340 295996
rect 212960 295888 238754 295916
rect 248386 295956 272340 295984
rect 212960 295876 212966 295888
rect 213178 295808 213184 295860
rect 213236 295848 213242 295860
rect 243078 295848 243084 295860
rect 213236 295820 243084 295848
rect 213236 295808 213242 295820
rect 243078 295808 243084 295820
rect 243136 295848 243142 295860
rect 248386 295848 248414 295956
rect 272334 295944 272340 295956
rect 272392 295944 272398 295996
rect 243136 295820 248414 295848
rect 243136 295808 243142 295820
rect 212994 295740 213000 295792
rect 213052 295780 213058 295792
rect 248598 295780 248604 295792
rect 213052 295752 248604 295780
rect 213052 295740 213058 295752
rect 248598 295740 248604 295752
rect 248656 295780 248662 295792
rect 249150 295780 249156 295792
rect 248656 295752 249156 295780
rect 248656 295740 248662 295752
rect 249150 295740 249156 295752
rect 249208 295740 249214 295792
rect 176746 295672 176752 295724
rect 176804 295712 176810 295724
rect 236822 295712 236828 295724
rect 176804 295684 236828 295712
rect 176804 295672 176810 295684
rect 236822 295672 236828 295684
rect 236880 295672 236886 295724
rect 173986 295604 173992 295656
rect 174044 295644 174050 295656
rect 233878 295644 233884 295656
rect 174044 295616 233884 295644
rect 174044 295604 174050 295616
rect 233878 295604 233884 295616
rect 233936 295604 233942 295656
rect 171134 295536 171140 295588
rect 171192 295576 171198 295588
rect 232406 295576 232412 295588
rect 171192 295548 232412 295576
rect 171192 295536 171198 295548
rect 232406 295536 232412 295548
rect 232464 295536 232470 295588
rect 172514 295468 172520 295520
rect 172572 295508 172578 295520
rect 233970 295508 233976 295520
rect 172572 295480 233976 295508
rect 172572 295468 172578 295480
rect 233970 295468 233976 295480
rect 234028 295468 234034 295520
rect 190454 295400 190460 295452
rect 190512 295440 190518 295452
rect 251174 295440 251180 295452
rect 190512 295412 251180 295440
rect 190512 295400 190518 295412
rect 251174 295400 251180 295412
rect 251232 295400 251238 295452
rect 297726 295400 297732 295452
rect 297784 295440 297790 295452
rect 305546 295440 305552 295452
rect 297784 295412 305552 295440
rect 297784 295400 297790 295412
rect 305546 295400 305552 295412
rect 305604 295400 305610 295452
rect 230934 295332 230940 295384
rect 230992 295372 230998 295384
rect 231670 295372 231676 295384
rect 230992 295344 231676 295372
rect 230992 295332 230998 295344
rect 231670 295332 231676 295344
rect 231728 295372 231734 295384
rect 231728 295344 233832 295372
rect 231728 295332 231734 295344
rect 233804 295304 233832 295344
rect 233878 295332 233884 295384
rect 233936 295372 233942 295384
rect 234522 295372 234528 295384
rect 233936 295344 234528 295372
rect 233936 295332 233942 295344
rect 234522 295332 234528 295344
rect 234580 295332 234586 295384
rect 577590 295372 577596 295384
rect 234632 295344 577596 295372
rect 234632 295304 234660 295344
rect 577590 295332 577596 295344
rect 577648 295332 577654 295384
rect 233804 295276 234660 295304
rect 288894 295264 288900 295316
rect 288952 295304 288958 295316
rect 347038 295304 347044 295316
rect 288952 295276 347044 295304
rect 288952 295264 288958 295276
rect 347038 295264 347044 295276
rect 347096 295264 347102 295316
rect 288618 295196 288624 295248
rect 288676 295236 288682 295248
rect 342898 295236 342904 295248
rect 288676 295208 342904 295236
rect 288676 295196 288682 295208
rect 342898 295196 342904 295208
rect 342956 295196 342962 295248
rect 287606 295128 287612 295180
rect 287664 295168 287670 295180
rect 340138 295168 340144 295180
rect 287664 295140 340144 295168
rect 287664 295128 287670 295140
rect 340138 295128 340144 295140
rect 340196 295128 340202 295180
rect 291654 295060 291660 295112
rect 291712 295100 291718 295112
rect 344278 295100 344284 295112
rect 291712 295072 344284 295100
rect 291712 295060 291718 295072
rect 344278 295060 344284 295072
rect 344336 295060 344342 295112
rect 166994 294788 167000 294840
rect 167052 294828 167058 294840
rect 228266 294828 228272 294840
rect 167052 294800 228272 294828
rect 167052 294788 167058 294800
rect 228266 294788 228272 294800
rect 228324 294788 228330 294840
rect 242802 294788 242808 294840
rect 242860 294828 242866 294840
rect 272426 294828 272432 294840
rect 242860 294800 272432 294828
rect 242860 294788 242866 294800
rect 272426 294788 272432 294800
rect 272484 294788 272490 294840
rect 168374 294720 168380 294772
rect 168432 294760 168438 294772
rect 229094 294760 229100 294772
rect 168432 294732 229100 294760
rect 168432 294720 168438 294732
rect 229094 294720 229100 294732
rect 229152 294760 229158 294772
rect 229830 294760 229836 294772
rect 229152 294732 229836 294760
rect 229152 294720 229158 294732
rect 229830 294720 229836 294732
rect 229888 294720 229894 294772
rect 235718 294720 235724 294772
rect 235776 294760 235782 294772
rect 267274 294760 267280 294772
rect 235776 294732 267280 294760
rect 235776 294720 235782 294732
rect 267274 294720 267280 294732
rect 267332 294720 267338 294772
rect 222470 294652 222476 294704
rect 222528 294692 222534 294704
rect 283006 294692 283012 294704
rect 222528 294664 283012 294692
rect 222528 294652 222534 294664
rect 283006 294652 283012 294664
rect 283064 294652 283070 294704
rect 164234 294584 164240 294636
rect 164292 294624 164298 294636
rect 224862 294624 224868 294636
rect 164292 294596 224868 294624
rect 164292 294584 164298 294596
rect 224862 294584 224868 294596
rect 224920 294584 224926 294636
rect 237466 294584 237472 294636
rect 237524 294624 237530 294636
rect 275094 294624 275100 294636
rect 237524 294596 275100 294624
rect 237524 294584 237530 294596
rect 275094 294584 275100 294596
rect 275152 294584 275158 294636
rect 213730 294516 213736 294568
rect 213788 294556 213794 294568
rect 232038 294556 232044 294568
rect 213788 294528 232044 294556
rect 213788 294516 213794 294528
rect 232038 294516 232044 294528
rect 232096 294556 232102 294568
rect 233142 294556 233148 294568
rect 232096 294528 233148 294556
rect 232096 294516 232102 294528
rect 233142 294516 233148 294528
rect 233200 294516 233206 294568
rect 171226 294448 171232 294500
rect 171284 294488 171290 294500
rect 231118 294488 231124 294500
rect 171284 294460 231124 294488
rect 171284 294448 171290 294460
rect 231118 294448 231124 294460
rect 231176 294448 231182 294500
rect 165890 294380 165896 294432
rect 165948 294420 165954 294432
rect 225598 294420 225604 294432
rect 165948 294392 225604 294420
rect 165948 294380 165954 294392
rect 225598 294380 225604 294392
rect 225656 294380 225662 294432
rect 169846 294312 169852 294364
rect 169904 294352 169910 294364
rect 229922 294352 229928 294364
rect 169904 294324 229928 294352
rect 169904 294312 169910 294324
rect 229922 294312 229928 294324
rect 229980 294352 229986 294364
rect 230198 294352 230204 294364
rect 229980 294324 230204 294352
rect 229980 294312 229986 294324
rect 230198 294312 230204 294324
rect 230256 294312 230262 294364
rect 287606 294312 287612 294364
rect 287664 294352 287670 294364
rect 288250 294352 288256 294364
rect 287664 294324 288256 294352
rect 287664 294312 287670 294324
rect 288250 294312 288256 294324
rect 288308 294312 288314 294364
rect 182174 294244 182180 294296
rect 182232 294284 182238 294296
rect 242710 294284 242716 294296
rect 182232 294256 242716 294284
rect 182232 294244 182238 294256
rect 242710 294244 242716 294256
rect 242768 294244 242774 294296
rect 176838 294176 176844 294228
rect 176896 294216 176902 294228
rect 237926 294216 237932 294228
rect 176896 294188 237932 294216
rect 176896 294176 176902 294188
rect 237926 294176 237932 294188
rect 237984 294176 237990 294228
rect 165706 294108 165712 294160
rect 165764 294148 165770 294160
rect 226886 294148 226892 294160
rect 165764 294120 226892 294148
rect 165764 294108 165770 294120
rect 226886 294108 226892 294120
rect 226944 294108 226950 294160
rect 225598 294040 225604 294092
rect 225656 294080 225662 294092
rect 225782 294080 225788 294092
rect 225656 294052 225788 294080
rect 225656 294040 225662 294052
rect 225782 294040 225788 294052
rect 225840 294040 225846 294092
rect 216490 293972 216496 294024
rect 216548 294012 216554 294024
rect 241974 294012 241980 294024
rect 216548 293984 241980 294012
rect 216548 293972 216554 293984
rect 241974 293972 241980 293984
rect 242032 294012 242038 294024
rect 242802 294012 242808 294024
rect 242032 293984 242808 294012
rect 242032 293972 242038 293984
rect 242802 293972 242808 293984
rect 242860 293972 242866 294024
rect 226334 293904 226340 293956
rect 226392 293944 226398 293956
rect 229738 293944 229744 293956
rect 226392 293916 229744 293944
rect 226392 293904 226398 293916
rect 229738 293904 229744 293916
rect 229796 293904 229802 293956
rect 198734 293428 198740 293480
rect 198792 293468 198798 293480
rect 253106 293468 253112 293480
rect 198792 293440 253112 293468
rect 198792 293428 198798 293440
rect 253106 293428 253112 293440
rect 253164 293428 253170 293480
rect 237374 293360 237380 293412
rect 237432 293400 237438 293412
rect 275186 293400 275192 293412
rect 237432 293372 275192 293400
rect 237432 293360 237438 293372
rect 275186 293360 275192 293372
rect 275244 293360 275250 293412
rect 164878 293292 164884 293344
rect 164936 293332 164942 293344
rect 225690 293332 225696 293344
rect 164936 293304 225696 293332
rect 164936 293292 164942 293304
rect 225690 293292 225696 293304
rect 225748 293292 225754 293344
rect 236086 293292 236092 293344
rect 236144 293332 236150 293344
rect 278222 293332 278228 293344
rect 236144 293304 278228 293332
rect 236144 293292 236150 293304
rect 278222 293292 278228 293304
rect 278280 293292 278286 293344
rect 157794 293224 157800 293276
rect 157852 293264 157858 293276
rect 226334 293264 226340 293276
rect 157852 293236 226340 293264
rect 157852 293224 157858 293236
rect 226334 293224 226340 293236
rect 226392 293224 226398 293276
rect 235350 293224 235356 293276
rect 235408 293264 235414 293276
rect 278130 293264 278136 293276
rect 235408 293236 278136 293264
rect 235408 293224 235414 293236
rect 278130 293224 278136 293236
rect 278188 293224 278194 293276
rect 188338 293156 188344 293208
rect 188396 293196 188402 293208
rect 237466 293196 237472 293208
rect 188396 293168 237472 293196
rect 188396 293156 188402 293168
rect 237466 293156 237472 293168
rect 237524 293196 237530 293208
rect 238478 293196 238484 293208
rect 237524 293168 238484 293196
rect 237524 293156 237530 293168
rect 238478 293156 238484 293168
rect 238536 293156 238542 293208
rect 172698 293088 172704 293140
rect 172756 293128 172762 293140
rect 233142 293128 233148 293140
rect 172756 293100 233148 293128
rect 172756 293088 172762 293100
rect 233142 293088 233148 293100
rect 233200 293088 233206 293140
rect 164326 293020 164332 293072
rect 164384 293060 164390 293072
rect 224218 293060 224224 293072
rect 164384 293032 224224 293060
rect 164384 293020 164390 293032
rect 224218 293020 224224 293032
rect 224276 293060 224282 293072
rect 224678 293060 224684 293072
rect 224276 293032 224684 293060
rect 224276 293020 224282 293032
rect 224678 293020 224684 293032
rect 224736 293020 224742 293072
rect 254026 293020 254032 293072
rect 254084 293060 254090 293072
rect 254302 293060 254308 293072
rect 254084 293032 254308 293060
rect 254084 293020 254090 293032
rect 254302 293020 254308 293032
rect 254360 293020 254366 293072
rect 259546 293020 259552 293072
rect 259604 293060 259610 293072
rect 260190 293060 260196 293072
rect 259604 293032 260196 293060
rect 259604 293020 259610 293032
rect 260190 293020 260196 293032
rect 260248 293020 260254 293072
rect 262490 293020 262496 293072
rect 262548 293060 262554 293072
rect 263134 293060 263140 293072
rect 262548 293032 263140 293060
rect 262548 293020 262554 293032
rect 263134 293020 263140 293032
rect 263192 293020 263198 293072
rect 263686 293020 263692 293072
rect 263744 293060 263750 293072
rect 264238 293060 264244 293072
rect 263744 293032 264244 293060
rect 263744 293020 263750 293032
rect 264238 293020 264244 293032
rect 264296 293020 264302 293072
rect 179414 292952 179420 293004
rect 179472 292992 179478 293004
rect 239766 292992 239772 293004
rect 179472 292964 239772 292992
rect 179472 292952 179478 292964
rect 239766 292952 239772 292964
rect 239824 292952 239830 293004
rect 263870 292952 263876 293004
rect 263928 292992 263934 293004
rect 264606 292992 264612 293004
rect 263928 292964 264612 292992
rect 263928 292952 263934 292964
rect 264606 292952 264612 292964
rect 264664 292952 264670 293004
rect 176930 292884 176936 292936
rect 176988 292924 176994 292936
rect 237374 292924 237380 292936
rect 176988 292896 237380 292924
rect 176988 292884 176994 292896
rect 237374 292884 237380 292896
rect 237432 292884 237438 292936
rect 172606 292816 172612 292868
rect 172664 292856 172670 292868
rect 232774 292856 232780 292868
rect 172664 292828 232780 292856
rect 172664 292816 172670 292828
rect 232774 292816 232780 292828
rect 232832 292816 232838 292868
rect 175274 292748 175280 292800
rect 175332 292788 175338 292800
rect 236086 292788 236092 292800
rect 175332 292760 236092 292788
rect 175332 292748 175338 292760
rect 236086 292748 236092 292760
rect 236144 292788 236150 292800
rect 236454 292788 236460 292800
rect 236144 292760 236460 292788
rect 236144 292748 236150 292760
rect 236454 292748 236460 292760
rect 236512 292748 236518 292800
rect 216582 292680 216588 292732
rect 216640 292720 216646 292732
rect 235350 292720 235356 292732
rect 216640 292692 235356 292720
rect 216640 292680 216646 292692
rect 235350 292680 235356 292692
rect 235408 292680 235414 292732
rect 210694 292612 210700 292664
rect 210752 292652 210758 292664
rect 210752 292624 241468 292652
rect 210752 292612 210758 292624
rect 3418 292544 3424 292596
rect 3476 292584 3482 292596
rect 198734 292584 198740 292596
rect 3476 292556 198740 292584
rect 3476 292544 3482 292556
rect 198734 292544 198740 292556
rect 198792 292544 198798 292596
rect 219250 292544 219256 292596
rect 219308 292584 219314 292596
rect 228726 292584 228732 292596
rect 219308 292556 228732 292584
rect 219308 292544 219314 292556
rect 228726 292544 228732 292556
rect 228784 292544 228790 292596
rect 235166 292476 235172 292528
rect 235224 292516 235230 292528
rect 236086 292516 236092 292528
rect 235224 292488 236092 292516
rect 235224 292476 235230 292488
rect 236086 292476 236092 292488
rect 236144 292476 236150 292528
rect 237466 292476 237472 292528
rect 237524 292516 237530 292528
rect 238570 292516 238576 292528
rect 237524 292488 238576 292516
rect 237524 292476 237530 292488
rect 238570 292476 238576 292488
rect 238628 292516 238634 292528
rect 239398 292516 239404 292528
rect 238628 292488 239404 292516
rect 238628 292476 238634 292488
rect 239398 292476 239404 292488
rect 239456 292476 239462 292528
rect 241440 292516 241468 292624
rect 242250 292516 242256 292528
rect 241440 292488 242256 292516
rect 242250 292476 242256 292488
rect 242308 292476 242314 292528
rect 261478 292476 261484 292528
rect 261536 292516 261542 292528
rect 262214 292516 262220 292528
rect 261536 292488 262220 292516
rect 261536 292476 261542 292488
rect 262214 292476 262220 292488
rect 262272 292476 262278 292528
rect 264422 292476 264428 292528
rect 264480 292516 264486 292528
rect 264974 292516 264980 292528
rect 264480 292488 264980 292516
rect 264480 292476 264486 292488
rect 264974 292476 264980 292488
rect 265032 292476 265038 292528
rect 311618 292476 311624 292528
rect 311676 292516 311682 292528
rect 376754 292516 376760 292528
rect 311676 292488 376760 292516
rect 311676 292476 311682 292488
rect 376754 292476 376760 292488
rect 376812 292516 376818 292528
rect 378134 292516 378140 292528
rect 376812 292488 378140 292516
rect 376812 292476 376818 292488
rect 378134 292476 378140 292488
rect 378192 292476 378198 292528
rect 240870 292408 240876 292460
rect 240928 292448 240934 292460
rect 275738 292448 275744 292460
rect 240928 292420 275744 292448
rect 240928 292408 240934 292420
rect 275738 292408 275744 292420
rect 275796 292408 275802 292460
rect 218882 292340 218888 292392
rect 218940 292380 218946 292392
rect 255958 292380 255964 292392
rect 218940 292352 255964 292380
rect 218940 292340 218946 292352
rect 255958 292340 255964 292352
rect 256016 292340 256022 292392
rect 246666 292272 246672 292324
rect 246724 292312 246730 292324
rect 267182 292312 267188 292324
rect 246724 292284 267188 292312
rect 246724 292272 246730 292284
rect 267182 292272 267188 292284
rect 267240 292272 267246 292324
rect 240502 292204 240508 292256
rect 240560 292244 240566 292256
rect 264514 292244 264520 292256
rect 240560 292216 264520 292244
rect 240560 292204 240566 292216
rect 264514 292204 264520 292216
rect 264572 292204 264578 292256
rect 245286 292136 245292 292188
rect 245344 292176 245350 292188
rect 269758 292176 269764 292188
rect 245344 292148 269764 292176
rect 245344 292136 245350 292148
rect 269758 292136 269764 292148
rect 269816 292136 269822 292188
rect 221458 292068 221464 292120
rect 221516 292108 221522 292120
rect 237374 292108 237380 292120
rect 221516 292080 237380 292108
rect 221516 292068 221522 292080
rect 237374 292068 237380 292080
rect 237432 292068 237438 292120
rect 252830 292068 252836 292120
rect 252888 292108 252894 292120
rect 279694 292108 279700 292120
rect 252888 292080 279700 292108
rect 252888 292068 252894 292080
rect 279694 292068 279700 292080
rect 279752 292068 279758 292120
rect 307110 292068 307116 292120
rect 307168 292108 307174 292120
rect 311618 292108 311624 292120
rect 307168 292080 311624 292108
rect 307168 292068 307174 292080
rect 311618 292068 311624 292080
rect 311676 292068 311682 292120
rect 220814 292000 220820 292052
rect 220872 292040 220878 292052
rect 237466 292040 237472 292052
rect 220872 292012 237472 292040
rect 220872 292000 220878 292012
rect 237466 292000 237472 292012
rect 237524 292000 237530 292052
rect 244182 292000 244188 292052
rect 244240 292040 244246 292052
rect 273070 292040 273076 292052
rect 244240 292012 273076 292040
rect 244240 292000 244246 292012
rect 273070 292000 273076 292012
rect 273128 292000 273134 292052
rect 218606 291932 218612 291984
rect 218664 291972 218670 291984
rect 220170 291972 220176 291984
rect 218664 291944 220176 291972
rect 218664 291932 218670 291944
rect 220170 291932 220176 291944
rect 220228 291972 220234 291984
rect 254854 291972 254860 291984
rect 220228 291944 254860 291972
rect 220228 291932 220234 291944
rect 254854 291932 254860 291944
rect 254912 291932 254918 291984
rect 218514 291864 218520 291916
rect 218572 291904 218578 291916
rect 222102 291904 222108 291916
rect 218572 291876 222108 291904
rect 218572 291864 218578 291876
rect 222102 291864 222108 291876
rect 222160 291904 222166 291916
rect 224402 291904 224408 291916
rect 222160 291876 224408 291904
rect 222160 291864 222166 291876
rect 224402 291864 224408 291876
rect 224460 291864 224466 291916
rect 237374 291864 237380 291916
rect 237432 291904 237438 291916
rect 238294 291904 238300 291916
rect 237432 291876 238300 291904
rect 237432 291864 237438 291876
rect 238294 291864 238300 291876
rect 238352 291904 238358 291916
rect 275646 291904 275652 291916
rect 238352 291876 275652 291904
rect 238352 291864 238358 291876
rect 275646 291864 275652 291876
rect 275704 291864 275710 291916
rect 215938 291796 215944 291848
rect 215996 291836 216002 291848
rect 221734 291836 221740 291848
rect 215996 291808 221740 291836
rect 215996 291796 216002 291808
rect 221734 291796 221740 291808
rect 221792 291796 221798 291848
rect 258166 291796 258172 291848
rect 258224 291836 258230 291848
rect 271046 291836 271052 291848
rect 258224 291808 271052 291836
rect 258224 291796 258230 291808
rect 271046 291796 271052 291808
rect 271104 291836 271110 291848
rect 272150 291836 272156 291848
rect 271104 291808 272156 291836
rect 271104 291796 271110 291808
rect 272150 291796 272156 291808
rect 272208 291796 272214 291848
rect 272334 291796 272340 291848
rect 272392 291836 272398 291848
rect 334158 291836 334164 291848
rect 272392 291808 334164 291836
rect 272392 291796 272398 291808
rect 334158 291796 334164 291808
rect 334216 291796 334222 291848
rect 219894 291728 219900 291780
rect 219952 291768 219958 291780
rect 249058 291768 249064 291780
rect 219952 291740 249064 291768
rect 219952 291728 219958 291740
rect 249058 291728 249064 291740
rect 249116 291728 249122 291780
rect 251910 291728 251916 291780
rect 251968 291768 251974 291780
rect 264146 291768 264152 291780
rect 251968 291740 264152 291768
rect 251968 291728 251974 291740
rect 264146 291728 264152 291740
rect 264204 291728 264210 291780
rect 217226 291660 217232 291712
rect 217284 291700 217290 291712
rect 229462 291700 229468 291712
rect 217284 291672 229468 291700
rect 217284 291660 217290 291672
rect 229462 291660 229468 291672
rect 229520 291700 229526 291712
rect 230014 291700 230020 291712
rect 229520 291672 230020 291700
rect 229520 291660 229526 291672
rect 230014 291660 230020 291672
rect 230072 291660 230078 291712
rect 232774 291660 232780 291712
rect 232832 291700 232838 291712
rect 275370 291700 275376 291712
rect 232832 291672 275376 291700
rect 232832 291660 232838 291672
rect 275370 291660 275376 291672
rect 275428 291660 275434 291712
rect 221274 291592 221280 291644
rect 221332 291632 221338 291644
rect 241882 291632 241888 291644
rect 221332 291604 241888 291632
rect 221332 291592 221338 291604
rect 241882 291592 241888 291604
rect 241940 291592 241946 291644
rect 255038 291592 255044 291644
rect 255096 291632 255102 291644
rect 272702 291632 272708 291644
rect 255096 291604 272708 291632
rect 255096 291592 255102 291604
rect 272702 291592 272708 291604
rect 272760 291592 272766 291644
rect 221366 291524 221372 291576
rect 221424 291564 221430 291576
rect 243630 291564 243636 291576
rect 221424 291536 243636 291564
rect 221424 291524 221430 291536
rect 243630 291524 243636 291536
rect 243688 291524 243694 291576
rect 253106 291524 253112 291576
rect 253164 291564 253170 291576
rect 258718 291564 258724 291576
rect 253164 291536 258724 291564
rect 253164 291524 253170 291536
rect 258718 291524 258724 291536
rect 258776 291524 258782 291576
rect 271966 291524 271972 291576
rect 272024 291564 272030 291576
rect 272610 291564 272616 291576
rect 272024 291536 272616 291564
rect 272024 291524 272030 291536
rect 272610 291524 272616 291536
rect 272668 291524 272674 291576
rect 220078 291456 220084 291508
rect 220136 291496 220142 291508
rect 244918 291496 244924 291508
rect 220136 291468 244924 291496
rect 220136 291456 220142 291468
rect 244918 291456 244924 291468
rect 244976 291456 244982 291508
rect 256694 291456 256700 291508
rect 256752 291496 256758 291508
rect 259270 291496 259276 291508
rect 256752 291468 259276 291496
rect 256752 291456 256758 291468
rect 259270 291456 259276 291468
rect 259328 291456 259334 291508
rect 220906 291388 220912 291440
rect 220964 291428 220970 291440
rect 246390 291428 246396 291440
rect 220964 291400 246396 291428
rect 220964 291388 220970 291400
rect 246390 291388 246396 291400
rect 246448 291388 246454 291440
rect 263686 291388 263692 291440
rect 263744 291428 263750 291440
rect 272058 291428 272064 291440
rect 263744 291400 272064 291428
rect 263744 291388 263750 291400
rect 272058 291388 272064 291400
rect 272116 291428 272122 291440
rect 272334 291428 272340 291440
rect 272116 291400 272340 291428
rect 272116 291388 272122 291400
rect 272334 291388 272340 291400
rect 272392 291388 272398 291440
rect 219802 291320 219808 291372
rect 219860 291360 219866 291372
rect 247402 291360 247408 291372
rect 219860 291332 247408 291360
rect 219860 291320 219866 291332
rect 247402 291320 247408 291332
rect 247460 291320 247466 291372
rect 262582 291320 262588 291372
rect 262640 291360 262646 291372
rect 270494 291360 270500 291372
rect 262640 291332 270500 291360
rect 262640 291320 262646 291332
rect 270494 291320 270500 291332
rect 270552 291360 270558 291372
rect 271230 291360 271236 291372
rect 270552 291332 271236 291360
rect 270552 291320 270558 291332
rect 271230 291320 271236 291332
rect 271288 291320 271294 291372
rect 217318 291252 217324 291304
rect 217376 291292 217382 291304
rect 227162 291292 227168 291304
rect 217376 291264 227168 291292
rect 217376 291252 217382 291264
rect 227162 291252 227168 291264
rect 227220 291252 227226 291304
rect 227714 291252 227720 291304
rect 227772 291292 227778 291304
rect 234246 291292 234252 291304
rect 227772 291264 234252 291292
rect 227772 291252 227778 291264
rect 234246 291252 234252 291264
rect 234304 291252 234310 291304
rect 244274 291252 244280 291304
rect 244332 291292 244338 291304
rect 246298 291292 246304 291304
rect 244332 291264 246304 291292
rect 244332 291252 244338 291264
rect 246298 291252 246304 291264
rect 246356 291292 246362 291304
rect 246758 291292 246764 291304
rect 246356 291264 246764 291292
rect 246356 291252 246362 291264
rect 246758 291252 246764 291264
rect 246816 291252 246822 291304
rect 246942 291252 246948 291304
rect 247000 291292 247006 291304
rect 249702 291292 249708 291304
rect 247000 291264 249708 291292
rect 247000 291252 247006 291264
rect 249702 291252 249708 291264
rect 249760 291252 249766 291304
rect 256142 291252 256148 291304
rect 256200 291292 256206 291304
rect 257798 291292 257804 291304
rect 256200 291264 257804 291292
rect 256200 291252 256206 291264
rect 257798 291252 257804 291264
rect 257856 291252 257862 291304
rect 261110 291252 261116 291304
rect 261168 291292 261174 291304
rect 270770 291292 270776 291304
rect 261168 291264 270776 291292
rect 261168 291252 261174 291264
rect 270770 291252 270776 291264
rect 270828 291292 270834 291304
rect 271138 291292 271144 291304
rect 270828 291264 271144 291292
rect 270828 291252 270834 291264
rect 271138 291252 271144 291264
rect 271196 291252 271202 291304
rect 227806 291184 227812 291236
rect 227864 291224 227870 291236
rect 229830 291224 229836 291236
rect 227864 291196 229836 291224
rect 227864 291184 227870 291196
rect 229830 291184 229836 291196
rect 229888 291184 229894 291236
rect 245010 291184 245016 291236
rect 245068 291224 245074 291236
rect 247862 291224 247868 291236
rect 245068 291196 247868 291224
rect 245068 291184 245074 291196
rect 247862 291184 247868 291196
rect 247920 291184 247926 291236
rect 259362 291184 259368 291236
rect 259420 291224 259426 291236
rect 260742 291224 260748 291236
rect 259420 291196 260748 291224
rect 259420 291184 259426 291196
rect 260742 291184 260748 291196
rect 260800 291184 260806 291236
rect 261478 291184 261484 291236
rect 261536 291224 261542 291236
rect 271966 291224 271972 291236
rect 261536 291196 271972 291224
rect 261536 291184 261542 291196
rect 271966 291184 271972 291196
rect 272024 291184 272030 291236
rect 239766 291116 239772 291168
rect 239824 291156 239830 291168
rect 279050 291156 279056 291168
rect 239824 291128 279056 291156
rect 239824 291116 239830 291128
rect 279050 291116 279056 291128
rect 279108 291116 279114 291168
rect 325694 291116 325700 291168
rect 325752 291156 325758 291168
rect 327534 291156 327540 291168
rect 325752 291128 327540 291156
rect 325752 291116 325758 291128
rect 327534 291116 327540 291128
rect 327592 291116 327598 291168
rect 233142 291048 233148 291100
rect 233200 291088 233206 291100
rect 268378 291088 268384 291100
rect 233200 291060 268384 291088
rect 233200 291048 233206 291060
rect 268378 291048 268384 291060
rect 268436 291048 268442 291100
rect 169938 290776 169944 290828
rect 169996 290816 170002 290828
rect 230934 290816 230940 290828
rect 169996 290788 230940 290816
rect 169996 290776 170002 290788
rect 230934 290776 230940 290788
rect 230992 290776 230998 290828
rect 173802 290708 173808 290760
rect 173860 290748 173866 290760
rect 220630 290748 220636 290760
rect 173860 290720 220636 290748
rect 173860 290708 173866 290720
rect 220630 290708 220636 290720
rect 220688 290748 220694 290760
rect 227806 290748 227812 290760
rect 220688 290720 227812 290748
rect 220688 290708 220694 290720
rect 227806 290708 227812 290720
rect 227864 290708 227870 290760
rect 168282 290640 168288 290692
rect 168340 290680 168346 290692
rect 220722 290680 220728 290692
rect 168340 290652 220728 290680
rect 168340 290640 168346 290652
rect 220722 290640 220728 290652
rect 220780 290640 220786 290692
rect 243446 290640 243452 290692
rect 243504 290680 243510 290692
rect 277210 290680 277216 290692
rect 243504 290652 277216 290680
rect 243504 290640 243510 290652
rect 277210 290640 277216 290652
rect 277268 290640 277274 290692
rect 200758 290572 200764 290624
rect 200816 290612 200822 290624
rect 259362 290612 259368 290624
rect 200816 290584 259368 290612
rect 200816 290572 200822 290584
rect 259362 290572 259368 290584
rect 259420 290572 259426 290624
rect 194686 290504 194692 290556
rect 194744 290544 194750 290556
rect 255038 290544 255044 290556
rect 194744 290516 255044 290544
rect 194744 290504 194750 290516
rect 255038 290504 255044 290516
rect 255096 290504 255102 290556
rect 191926 290436 191932 290488
rect 191984 290476 191990 290488
rect 252830 290476 252836 290488
rect 191984 290448 252836 290476
rect 191984 290436 191990 290448
rect 252830 290436 252836 290448
rect 252888 290436 252894 290488
rect 327534 290436 327540 290488
rect 327592 290476 327598 290488
rect 394694 290476 394700 290488
rect 327592 290448 394700 290476
rect 327592 290436 327598 290448
rect 394694 290436 394700 290448
rect 394752 290476 394758 290488
rect 569954 290476 569960 290488
rect 394752 290448 569960 290476
rect 394752 290436 394758 290448
rect 569954 290436 569960 290448
rect 570012 290436 570018 290488
rect 182266 290368 182272 290420
rect 182324 290408 182330 290420
rect 243446 290408 243452 290420
rect 182324 290380 243452 290408
rect 182324 290368 182330 290380
rect 243446 290368 243452 290380
rect 243504 290368 243510 290420
rect 221550 290300 221556 290352
rect 221608 290340 221614 290352
rect 254118 290340 254124 290352
rect 221608 290312 254124 290340
rect 221608 290300 221614 290312
rect 254118 290300 254124 290312
rect 254176 290300 254182 290352
rect 221642 290232 221648 290284
rect 221700 290272 221706 290284
rect 256786 290272 256792 290284
rect 221700 290244 256792 290272
rect 221700 290232 221706 290244
rect 256786 290232 256792 290244
rect 256844 290272 256850 290284
rect 257062 290272 257068 290284
rect 256844 290244 257068 290272
rect 256844 290232 256850 290244
rect 257062 290232 257068 290244
rect 257120 290232 257126 290284
rect 220354 290164 220360 290216
rect 220412 290204 220418 290216
rect 259638 290204 259644 290216
rect 220412 290176 259644 290204
rect 220412 290164 220418 290176
rect 259638 290164 259644 290176
rect 259696 290164 259702 290216
rect 197538 290096 197544 290148
rect 197596 290136 197602 290148
rect 257246 290136 257252 290148
rect 197596 290108 257252 290136
rect 197596 290096 197602 290108
rect 257246 290096 257252 290108
rect 257304 290136 257310 290148
rect 257430 290136 257436 290148
rect 257304 290108 257436 290136
rect 257304 290096 257310 290108
rect 257430 290096 257436 290108
rect 257488 290096 257494 290148
rect 196066 290028 196072 290080
rect 196124 290068 196130 290080
rect 255498 290068 255504 290080
rect 196124 290040 255504 290068
rect 196124 290028 196130 290040
rect 255498 290028 255504 290040
rect 255556 290068 255562 290080
rect 256142 290068 256148 290080
rect 255556 290040 256148 290068
rect 255556 290028 255562 290040
rect 256142 290028 256148 290040
rect 256200 290028 256206 290080
rect 201494 289960 201500 290012
rect 201552 290000 201558 290012
rect 261662 290000 261668 290012
rect 201552 289972 261668 290000
rect 201552 289960 201558 289972
rect 261662 289960 261668 289972
rect 261720 289960 261726 290012
rect 221734 289892 221740 289944
rect 221792 289932 221798 289944
rect 240410 289932 240416 289944
rect 221792 289904 240416 289932
rect 221792 289892 221798 289904
rect 240410 289892 240416 289904
rect 240468 289892 240474 289944
rect 178034 289824 178040 289876
rect 178092 289864 178098 289876
rect 238846 289864 238852 289876
rect 178092 289836 238852 289864
rect 178092 289824 178098 289836
rect 238846 289824 238852 289836
rect 238904 289824 238910 289876
rect 219710 289756 219716 289808
rect 219768 289796 219774 289808
rect 223574 289796 223580 289808
rect 219768 289768 223580 289796
rect 219768 289756 219774 289768
rect 223574 289756 223580 289768
rect 223632 289756 223638 289808
rect 244826 289756 244832 289808
rect 244884 289796 244890 289808
rect 246206 289796 246212 289808
rect 244884 289768 246212 289796
rect 244884 289756 244890 289768
rect 246206 289756 246212 289768
rect 246264 289756 246270 289808
rect 300578 289552 300584 289604
rect 300636 289592 300642 289604
rect 306190 289592 306196 289604
rect 300636 289564 306196 289592
rect 300636 289552 300642 289564
rect 306190 289552 306196 289564
rect 306248 289552 306254 289604
rect 242618 289416 242624 289468
rect 242676 289456 242682 289468
rect 242676 289428 253934 289456
rect 242676 289416 242682 289428
rect 235534 289388 235540 289400
rect 219406 289360 235540 289388
rect 174078 289280 174084 289332
rect 174136 289320 174142 289332
rect 218054 289320 218060 289332
rect 174136 289292 218060 289320
rect 174136 289280 174142 289292
rect 218054 289280 218060 289292
rect 218112 289280 218118 289332
rect 180058 289212 180064 289264
rect 180116 289252 180122 289264
rect 219406 289252 219434 289360
rect 235534 289348 235540 289360
rect 235592 289348 235598 289400
rect 243998 289388 244004 289400
rect 238726 289360 244004 289388
rect 180116 289224 219434 289252
rect 180116 289212 180122 289224
rect 183646 289144 183652 289196
rect 183704 289184 183710 289196
rect 238726 289184 238754 289360
rect 243998 289348 244004 289360
rect 244056 289348 244062 289400
rect 245562 289388 245568 289400
rect 244108 289360 245568 289388
rect 244108 289320 244136 289360
rect 245562 289348 245568 289360
rect 245620 289348 245626 289400
rect 183704 289156 238754 289184
rect 244016 289292 244136 289320
rect 183704 289144 183710 289156
rect 184934 289076 184940 289128
rect 184992 289116 184998 289128
rect 244016 289116 244044 289292
rect 184992 289088 244044 289116
rect 184992 289076 184998 289088
rect 253906 288436 253934 289428
rect 274266 288436 274272 288448
rect 253906 288408 274272 288436
rect 274266 288396 274272 288408
rect 274324 288396 274330 288448
rect 269022 287648 269028 287700
rect 269080 287688 269086 287700
rect 319714 287688 319720 287700
rect 269080 287660 319720 287688
rect 269080 287648 269086 287660
rect 319714 287648 319720 287660
rect 319772 287648 319778 287700
rect 349246 286492 349252 286544
rect 349304 286532 349310 286544
rect 350258 286532 350264 286544
rect 349304 286504 350264 286532
rect 349304 286492 349310 286504
rect 350258 286492 350264 286504
rect 350316 286492 350322 286544
rect 169662 286288 169668 286340
rect 169720 286328 169726 286340
rect 219250 286328 219256 286340
rect 169720 286300 219256 286328
rect 169720 286288 169726 286300
rect 219250 286288 219256 286300
rect 219308 286288 219314 286340
rect 310238 286288 310244 286340
rect 310296 286328 310302 286340
rect 349246 286328 349252 286340
rect 310296 286300 349252 286328
rect 310296 286288 310302 286300
rect 349246 286288 349252 286300
rect 349304 286288 349310 286340
rect 310054 285676 310060 285728
rect 310112 285716 310118 285728
rect 310238 285716 310244 285728
rect 310112 285688 310244 285716
rect 310112 285676 310118 285688
rect 310238 285676 310244 285688
rect 310296 285676 310302 285728
rect 268930 285064 268936 285116
rect 268988 285104 268994 285116
rect 268988 285076 277394 285104
rect 268988 285064 268994 285076
rect 277366 285036 277394 285076
rect 315482 285036 315488 285048
rect 277366 285008 315488 285036
rect 315482 284996 315488 285008
rect 315540 284996 315546 285048
rect 185118 284928 185124 284980
rect 185176 284968 185182 284980
rect 220906 284968 220912 284980
rect 185176 284940 220912 284968
rect 185176 284928 185182 284940
rect 220906 284928 220912 284940
rect 220964 284928 220970 284980
rect 268930 284928 268936 284980
rect 268988 284968 268994 284980
rect 326706 284968 326712 284980
rect 268988 284940 326712 284968
rect 268988 284928 268994 284940
rect 326706 284928 326712 284940
rect 326764 284928 326770 284980
rect 180794 283568 180800 283620
rect 180852 283608 180858 283620
rect 220906 283608 220912 283620
rect 180852 283580 220912 283608
rect 180852 283568 180858 283580
rect 220906 283568 220912 283580
rect 220964 283568 220970 283620
rect 269758 283568 269764 283620
rect 269816 283608 269822 283620
rect 325234 283608 325240 283620
rect 269816 283580 325240 283608
rect 269816 283568 269822 283580
rect 325234 283568 325240 283580
rect 325292 283568 325298 283620
rect 183738 282140 183744 282192
rect 183796 282180 183802 282192
rect 220906 282180 220912 282192
rect 183796 282152 220912 282180
rect 183796 282140 183802 282152
rect 220906 282140 220912 282152
rect 220964 282140 220970 282192
rect 179506 280780 179512 280832
rect 179564 280820 179570 280832
rect 220814 280820 220820 280832
rect 179564 280792 220820 280820
rect 179564 280780 179570 280792
rect 220814 280780 220820 280792
rect 220872 280780 220878 280832
rect 271138 280780 271144 280832
rect 271196 280820 271202 280832
rect 291194 280820 291200 280832
rect 271196 280792 291200 280820
rect 271196 280780 271202 280792
rect 291194 280780 291200 280792
rect 291252 280780 291258 280832
rect 178126 279420 178132 279472
rect 178184 279460 178190 279472
rect 220906 279460 220912 279472
rect 178184 279432 220912 279460
rect 178184 279420 178190 279432
rect 220906 279420 220912 279432
rect 220964 279420 220970 279472
rect 271230 279420 271236 279472
rect 271288 279460 271294 279472
rect 291746 279460 291752 279472
rect 271288 279432 291752 279460
rect 271288 279420 271294 279432
rect 291746 279420 291752 279432
rect 291804 279420 291810 279472
rect 186406 273912 186412 273964
rect 186464 273952 186470 273964
rect 219802 273952 219808 273964
rect 186464 273924 219808 273952
rect 186464 273912 186470 273924
rect 219802 273912 219808 273924
rect 219860 273912 219866 273964
rect 322934 273912 322940 273964
rect 322992 273952 322998 273964
rect 324038 273952 324044 273964
rect 322992 273924 324044 273952
rect 322992 273912 322998 273924
rect 324038 273912 324044 273924
rect 324096 273952 324102 273964
rect 531314 273952 531320 273964
rect 324096 273924 531320 273952
rect 324096 273912 324102 273924
rect 531314 273912 531320 273924
rect 531372 273912 531378 273964
rect 189258 272484 189264 272536
rect 189316 272524 189322 272536
rect 219894 272524 219900 272536
rect 189316 272496 219900 272524
rect 189316 272484 189322 272496
rect 219894 272484 219900 272496
rect 219952 272484 219958 272536
rect 315482 272484 315488 272536
rect 315540 272524 315546 272536
rect 348878 272524 348884 272536
rect 315540 272496 348884 272524
rect 315540 272484 315546 272496
rect 348878 272484 348884 272496
rect 348936 272524 348942 272536
rect 416774 272524 416780 272536
rect 348936 272496 416780 272524
rect 348936 272484 348942 272496
rect 416774 272484 416780 272496
rect 416832 272484 416838 272536
rect 194778 271124 194784 271176
rect 194836 271164 194842 271176
rect 218606 271164 218612 271176
rect 194836 271136 218612 271164
rect 194836 271124 194842 271136
rect 218606 271124 218612 271136
rect 218664 271124 218670 271176
rect 289630 271124 289636 271176
rect 289688 271164 289694 271176
rect 318334 271164 318340 271176
rect 289688 271136 318340 271164
rect 289688 271124 289694 271136
rect 318334 271124 318340 271136
rect 318392 271124 318398 271176
rect 196158 269764 196164 269816
rect 196216 269804 196222 269816
rect 218882 269804 218888 269816
rect 196216 269776 218888 269804
rect 196216 269764 196222 269776
rect 218882 269764 218888 269776
rect 218940 269764 218946 269816
rect 323670 268200 323676 268252
rect 323728 268240 323734 268252
rect 324130 268240 324136 268252
rect 323728 268212 324136 268240
rect 323728 268200 323734 268212
rect 324130 268200 324136 268212
rect 324188 268200 324194 268252
rect 323670 267724 323676 267776
rect 323728 267764 323734 267776
rect 523126 267764 523132 267776
rect 323728 267736 523132 267764
rect 323728 267724 323734 267736
rect 523126 267724 523132 267736
rect 523184 267724 523190 267776
rect 3050 266364 3056 266416
rect 3108 266404 3114 266416
rect 14458 266404 14464 266416
rect 3108 266376 14464 266404
rect 3108 266364 3114 266376
rect 14458 266364 14464 266376
rect 14516 266364 14522 266416
rect 269114 265616 269120 265668
rect 269172 265656 269178 265668
rect 322658 265656 322664 265668
rect 269172 265628 322664 265656
rect 269172 265616 269178 265628
rect 322658 265616 322664 265628
rect 322716 265616 322722 265668
rect 311342 262148 311348 262200
rect 311400 262188 311406 262200
rect 311710 262188 311716 262200
rect 311400 262160 311716 262188
rect 311400 262148 311406 262160
rect 311710 262148 311716 262160
rect 311768 262148 311774 262200
rect 275370 261468 275376 261520
rect 275428 261508 275434 261520
rect 307202 261508 307208 261520
rect 275428 261480 307208 261508
rect 275428 261468 275434 261480
rect 307202 261468 307208 261480
rect 307260 261468 307266 261520
rect 311342 260924 311348 260976
rect 311400 260964 311406 260976
rect 374086 260964 374092 260976
rect 311400 260936 374092 260964
rect 311400 260924 311406 260936
rect 374086 260924 374092 260936
rect 374144 260924 374150 260976
rect 318518 260856 318524 260908
rect 318576 260896 318582 260908
rect 463694 260896 463700 260908
rect 318576 260868 463700 260896
rect 318576 260856 318582 260868
rect 463694 260856 463700 260868
rect 463752 260856 463758 260908
rect 312906 259428 312912 259480
rect 312964 259468 312970 259480
rect 396074 259468 396080 259480
rect 312964 259440 396080 259468
rect 312964 259428 312970 259440
rect 396074 259428 396080 259440
rect 396132 259428 396138 259480
rect 310330 258068 310336 258120
rect 310388 258108 310394 258120
rect 357434 258108 357440 258120
rect 310388 258080 357440 258108
rect 310388 258068 310394 258080
rect 357434 258068 357440 258080
rect 357492 258068 357498 258120
rect 269114 257388 269120 257440
rect 269172 257428 269178 257440
rect 290734 257428 290740 257440
rect 269172 257400 290740 257428
rect 269172 257388 269178 257400
rect 290734 257388 290740 257400
rect 290792 257388 290798 257440
rect 269574 257320 269580 257372
rect 269632 257360 269638 257372
rect 318610 257360 318616 257372
rect 269632 257332 318616 257360
rect 269632 257320 269638 257332
rect 318610 257320 318616 257332
rect 318668 257360 318674 257372
rect 459554 257360 459560 257372
rect 318668 257332 459560 257360
rect 318668 257320 318674 257332
rect 459554 257320 459560 257332
rect 459612 257320 459618 257372
rect 389174 256816 389180 256828
rect 316006 256788 389180 256816
rect 273806 256708 273812 256760
rect 273864 256748 273870 256760
rect 274634 256748 274640 256760
rect 273864 256720 274640 256748
rect 273864 256708 273870 256720
rect 274634 256708 274640 256720
rect 274692 256708 274698 256760
rect 312906 256708 312912 256760
rect 312964 256748 312970 256760
rect 313090 256748 313096 256760
rect 312964 256720 313096 256748
rect 312964 256708 312970 256720
rect 313090 256708 313096 256720
rect 313148 256748 313154 256760
rect 316006 256748 316034 256788
rect 389174 256776 389180 256788
rect 389232 256776 389238 256828
rect 313148 256720 316034 256748
rect 313148 256708 313154 256720
rect 318150 256708 318156 256760
rect 318208 256748 318214 256760
rect 318702 256748 318708 256760
rect 318208 256720 318708 256748
rect 318208 256708 318214 256720
rect 318702 256708 318708 256720
rect 318760 256748 318766 256760
rect 456794 256748 456800 256760
rect 318760 256720 456800 256748
rect 318760 256708 318766 256720
rect 456794 256708 456800 256720
rect 456852 256708 456858 256760
rect 311526 255348 311532 255400
rect 311584 255388 311590 255400
rect 371234 255388 371240 255400
rect 311584 255360 371240 255388
rect 311584 255348 311590 255360
rect 371234 255348 371240 255360
rect 371292 255348 371298 255400
rect 316954 255280 316960 255332
rect 317012 255320 317018 255332
rect 445754 255320 445760 255332
rect 317012 255292 445760 255320
rect 317012 255280 317018 255292
rect 445754 255280 445760 255292
rect 445812 255280 445818 255332
rect 284202 254532 284208 254584
rect 284260 254572 284266 254584
rect 308490 254572 308496 254584
rect 284260 254544 308496 254572
rect 284260 254532 284266 254544
rect 308490 254532 308496 254544
rect 308548 254532 308554 254584
rect 3418 253920 3424 253972
rect 3476 253960 3482 253972
rect 199930 253960 199936 253972
rect 3476 253932 199936 253960
rect 3476 253920 3482 253932
rect 199930 253920 199936 253932
rect 199988 253960 199994 253972
rect 199988 253932 200114 253960
rect 199988 253920 199994 253932
rect 200086 253892 200114 253932
rect 312722 253920 312728 253972
rect 312780 253960 312786 253972
rect 313182 253960 313188 253972
rect 312780 253932 313188 253960
rect 312780 253920 312786 253932
rect 313182 253920 313188 253932
rect 313240 253960 313246 253972
rect 391934 253960 391940 253972
rect 313240 253932 391940 253960
rect 313240 253920 313246 253932
rect 391934 253920 391940 253932
rect 391992 253920 391998 253972
rect 213270 253892 213276 253904
rect 200086 253864 213276 253892
rect 213270 253852 213276 253864
rect 213328 253852 213334 253904
rect 270402 253308 270408 253360
rect 270460 253348 270466 253360
rect 292482 253348 292488 253360
rect 270460 253320 292488 253348
rect 270460 253308 270466 253320
rect 292482 253308 292488 253320
rect 292540 253308 292546 253360
rect 289722 253240 289728 253292
rect 289780 253280 289786 253292
rect 322382 253280 322388 253292
rect 289780 253252 322388 253280
rect 289780 253240 289786 253252
rect 322382 253240 322388 253252
rect 322440 253240 322446 253292
rect 286870 253172 286876 253224
rect 286928 253212 286934 253224
rect 311434 253212 311440 253224
rect 286928 253184 311440 253212
rect 286928 253172 286934 253184
rect 311434 253172 311440 253184
rect 311492 253172 311498 253224
rect 312814 253172 312820 253224
rect 312872 253212 312878 253224
rect 347590 253212 347596 253224
rect 312872 253184 347596 253212
rect 312872 253172 312878 253184
rect 347590 253172 347596 253184
rect 347648 253212 347654 253224
rect 385034 253212 385040 253224
rect 347648 253184 385040 253212
rect 347648 253172 347654 253184
rect 385034 253172 385040 253184
rect 385092 253172 385098 253224
rect 319714 253036 319720 253088
rect 319772 253076 319778 253088
rect 319990 253076 319996 253088
rect 319772 253048 319996 253076
rect 319772 253036 319778 253048
rect 319990 253036 319996 253048
rect 320048 253036 320054 253088
rect 319714 252628 319720 252680
rect 319772 252668 319778 252680
rect 471238 252668 471244 252680
rect 319772 252640 471244 252668
rect 319772 252628 319778 252640
rect 471238 252628 471244 252640
rect 471296 252628 471302 252680
rect 321462 252560 321468 252612
rect 321520 252600 321526 252612
rect 491294 252600 491300 252612
rect 321520 252572 491300 252600
rect 321520 252560 321526 252572
rect 491294 252560 491300 252572
rect 491352 252560 491358 252612
rect 316770 251812 316776 251864
rect 316828 251852 316834 251864
rect 351454 251852 351460 251864
rect 316828 251824 351460 251852
rect 316828 251812 316834 251824
rect 351454 251812 351460 251824
rect 351512 251852 351518 251864
rect 434714 251852 434720 251864
rect 351512 251824 434720 251852
rect 351512 251812 351518 251824
rect 434714 251812 434720 251824
rect 434772 251812 434778 251864
rect 312998 251268 313004 251320
rect 313056 251308 313062 251320
rect 382274 251308 382280 251320
rect 313056 251280 382280 251308
rect 313056 251268 313062 251280
rect 382274 251268 382280 251280
rect 382332 251268 382338 251320
rect 323762 251200 323768 251252
rect 323820 251240 323826 251252
rect 324222 251240 324228 251252
rect 323820 251212 324228 251240
rect 323820 251200 323826 251212
rect 324222 251200 324228 251212
rect 324280 251240 324286 251252
rect 538214 251240 538220 251252
rect 324280 251212 538220 251240
rect 324280 251200 324286 251212
rect 538214 251200 538220 251212
rect 538272 251200 538278 251252
rect 319806 251132 319812 251184
rect 319864 251172 319870 251184
rect 320082 251172 320088 251184
rect 319864 251144 320088 251172
rect 319864 251132 319870 251144
rect 320082 251132 320088 251144
rect 320140 251132 320146 251184
rect 309042 250452 309048 250504
rect 309100 250492 309106 250504
rect 332594 250492 332600 250504
rect 309100 250464 332600 250492
rect 309100 250452 309106 250464
rect 332594 250452 332600 250464
rect 332652 250452 332658 250504
rect 319806 249772 319812 249824
rect 319864 249812 319870 249824
rect 470594 249812 470600 249824
rect 319864 249784 470600 249812
rect 319864 249772 319870 249784
rect 470594 249772 470600 249784
rect 470652 249772 470658 249824
rect 314562 248548 314568 248600
rect 314620 248588 314626 248600
rect 407114 248588 407120 248600
rect 314620 248560 407120 248588
rect 314620 248548 314626 248560
rect 407114 248548 407120 248560
rect 407172 248548 407178 248600
rect 316034 248480 316040 248532
rect 316092 248520 316098 248532
rect 317138 248520 317144 248532
rect 316092 248492 317144 248520
rect 316092 248480 316098 248492
rect 317138 248480 317144 248492
rect 317196 248520 317202 248532
rect 441614 248520 441620 248532
rect 317196 248492 441620 248520
rect 317196 248480 317202 248492
rect 441614 248480 441620 248492
rect 441672 248480 441678 248532
rect 320082 248412 320088 248464
rect 320140 248452 320146 248464
rect 484394 248452 484400 248464
rect 320140 248424 484400 248452
rect 320140 248412 320146 248424
rect 484394 248412 484400 248424
rect 484452 248412 484458 248464
rect 271046 247868 271052 247920
rect 271104 247908 271110 247920
rect 319898 247908 319904 247920
rect 271104 247880 319904 247908
rect 271104 247868 271110 247880
rect 319898 247868 319904 247880
rect 319956 247868 319962 247920
rect 275738 247800 275744 247852
rect 275796 247840 275802 247852
rect 303246 247840 303252 247852
rect 275796 247812 303252 247840
rect 275796 247800 275802 247812
rect 303246 247800 303252 247812
rect 303304 247800 303310 247852
rect 307662 247800 307668 247852
rect 307720 247840 307726 247852
rect 317414 247840 317420 247852
rect 307720 247812 317420 247840
rect 307720 247800 307726 247812
rect 317414 247800 317420 247812
rect 317472 247800 317478 247852
rect 272242 247732 272248 247784
rect 272300 247772 272306 247784
rect 316034 247772 316040 247784
rect 272300 247744 316040 247772
rect 272300 247732 272306 247744
rect 316034 247732 316040 247744
rect 316092 247732 316098 247784
rect 168558 247664 168564 247716
rect 168616 247704 168622 247716
rect 217226 247704 217232 247716
rect 168616 247676 217232 247704
rect 168616 247664 168622 247676
rect 217226 247664 217232 247676
rect 217284 247664 217290 247716
rect 318242 247664 318248 247716
rect 318300 247704 318306 247716
rect 345934 247704 345940 247716
rect 318300 247676 345940 247704
rect 318300 247664 318306 247676
rect 345934 247664 345940 247676
rect 345992 247704 345998 247716
rect 452654 247704 452660 247716
rect 345992 247676 452660 247704
rect 345992 247664 345998 247676
rect 452654 247664 452660 247676
rect 452712 247664 452718 247716
rect 315390 247052 315396 247104
rect 315448 247092 315454 247104
rect 315850 247092 315856 247104
rect 315448 247064 315856 247092
rect 315448 247052 315454 247064
rect 315850 247052 315856 247064
rect 315908 247092 315914 247104
rect 423766 247092 423772 247104
rect 315908 247064 423772 247092
rect 315908 247052 315914 247064
rect 423766 247052 423772 247064
rect 423824 247052 423830 247104
rect 269758 246372 269764 246424
rect 269816 246412 269822 246424
rect 292206 246412 292212 246424
rect 269816 246384 292212 246412
rect 269816 246372 269822 246384
rect 292206 246372 292212 246384
rect 292264 246372 292270 246424
rect 198826 246304 198832 246356
rect 198884 246344 198890 246356
rect 215938 246344 215944 246356
rect 198884 246316 215944 246344
rect 198884 246304 198890 246316
rect 215938 246304 215944 246316
rect 215996 246304 216002 246356
rect 288986 246304 288992 246356
rect 289044 246344 289050 246356
rect 315298 246344 315304 246356
rect 289044 246316 315304 246344
rect 289044 246304 289050 246316
rect 315298 246304 315304 246316
rect 315356 246304 315362 246356
rect 270862 245692 270868 245744
rect 270920 245732 270926 245744
rect 271506 245732 271512 245744
rect 270920 245704 271512 245732
rect 270920 245692 270926 245704
rect 271506 245692 271512 245704
rect 271564 245692 271570 245744
rect 316678 245624 316684 245676
rect 316736 245664 316742 245676
rect 317230 245664 317236 245676
rect 316736 245636 317236 245664
rect 316736 245624 316742 245636
rect 317230 245624 317236 245636
rect 317288 245664 317294 245676
rect 438854 245664 438860 245676
rect 317288 245636 438860 245664
rect 317288 245624 317294 245636
rect 438854 245624 438860 245636
rect 438912 245624 438918 245676
rect 577590 245556 577596 245608
rect 577648 245596 577654 245608
rect 579614 245596 579620 245608
rect 577648 245568 579620 245596
rect 577648 245556 577654 245568
rect 579614 245556 579620 245568
rect 579672 245556 579678 245608
rect 268930 244944 268936 244996
rect 268988 244984 268994 244996
rect 271230 244984 271236 244996
rect 268988 244956 271236 244984
rect 268988 244944 268994 244956
rect 271230 244944 271236 244956
rect 271288 244944 271294 244996
rect 167086 244876 167092 244928
rect 167144 244916 167150 244928
rect 217318 244916 217324 244928
rect 167144 244888 217324 244916
rect 167144 244876 167150 244888
rect 217318 244876 217324 244888
rect 217376 244876 217382 244928
rect 283466 244876 283472 244928
rect 283524 244916 283530 244928
rect 304534 244916 304540 244928
rect 283524 244888 304540 244916
rect 283524 244876 283530 244888
rect 304534 244876 304540 244888
rect 304592 244876 304598 244928
rect 317322 244468 317328 244520
rect 317380 244508 317386 244520
rect 448514 244508 448520 244520
rect 317380 244480 448520 244508
rect 317380 244468 317386 244480
rect 448514 244468 448520 244480
rect 448572 244468 448578 244520
rect 322382 244400 322388 244452
rect 322440 244440 322446 244452
rect 322842 244440 322848 244452
rect 322440 244412 322848 244440
rect 322440 244400 322446 244412
rect 322842 244400 322848 244412
rect 322900 244440 322906 244452
rect 516134 244440 516140 244452
rect 322900 244412 516140 244440
rect 322900 244400 322906 244412
rect 516134 244400 516140 244412
rect 516192 244400 516198 244452
rect 325142 244332 325148 244384
rect 325200 244372 325206 244384
rect 325510 244372 325516 244384
rect 325200 244344 325516 244372
rect 325200 244332 325206 244344
rect 325510 244332 325516 244344
rect 325568 244372 325574 244384
rect 540974 244372 540980 244384
rect 325568 244344 540980 244372
rect 325568 244332 325574 244344
rect 540974 244332 540980 244344
rect 541032 244332 541038 244384
rect 316862 244264 316868 244316
rect 316920 244304 316926 244316
rect 317322 244304 317328 244316
rect 316920 244276 317328 244304
rect 316920 244264 316926 244276
rect 317322 244264 317328 244276
rect 317380 244264 317386 244316
rect 326338 244264 326344 244316
rect 326396 244304 326402 244316
rect 326982 244304 326988 244316
rect 326396 244276 326988 244304
rect 326396 244264 326402 244276
rect 326982 244264 326988 244276
rect 327040 244304 327046 244316
rect 558914 244304 558920 244316
rect 327040 244276 558920 244304
rect 327040 244264 327046 244276
rect 558914 244264 558920 244276
rect 558972 244264 558978 244316
rect 206462 243584 206468 243636
rect 206520 243624 206526 243636
rect 206646 243624 206652 243636
rect 206520 243596 206652 243624
rect 206520 243584 206526 243596
rect 206646 243584 206652 243596
rect 206704 243584 206710 243636
rect 271782 243516 271788 243568
rect 271840 243556 271846 243568
rect 285030 243556 285036 243568
rect 271840 243528 285036 243556
rect 271840 243516 271846 243528
rect 285030 243516 285036 243528
rect 285088 243516 285094 243568
rect 315298 243040 315304 243092
rect 315356 243080 315362 243092
rect 315942 243080 315948 243092
rect 315356 243052 315948 243080
rect 315356 243040 315362 243052
rect 315942 243040 315948 243052
rect 316000 243080 316006 243092
rect 420914 243080 420920 243092
rect 316000 243052 420920 243080
rect 316000 243040 316006 243052
rect 420914 243040 420920 243052
rect 420972 243040 420978 243092
rect 325050 242972 325056 243024
rect 325108 243012 325114 243024
rect 325602 243012 325608 243024
rect 325108 242984 325608 243012
rect 325108 242972 325114 242984
rect 325602 242972 325608 242984
rect 325660 243012 325666 243024
rect 542998 243012 543004 243024
rect 325660 242984 543004 243012
rect 325660 242972 325666 242984
rect 542998 242972 543004 242984
rect 543056 242972 543062 243024
rect 326246 242904 326252 242956
rect 326304 242944 326310 242956
rect 326890 242944 326896 242956
rect 326304 242916 326896 242944
rect 326304 242904 326310 242916
rect 326890 242904 326896 242916
rect 326948 242944 326954 242956
rect 563054 242944 563060 242956
rect 326948 242916 563060 242944
rect 326948 242904 326954 242916
rect 563054 242904 563060 242916
rect 563112 242904 563118 242956
rect 321462 242836 321468 242888
rect 321520 242876 321526 242888
rect 322290 242876 322296 242888
rect 321520 242848 322296 242876
rect 321520 242836 321526 242848
rect 322290 242836 322296 242848
rect 322348 242836 322354 242888
rect 276198 242292 276204 242344
rect 276256 242332 276262 242344
rect 320910 242332 320916 242344
rect 276256 242304 320916 242332
rect 276256 242292 276262 242304
rect 320910 242292 320916 242304
rect 320968 242292 320974 242344
rect 187878 242224 187884 242276
rect 187936 242264 187942 242276
rect 219986 242264 219992 242276
rect 187936 242236 219992 242264
rect 187936 242224 187942 242236
rect 219986 242224 219992 242236
rect 220044 242224 220050 242276
rect 278774 242224 278780 242276
rect 278832 242264 278838 242276
rect 326246 242264 326252 242276
rect 278832 242236 326252 242264
rect 278832 242224 278838 242236
rect 326246 242224 326252 242236
rect 326304 242224 326310 242276
rect 154390 242156 154396 242208
rect 154448 242196 154454 242208
rect 154448 242168 200114 242196
rect 154448 242156 154454 242168
rect 200086 242060 200114 242168
rect 277854 242156 277860 242208
rect 277912 242196 277918 242208
rect 324958 242196 324964 242208
rect 277912 242168 324964 242196
rect 277912 242156 277918 242168
rect 324958 242156 324964 242168
rect 325016 242156 325022 242208
rect 211982 242060 211988 242072
rect 200086 242032 211988 242060
rect 211982 242020 211988 242032
rect 212040 242060 212046 242072
rect 221090 242060 221096 242072
rect 212040 242032 221096 242060
rect 212040 242020 212046 242032
rect 221090 242020 221096 242032
rect 221148 242020 221154 242072
rect 221182 242020 221188 242072
rect 221240 242060 221246 242072
rect 222470 242060 222476 242072
rect 221240 242032 222476 242060
rect 221240 242020 221246 242032
rect 222470 242020 222476 242032
rect 222528 242020 222534 242072
rect 269022 241612 269028 241664
rect 269080 241652 269086 241664
rect 271138 241652 271144 241664
rect 269080 241624 271144 241652
rect 269080 241612 269086 241624
rect 271138 241612 271144 241624
rect 271196 241612 271202 241664
rect 160002 241544 160008 241596
rect 160060 241584 160066 241596
rect 204898 241584 204904 241596
rect 160060 241556 204904 241584
rect 160060 241544 160066 241556
rect 204898 241544 204904 241556
rect 204956 241544 204962 241596
rect 154482 241476 154488 241528
rect 154540 241516 154546 241528
rect 209038 241516 209044 241528
rect 154540 241488 209044 241516
rect 154540 241476 154546 241488
rect 209038 241476 209044 241488
rect 209096 241476 209102 241528
rect 277394 241476 277400 241528
rect 277452 241516 277458 241528
rect 321462 241516 321468 241528
rect 277452 241488 321468 241516
rect 277452 241476 277458 241488
rect 321462 241476 321468 241488
rect 321520 241476 321526 241528
rect 215754 241408 215760 241460
rect 215812 241448 215818 241460
rect 216306 241448 216312 241460
rect 215812 241420 216312 241448
rect 215812 241408 215818 241420
rect 216306 241408 216312 241420
rect 216364 241408 216370 241460
rect 288434 241408 288440 241460
rect 288492 241448 288498 241460
rect 289630 241448 289636 241460
rect 288492 241420 289636 241448
rect 288492 241408 288498 241420
rect 289630 241408 289636 241420
rect 289688 241408 289694 241460
rect 267550 241340 267556 241392
rect 267608 241380 267614 241392
rect 271138 241380 271144 241392
rect 267608 241352 271144 241380
rect 267608 241340 267614 241352
rect 271138 241340 271144 241352
rect 271196 241340 271202 241392
rect 270586 241272 270592 241324
rect 270644 241312 270650 241324
rect 270954 241312 270960 241324
rect 270644 241284 270960 241312
rect 270644 241272 270650 241284
rect 270954 241272 270960 241284
rect 271012 241272 271018 241324
rect 217594 241204 217600 241256
rect 217652 241244 217658 241256
rect 217652 241216 237374 241244
rect 217652 241204 217658 241216
rect 210418 241136 210424 241188
rect 210476 241176 210482 241188
rect 217686 241176 217692 241188
rect 210476 241148 217692 241176
rect 210476 241136 210482 241148
rect 217686 241136 217692 241148
rect 217744 241176 217750 241188
rect 217744 241148 234384 241176
rect 217744 241136 217750 241148
rect 212258 241000 212264 241052
rect 212316 241040 212322 241052
rect 212316 241012 234292 241040
rect 212316 241000 212322 241012
rect 214926 240864 214932 240916
rect 214984 240904 214990 240916
rect 214984 240876 234108 240904
rect 214984 240864 214990 240876
rect 153102 240796 153108 240848
rect 153160 240836 153166 240848
rect 207750 240836 207756 240848
rect 153160 240808 207756 240836
rect 153160 240796 153166 240808
rect 207750 240796 207756 240808
rect 207808 240836 207814 240848
rect 218606 240836 218612 240848
rect 207808 240808 218612 240836
rect 207808 240796 207814 240808
rect 218606 240796 218612 240808
rect 218664 240796 218670 240848
rect 14458 240728 14464 240780
rect 14516 240768 14522 240780
rect 199378 240768 199384 240780
rect 14516 240740 199384 240768
rect 14516 240728 14522 240740
rect 199378 240728 199384 240740
rect 199436 240728 199442 240780
rect 215266 240672 227898 240700
rect 213362 240388 213368 240440
rect 213420 240428 213426 240440
rect 215266 240428 215294 240672
rect 220538 240592 220544 240644
rect 220596 240632 220602 240644
rect 220596 240604 227714 240632
rect 220596 240592 220602 240604
rect 219158 240456 219164 240508
rect 219216 240496 219222 240508
rect 222194 240496 222200 240508
rect 219216 240468 222200 240496
rect 219216 240456 219222 240468
rect 222194 240456 222200 240468
rect 222252 240456 222258 240508
rect 213420 240400 215294 240428
rect 221016 240400 227622 240428
rect 213420 240388 213426 240400
rect 214834 240320 214840 240372
rect 214892 240360 214898 240372
rect 221016 240360 221044 240400
rect 214892 240332 221044 240360
rect 214892 240320 214898 240332
rect 221090 240320 221096 240372
rect 221148 240360 221154 240372
rect 222194 240360 222200 240372
rect 221148 240332 222200 240360
rect 221148 240320 221154 240332
rect 222194 240320 222200 240332
rect 222252 240320 222258 240372
rect 222286 240320 222292 240372
rect 222344 240360 222350 240372
rect 222344 240332 227530 240360
rect 222344 240320 222350 240332
rect 218606 240252 218612 240304
rect 218664 240292 218670 240304
rect 218664 240264 225782 240292
rect 218664 240252 218670 240264
rect 199930 240184 199936 240236
rect 199988 240224 199994 240236
rect 200298 240224 200304 240236
rect 199988 240196 200304 240224
rect 199988 240184 199994 240196
rect 200298 240184 200304 240196
rect 200356 240184 200362 240236
rect 221366 240184 221372 240236
rect 221424 240224 221430 240236
rect 225754 240224 225782 240264
rect 221424 240196 225690 240224
rect 225754 240196 227438 240224
rect 221424 240184 221430 240196
rect 155678 240116 155684 240168
rect 155736 240156 155742 240168
rect 218698 240156 218704 240168
rect 155736 240128 218704 240156
rect 155736 240116 155742 240128
rect 218698 240116 218704 240128
rect 218756 240116 218762 240168
rect 222194 240116 222200 240168
rect 222252 240156 222258 240168
rect 225662 240156 225690 240196
rect 222252 240128 225598 240156
rect 225662 240128 227346 240156
rect 222252 240116 222258 240128
rect 221274 240048 221280 240100
rect 221332 240088 221338 240100
rect 221332 240060 225322 240088
rect 221332 240048 221338 240060
rect 221458 239980 221464 240032
rect 221516 240020 221522 240032
rect 221516 239992 224126 240020
rect 221516 239980 221522 239992
rect 224098 239964 224126 239992
rect 225294 239964 225322 240060
rect 225570 239964 225598 240128
rect 225662 240060 227254 240088
rect 218698 239912 218704 239964
rect 218756 239952 218762 239964
rect 223068 239952 223074 239964
rect 218756 239924 223074 239952
rect 218756 239912 218762 239924
rect 223068 239912 223074 239924
rect 223126 239912 223132 239964
rect 223344 239912 223350 239964
rect 223402 239912 223408 239964
rect 223712 239912 223718 239964
rect 223770 239912 223776 239964
rect 223896 239912 223902 239964
rect 223954 239912 223960 239964
rect 224080 239912 224086 239964
rect 224138 239912 224144 239964
rect 224172 239912 224178 239964
rect 224230 239912 224236 239964
rect 224540 239912 224546 239964
rect 224598 239912 224604 239964
rect 224816 239912 224822 239964
rect 224874 239912 224880 239964
rect 225276 239952 225282 239964
rect 224926 239924 225282 239952
rect 222286 239844 222292 239896
rect 222344 239884 222350 239896
rect 222792 239884 222798 239896
rect 222344 239856 222798 239884
rect 222344 239844 222350 239856
rect 222792 239844 222798 239856
rect 222850 239844 222856 239896
rect 222884 239844 222890 239896
rect 222942 239844 222948 239896
rect 223160 239844 223166 239896
rect 223218 239884 223224 239896
rect 223218 239856 223298 239884
rect 223218 239844 223224 239856
rect 214558 239776 214564 239828
rect 214616 239816 214622 239828
rect 217594 239816 217600 239828
rect 214616 239788 217600 239816
rect 214616 239776 214622 239788
rect 217594 239776 217600 239788
rect 217652 239776 217658 239828
rect 221090 239776 221096 239828
rect 221148 239816 221154 239828
rect 222700 239816 222706 239828
rect 221148 239788 222706 239816
rect 221148 239776 221154 239788
rect 222700 239776 222706 239788
rect 222758 239776 222764 239828
rect 222902 239816 222930 239844
rect 222902 239788 223022 239816
rect 213086 239708 213092 239760
rect 213144 239748 213150 239760
rect 213144 239720 222792 239748
rect 213144 239708 213150 239720
rect 222764 239692 222792 239720
rect 156506 239640 156512 239692
rect 156564 239680 156570 239692
rect 219986 239680 219992 239692
rect 156564 239652 219992 239680
rect 156564 239640 156570 239652
rect 219986 239640 219992 239652
rect 220044 239640 220050 239692
rect 220078 239640 220084 239692
rect 220136 239640 220142 239692
rect 222746 239640 222752 239692
rect 222804 239640 222810 239692
rect 185210 239572 185216 239624
rect 185268 239612 185274 239624
rect 220096 239612 220124 239640
rect 185268 239584 220124 239612
rect 185268 239572 185274 239584
rect 222286 239572 222292 239624
rect 222344 239612 222350 239624
rect 222994 239612 223022 239788
rect 223114 239640 223120 239692
rect 223172 239680 223178 239692
rect 223270 239680 223298 239856
rect 223172 239652 223298 239680
rect 223172 239640 223178 239652
rect 222344 239584 223022 239612
rect 222344 239572 222350 239584
rect 223206 239572 223212 239624
rect 223264 239612 223270 239624
rect 223362 239612 223390 239912
rect 223436 239844 223442 239896
rect 223494 239884 223500 239896
rect 223620 239884 223626 239896
rect 223494 239844 223528 239884
rect 223500 239624 223528 239844
rect 223592 239844 223626 239884
rect 223678 239844 223684 239896
rect 223592 239680 223620 239844
rect 223730 239760 223758 239912
rect 223666 239708 223672 239760
rect 223724 239720 223758 239760
rect 223914 239760 223942 239912
rect 224190 239828 224218 239912
rect 224264 239844 224270 239896
rect 224322 239844 224328 239896
rect 224126 239776 224132 239828
rect 224184 239788 224218 239828
rect 224184 239776 224190 239788
rect 224282 239760 224310 239844
rect 223914 239720 223948 239760
rect 223724 239708 223730 239720
rect 223942 239708 223948 239720
rect 224000 239708 224006 239760
rect 224218 239708 224224 239760
rect 224276 239720 224310 239760
rect 224276 239708 224282 239720
rect 223850 239680 223856 239692
rect 223592 239652 223856 239680
rect 223592 239624 223620 239652
rect 223850 239640 223856 239652
rect 223908 239640 223914 239692
rect 224034 239640 224040 239692
rect 224092 239680 224098 239692
rect 224558 239680 224586 239912
rect 224834 239816 224862 239912
rect 224696 239788 224862 239816
rect 224696 239692 224724 239788
rect 224926 239692 224954 239924
rect 225276 239912 225282 239924
rect 225334 239912 225340 239964
rect 225460 239912 225466 239964
rect 225518 239912 225524 239964
rect 225552 239912 225558 239964
rect 225610 239912 225616 239964
rect 225478 239884 225506 239912
rect 224092 239652 224586 239680
rect 224092 239640 224098 239652
rect 224678 239640 224684 239692
rect 224736 239640 224742 239692
rect 224862 239640 224868 239692
rect 224920 239652 224954 239692
rect 225156 239856 225506 239884
rect 225662 239884 225690 240060
rect 225754 239992 226610 240020
rect 225754 239964 225782 239992
rect 225736 239912 225742 239964
rect 225794 239912 225800 239964
rect 225828 239912 225834 239964
rect 225886 239912 225892 239964
rect 226012 239912 226018 239964
rect 226070 239912 226076 239964
rect 226288 239912 226294 239964
rect 226346 239912 226352 239964
rect 225846 239884 225874 239912
rect 225662 239856 225874 239884
rect 224920 239640 224926 239652
rect 223264 239584 223390 239612
rect 223264 239572 223270 239584
rect 223482 239572 223488 239624
rect 223540 239572 223546 239624
rect 223574 239572 223580 239624
rect 223632 239572 223638 239624
rect 224310 239572 224316 239624
rect 224368 239612 224374 239624
rect 225156 239612 225184 239856
rect 224368 239584 225184 239612
rect 224368 239572 224374 239584
rect 158438 239504 158444 239556
rect 158496 239544 158502 239556
rect 215018 239544 215024 239556
rect 158496 239516 215024 239544
rect 158496 239504 158502 239516
rect 215018 239504 215024 239516
rect 215076 239544 215082 239556
rect 218882 239544 218888 239556
rect 215076 239516 218888 239544
rect 215076 239504 215082 239516
rect 218882 239504 218888 239516
rect 218940 239504 218946 239556
rect 219066 239504 219072 239556
rect 219124 239544 219130 239556
rect 220630 239544 220636 239556
rect 219124 239516 220636 239544
rect 219124 239504 219130 239516
rect 220630 239504 220636 239516
rect 220688 239504 220694 239556
rect 220722 239504 220728 239556
rect 220780 239544 220786 239556
rect 222746 239544 222752 239556
rect 220780 239516 222752 239544
rect 220780 239504 220786 239516
rect 222746 239504 222752 239516
rect 222804 239504 222810 239556
rect 223850 239504 223856 239556
rect 223908 239544 223914 239556
rect 225046 239544 225052 239556
rect 223908 239516 225052 239544
rect 223908 239504 223914 239516
rect 225046 239504 225052 239516
rect 225104 239504 225110 239556
rect 225156 239544 225184 239584
rect 225230 239572 225236 239624
rect 225288 239612 225294 239624
rect 225782 239612 225788 239624
rect 225288 239584 225788 239612
rect 225288 239572 225294 239584
rect 225782 239572 225788 239584
rect 225840 239612 225846 239624
rect 226030 239612 226058 239912
rect 225840 239584 226058 239612
rect 225840 239572 225846 239584
rect 225506 239544 225512 239556
rect 225156 239516 225512 239544
rect 225506 239504 225512 239516
rect 225564 239504 225570 239556
rect 225690 239504 225696 239556
rect 225748 239544 225754 239556
rect 226306 239544 226334 239912
rect 226472 239844 226478 239896
rect 226530 239844 226536 239896
rect 226490 239760 226518 239844
rect 226582 239760 226610 239992
rect 226858 239992 227162 240020
rect 226858 239964 226886 239992
rect 226840 239912 226846 239964
rect 226898 239912 226904 239964
rect 226656 239844 226662 239896
rect 226714 239844 226720 239896
rect 226426 239708 226432 239760
rect 226484 239720 226518 239760
rect 226484 239708 226490 239720
rect 226564 239708 226570 239760
rect 226622 239708 226628 239760
rect 226674 239680 226702 239844
rect 227134 239748 227162 239992
rect 225748 239516 226334 239544
rect 226628 239652 226702 239680
rect 226904 239720 227162 239748
rect 225748 239504 225754 239516
rect 158530 239436 158536 239488
rect 158588 239476 158594 239488
rect 216306 239476 216312 239488
rect 158588 239448 216312 239476
rect 158588 239436 158594 239448
rect 216306 239436 216312 239448
rect 216364 239476 216370 239488
rect 218606 239476 218612 239488
rect 216364 239448 218612 239476
rect 216364 239436 216370 239448
rect 218606 239436 218612 239448
rect 218664 239436 218670 239488
rect 218698 239436 218704 239488
rect 218756 239476 218762 239488
rect 219342 239476 219348 239488
rect 218756 239448 219348 239476
rect 218756 239436 218762 239448
rect 219342 239436 219348 239448
rect 219400 239436 219406 239488
rect 220906 239436 220912 239488
rect 220964 239476 220970 239488
rect 226628 239476 226656 239652
rect 220964 239448 226656 239476
rect 226904 239476 226932 239720
rect 227226 239680 227254 240060
rect 227318 239952 227346 240128
rect 227410 240088 227438 240196
rect 227502 240156 227530 240332
rect 227594 240224 227622 240400
rect 227686 240292 227714 240604
rect 227870 240360 227898 240672
rect 227870 240332 233050 240360
rect 227686 240264 232958 240292
rect 227594 240196 232406 240224
rect 227502 240128 231854 240156
rect 227410 240060 230566 240088
rect 227962 239992 228358 240020
rect 227962 239964 227990 239992
rect 227392 239952 227398 239964
rect 227318 239924 227398 239952
rect 227392 239912 227398 239924
rect 227450 239912 227456 239964
rect 227576 239912 227582 239964
rect 227634 239952 227640 239964
rect 227634 239912 227668 239952
rect 227944 239912 227950 239964
rect 228002 239912 228008 239964
rect 228036 239912 228042 239964
rect 228094 239952 228100 239964
rect 228220 239952 228226 239964
rect 228094 239912 228128 239952
rect 227410 239884 227438 239912
rect 227410 239856 227576 239884
rect 227438 239680 227444 239692
rect 227226 239652 227444 239680
rect 227438 239640 227444 239652
rect 227496 239640 227502 239692
rect 226978 239572 226984 239624
rect 227036 239612 227042 239624
rect 227548 239612 227576 239856
rect 227640 239624 227668 239912
rect 228100 239692 228128 239912
rect 228192 239912 228226 239952
rect 228278 239912 228284 239964
rect 228082 239640 228088 239692
rect 228140 239640 228146 239692
rect 227036 239584 227576 239612
rect 227036 239572 227042 239584
rect 227622 239572 227628 239624
rect 227680 239572 227686 239624
rect 228192 239612 228220 239912
rect 228008 239584 228220 239612
rect 227070 239476 227076 239488
rect 226904 239448 227076 239476
rect 220964 239436 220970 239448
rect 227070 239436 227076 239448
rect 227128 239476 227134 239488
rect 227438 239476 227444 239488
rect 227128 239448 227444 239476
rect 227128 239436 227134 239448
rect 227438 239436 227444 239448
rect 227496 239436 227502 239488
rect 228008 239476 228036 239584
rect 228330 239556 228358 239992
rect 230538 239964 230566 240060
rect 228404 239912 228410 239964
rect 228462 239912 228468 239964
rect 228496 239912 228502 239964
rect 228554 239952 228560 239964
rect 229048 239952 229054 239964
rect 228554 239924 228910 239952
rect 228554 239912 228560 239924
rect 228422 239612 228450 239912
rect 228588 239844 228594 239896
rect 228646 239844 228652 239896
rect 228680 239844 228686 239896
rect 228738 239844 228744 239896
rect 228772 239844 228778 239896
rect 228830 239844 228836 239896
rect 228606 239816 228634 239844
rect 228560 239788 228634 239816
rect 228560 239624 228588 239788
rect 228698 239760 228726 239844
rect 228634 239708 228640 239760
rect 228692 239720 228726 239760
rect 228692 239708 228698 239720
rect 228422 239584 228496 239612
rect 228330 239516 228364 239556
rect 228358 239504 228364 239516
rect 228416 239504 228422 239556
rect 228082 239476 228088 239488
rect 228008 239448 228088 239476
rect 228082 239436 228088 239448
rect 228140 239436 228146 239488
rect 228468 239476 228496 239584
rect 228542 239572 228548 239624
rect 228600 239572 228606 239624
rect 228238 239448 228496 239476
rect 3326 239368 3332 239420
rect 3384 239408 3390 239420
rect 198918 239408 198924 239420
rect 3384 239380 198924 239408
rect 3384 239368 3390 239380
rect 198918 239368 198924 239380
rect 198976 239408 198982 239420
rect 216030 239408 216036 239420
rect 198976 239380 216036 239408
rect 198976 239368 198982 239380
rect 216030 239368 216036 239380
rect 216088 239368 216094 239420
rect 217410 239368 217416 239420
rect 217468 239408 217474 239420
rect 217594 239408 217600 239420
rect 217468 239380 217600 239408
rect 217468 239368 217474 239380
rect 217594 239368 217600 239380
rect 217652 239368 217658 239420
rect 226426 239408 226432 239420
rect 219360 239380 226432 239408
rect 213638 239300 213644 239352
rect 213696 239340 213702 239352
rect 217870 239340 217876 239352
rect 213696 239312 217876 239340
rect 213696 239300 213702 239312
rect 217870 239300 217876 239312
rect 217928 239340 217934 239352
rect 219360 239340 219388 239380
rect 226426 239368 226432 239380
rect 226484 239368 226490 239420
rect 227898 239368 227904 239420
rect 227956 239408 227962 239420
rect 228238 239408 228266 239448
rect 228634 239436 228640 239488
rect 228692 239476 228698 239488
rect 228790 239476 228818 239844
rect 228882 239544 228910 239924
rect 229020 239912 229054 239952
rect 229106 239912 229112 239964
rect 229140 239912 229146 239964
rect 229198 239912 229204 239964
rect 229416 239952 229422 239964
rect 229388 239912 229422 239952
rect 229474 239912 229480 239964
rect 229508 239912 229514 239964
rect 229566 239912 229572 239964
rect 229600 239912 229606 239964
rect 229658 239912 229664 239964
rect 229968 239912 229974 239964
rect 230026 239912 230032 239964
rect 230244 239912 230250 239964
rect 230302 239912 230308 239964
rect 230520 239912 230526 239964
rect 230578 239912 230584 239964
rect 231256 239912 231262 239964
rect 231314 239952 231320 239964
rect 231440 239952 231446 239964
rect 231314 239912 231348 239952
rect 229020 239680 229048 239912
rect 229158 239884 229186 239912
rect 229112 239856 229186 239884
rect 229112 239760 229140 239856
rect 229388 239816 229416 239912
rect 229526 239828 229554 239912
rect 229296 239788 229416 239816
rect 229094 239708 229100 239760
rect 229152 239708 229158 239760
rect 229296 239692 229324 239788
rect 229462 239776 229468 239828
rect 229520 239788 229554 239828
rect 229520 239776 229526 239788
rect 229186 239680 229192 239692
rect 229020 239652 229192 239680
rect 229186 239640 229192 239652
rect 229244 239640 229250 239692
rect 229278 239640 229284 239692
rect 229336 239640 229342 239692
rect 229618 239680 229646 239912
rect 229876 239844 229882 239896
rect 229934 239844 229940 239896
rect 229738 239708 229744 239760
rect 229796 239748 229802 239760
rect 229894 239748 229922 239844
rect 229796 239720 229922 239748
rect 229796 239708 229802 239720
rect 229986 239692 230014 239912
rect 229830 239680 229836 239692
rect 229618 239652 229836 239680
rect 229830 239640 229836 239652
rect 229888 239640 229894 239692
rect 229922 239640 229928 239692
rect 229980 239652 230014 239692
rect 230262 239680 230290 239912
rect 230796 239844 230802 239896
rect 230854 239844 230860 239896
rect 230888 239844 230894 239896
rect 230946 239844 230952 239896
rect 230980 239844 230986 239896
rect 231038 239844 231044 239896
rect 231072 239844 231078 239896
rect 231130 239844 231136 239896
rect 230814 239816 230842 239844
rect 230400 239788 230842 239816
rect 230400 239760 230428 239788
rect 230906 239760 230934 239844
rect 230382 239708 230388 239760
rect 230440 239708 230446 239760
rect 230842 239708 230848 239760
rect 230900 239720 230934 239760
rect 230900 239708 230906 239720
rect 230262 239652 230428 239680
rect 229980 239640 229986 239652
rect 229646 239572 229652 239624
rect 229704 239612 229710 239624
rect 230290 239612 230296 239624
rect 229704 239584 230296 239612
rect 229704 239572 229710 239584
rect 230290 239572 230296 239584
rect 230348 239572 230354 239624
rect 229278 239544 229284 239556
rect 228882 239516 229284 239544
rect 229278 239504 229284 239516
rect 229336 239504 229342 239556
rect 230198 239504 230204 239556
rect 230256 239544 230262 239556
rect 230400 239544 230428 239652
rect 230842 239572 230848 239624
rect 230900 239612 230906 239624
rect 230998 239612 231026 239844
rect 231090 239748 231118 239844
rect 231210 239748 231216 239760
rect 231090 239720 231216 239748
rect 231210 239708 231216 239720
rect 231268 239708 231274 239760
rect 231320 239692 231348 239912
rect 231412 239912 231446 239952
rect 231498 239912 231504 239964
rect 231532 239912 231538 239964
rect 231590 239912 231596 239964
rect 231716 239912 231722 239964
rect 231774 239912 231780 239964
rect 231302 239640 231308 239692
rect 231360 239640 231366 239692
rect 230900 239584 231026 239612
rect 230900 239572 230906 239584
rect 231118 239572 231124 239624
rect 231176 239612 231182 239624
rect 231412 239612 231440 239912
rect 231550 239624 231578 239912
rect 231176 239584 231440 239612
rect 231176 239572 231182 239584
rect 231486 239572 231492 239624
rect 231544 239584 231578 239624
rect 231734 239624 231762 239912
rect 231826 239680 231854 240128
rect 232378 239964 232406 240196
rect 231992 239912 231998 239964
rect 232050 239912 232056 239964
rect 232084 239912 232090 239964
rect 232142 239952 232148 239964
rect 232142 239912 232176 239952
rect 232268 239912 232274 239964
rect 232326 239912 232332 239964
rect 232360 239912 232366 239964
rect 232418 239912 232424 239964
rect 232728 239912 232734 239964
rect 232786 239912 232792 239964
rect 232820 239912 232826 239964
rect 232878 239912 232884 239964
rect 232010 239884 232038 239912
rect 232010 239856 232084 239884
rect 232056 239828 232084 239856
rect 232038 239776 232044 239828
rect 232096 239776 232102 239828
rect 232148 239760 232176 239912
rect 232286 239884 232314 239912
rect 232286 239856 232360 239884
rect 232332 239828 232360 239856
rect 232314 239776 232320 239828
rect 232372 239776 232378 239828
rect 232130 239708 232136 239760
rect 232188 239708 232194 239760
rect 231826 239652 232636 239680
rect 232608 239624 232636 239652
rect 231734 239584 231768 239624
rect 231544 239572 231550 239584
rect 231762 239572 231768 239584
rect 231820 239572 231826 239624
rect 232590 239572 232596 239624
rect 232648 239572 232654 239624
rect 230256 239516 230428 239544
rect 230256 239504 230262 239516
rect 230658 239504 230664 239556
rect 230716 239544 230722 239556
rect 232746 239544 232774 239912
rect 230716 239516 232774 239544
rect 230716 239504 230722 239516
rect 230290 239476 230296 239488
rect 228692 239448 230296 239476
rect 228692 239436 228698 239448
rect 230290 239436 230296 239448
rect 230348 239436 230354 239488
rect 231854 239436 231860 239488
rect 231912 239476 231918 239488
rect 232838 239476 232866 239912
rect 232930 239544 232958 240264
rect 233022 240020 233050 240332
rect 234080 240156 234108 240876
rect 234264 240224 234292 241012
rect 234356 240564 234384 241148
rect 237346 240632 237374 241216
rect 267550 241176 267556 241188
rect 248248 241148 267556 241176
rect 237346 240604 238938 240632
rect 234356 240536 237374 240564
rect 234264 240196 235166 240224
rect 235138 240156 235166 240196
rect 237346 240156 237374 240536
rect 238910 240224 238938 240604
rect 248248 240360 248276 241148
rect 267550 241136 267556 241148
rect 267608 241136 267614 241188
rect 269206 241108 269212 241120
rect 246454 240332 248276 240360
rect 248340 241080 269212 241108
rect 238910 240196 240502 240224
rect 234080 240128 235074 240156
rect 235138 240128 237006 240156
rect 237346 240128 239398 240156
rect 234034 240060 234706 240088
rect 233022 239992 233418 240020
rect 233390 239964 233418 239992
rect 234034 239964 234062 240060
rect 233096 239912 233102 239964
rect 233154 239912 233160 239964
rect 233372 239912 233378 239964
rect 233430 239912 233436 239964
rect 233464 239912 233470 239964
rect 233522 239912 233528 239964
rect 233648 239952 233654 239964
rect 233620 239912 233654 239952
rect 233706 239912 233712 239964
rect 233740 239912 233746 239964
rect 233798 239912 233804 239964
rect 234016 239912 234022 239964
rect 234074 239912 234080 239964
rect 234200 239912 234206 239964
rect 234258 239912 234264 239964
rect 234568 239912 234574 239964
rect 234626 239912 234632 239964
rect 233114 239624 233142 239912
rect 233482 239884 233510 239912
rect 233620 239884 233648 239912
rect 233758 239884 233786 239912
rect 233436 239856 233510 239884
rect 233574 239856 233648 239884
rect 233712 239856 233786 239884
rect 233436 239828 233464 239856
rect 233418 239776 233424 239828
rect 233476 239776 233482 239828
rect 233574 239748 233602 239856
rect 233712 239828 233740 239856
rect 233924 239844 233930 239896
rect 233982 239844 233988 239896
rect 233694 239776 233700 239828
rect 233752 239776 233758 239828
rect 233252 239720 233602 239748
rect 233252 239624 233280 239720
rect 233942 239692 233970 239844
rect 234218 239760 234246 239912
rect 234384 239844 234390 239896
rect 234442 239844 234448 239896
rect 234218 239720 234252 239760
rect 234246 239708 234252 239720
rect 234304 239708 234310 239760
rect 234402 239692 234430 239844
rect 233942 239652 233976 239692
rect 233970 239640 233976 239652
rect 234028 239640 234034 239692
rect 234338 239640 234344 239692
rect 234396 239652 234430 239692
rect 234396 239640 234402 239652
rect 233050 239572 233056 239624
rect 233108 239584 233142 239624
rect 233108 239572 233114 239584
rect 233234 239572 233240 239624
rect 233292 239572 233298 239624
rect 234154 239612 234160 239624
rect 233344 239584 234160 239612
rect 233344 239544 233372 239584
rect 234154 239572 234160 239584
rect 234212 239572 234218 239624
rect 234430 239572 234436 239624
rect 234488 239612 234494 239624
rect 234586 239612 234614 239912
rect 234488 239584 234614 239612
rect 234678 239612 234706 240060
rect 235046 240020 235074 240128
rect 234770 239992 235074 240020
rect 236196 239992 236638 240020
rect 234770 239964 234798 239992
rect 234752 239912 234758 239964
rect 234810 239912 234816 239964
rect 235028 239912 235034 239964
rect 235086 239952 235092 239964
rect 235086 239912 235120 239952
rect 235212 239912 235218 239964
rect 235270 239912 235276 239964
rect 235396 239912 235402 239964
rect 235454 239952 235460 239964
rect 235454 239912 235488 239952
rect 235580 239912 235586 239964
rect 235638 239912 235644 239964
rect 235672 239912 235678 239964
rect 235730 239912 235736 239964
rect 235764 239912 235770 239964
rect 235822 239912 235828 239964
rect 235948 239912 235954 239964
rect 236006 239912 236012 239964
rect 234890 239612 234896 239624
rect 234678 239584 234896 239612
rect 234488 239572 234494 239584
rect 234890 239572 234896 239584
rect 234948 239572 234954 239624
rect 232930 239516 233372 239544
rect 233418 239504 233424 239556
rect 233476 239544 233482 239556
rect 235092 239544 235120 239912
rect 235230 239760 235258 239912
rect 235230 239720 235264 239760
rect 235258 239708 235264 239720
rect 235316 239708 235322 239760
rect 235460 239692 235488 239912
rect 235442 239640 235448 239692
rect 235500 239640 235506 239692
rect 235166 239572 235172 239624
rect 235224 239612 235230 239624
rect 235598 239612 235626 239912
rect 235224 239584 235626 239612
rect 235224 239572 235230 239584
rect 233476 239516 235120 239544
rect 233476 239504 233482 239516
rect 235534 239504 235540 239556
rect 235592 239544 235598 239556
rect 235690 239544 235718 239912
rect 235592 239516 235718 239544
rect 235782 239544 235810 239912
rect 235966 239760 235994 239912
rect 236040 239844 236046 239896
rect 236098 239884 236104 239896
rect 236098 239844 236132 239884
rect 235966 239720 236000 239760
rect 235994 239708 236000 239720
rect 236052 239708 236058 239760
rect 236104 239624 236132 239844
rect 236086 239572 236092 239624
rect 236144 239572 236150 239624
rect 236196 239544 236224 239992
rect 236610 239964 236638 239992
rect 236592 239912 236598 239964
rect 236650 239912 236656 239964
rect 236868 239952 236874 239964
rect 236794 239924 236874 239952
rect 236684 239844 236690 239896
rect 236742 239844 236748 239896
rect 236702 239680 236730 239844
rect 236564 239652 236730 239680
rect 236454 239544 236460 239556
rect 235782 239516 236132 239544
rect 236196 239516 236460 239544
rect 235592 239504 235598 239516
rect 235994 239476 236000 239488
rect 231912 239448 236000 239476
rect 231912 239436 231918 239448
rect 235994 239436 236000 239448
rect 236052 239436 236058 239488
rect 227956 239380 228266 239408
rect 227956 239368 227962 239380
rect 228726 239368 228732 239420
rect 228784 239408 228790 239420
rect 229002 239408 229008 239420
rect 228784 239380 229008 239408
rect 228784 239368 228790 239380
rect 229002 239368 229008 239380
rect 229060 239368 229066 239420
rect 229094 239368 229100 239420
rect 229152 239408 229158 239420
rect 233418 239408 233424 239420
rect 229152 239380 233424 239408
rect 229152 239368 229158 239380
rect 233418 239368 233424 239380
rect 233476 239368 233482 239420
rect 233786 239368 233792 239420
rect 233844 239408 233850 239420
rect 235534 239408 235540 239420
rect 233844 239380 235540 239408
rect 233844 239368 233850 239380
rect 235534 239368 235540 239380
rect 235592 239368 235598 239420
rect 235718 239368 235724 239420
rect 235776 239408 235782 239420
rect 236104 239408 236132 239516
rect 236454 239504 236460 239516
rect 236512 239504 236518 239556
rect 235776 239380 236132 239408
rect 235776 239368 235782 239380
rect 217928 239312 219388 239340
rect 217928 239300 217934 239312
rect 222010 239300 222016 239352
rect 222068 239340 222074 239352
rect 223390 239340 223396 239352
rect 222068 239312 223396 239340
rect 222068 239300 222074 239312
rect 223390 239300 223396 239312
rect 223448 239300 223454 239352
rect 232774 239300 232780 239352
rect 232832 239340 232838 239352
rect 236564 239340 236592 239652
rect 236794 239624 236822 239924
rect 236868 239912 236874 239924
rect 236926 239912 236932 239964
rect 236978 239828 237006 240128
rect 237208 240060 237558 240088
rect 237052 239912 237058 239964
rect 237110 239912 237116 239964
rect 237070 239884 237098 239912
rect 237070 239856 237144 239884
rect 236978 239788 237012 239828
rect 237006 239776 237012 239788
rect 237064 239776 237070 239828
rect 236914 239708 236920 239760
rect 236972 239708 236978 239760
rect 237116 239748 237144 239856
rect 237024 239720 237144 239748
rect 236932 239624 236960 239708
rect 236794 239584 236828 239624
rect 236822 239572 236828 239584
rect 236880 239572 236886 239624
rect 236914 239572 236920 239624
rect 236972 239572 236978 239624
rect 237024 239556 237052 239720
rect 237006 239504 237012 239556
rect 237064 239504 237070 239556
rect 237208 239544 237236 240060
rect 237530 239964 237558 240060
rect 239370 239964 239398 240128
rect 240474 239964 240502 240196
rect 246454 240088 246482 240332
rect 245994 240060 246482 240088
rect 244798 239992 245194 240020
rect 244798 239964 244826 239992
rect 237420 239912 237426 239964
rect 237478 239912 237484 239964
rect 237512 239912 237518 239964
rect 237570 239912 237576 239964
rect 237788 239912 237794 239964
rect 237846 239912 237852 239964
rect 238156 239912 238162 239964
rect 238214 239912 238220 239964
rect 238248 239912 238254 239964
rect 238306 239912 238312 239964
rect 238432 239912 238438 239964
rect 238490 239912 238496 239964
rect 238616 239912 238622 239964
rect 238674 239952 238680 239964
rect 239260 239952 239266 239964
rect 238674 239924 238846 239952
rect 238674 239912 238680 239924
rect 237438 239816 237466 239912
rect 237604 239844 237610 239896
rect 237662 239884 237668 239896
rect 237662 239844 237696 239884
rect 237438 239788 237604 239816
rect 237576 239692 237604 239788
rect 237558 239640 237564 239692
rect 237616 239640 237622 239692
rect 237466 239572 237472 239624
rect 237524 239612 237530 239624
rect 237668 239612 237696 239844
rect 237524 239584 237696 239612
rect 237806 239624 237834 239912
rect 237880 239844 237886 239896
rect 237938 239844 237944 239896
rect 237972 239844 237978 239896
rect 238030 239884 238036 239896
rect 238030 239844 238064 239884
rect 237898 239692 237926 239844
rect 238036 239692 238064 239844
rect 237898 239652 237932 239692
rect 237926 239640 237932 239652
rect 237984 239640 237990 239692
rect 238018 239640 238024 239692
rect 238076 239640 238082 239692
rect 237806 239584 237840 239624
rect 237524 239572 237530 239584
rect 237834 239572 237840 239584
rect 237892 239572 237898 239624
rect 237116 239516 237236 239544
rect 232832 239312 236592 239340
rect 232832 239300 232838 239312
rect 237006 239300 237012 239352
rect 237064 239340 237070 239352
rect 237116 239340 237144 239516
rect 237650 239504 237656 239556
rect 237708 239544 237714 239556
rect 238174 239544 238202 239912
rect 238266 239692 238294 239912
rect 238450 239884 238478 239912
rect 238404 239856 238478 239884
rect 238266 239652 238300 239692
rect 238294 239640 238300 239652
rect 238352 239640 238358 239692
rect 237708 239516 238202 239544
rect 237708 239504 237714 239516
rect 238110 239436 238116 239488
rect 238168 239436 238174 239488
rect 237282 239368 237288 239420
rect 237340 239408 237346 239420
rect 238128 239408 238156 239436
rect 237340 239380 238156 239408
rect 237340 239368 237346 239380
rect 237064 239312 237144 239340
rect 237064 239300 237070 239312
rect 237374 239300 237380 239352
rect 237432 239340 237438 239352
rect 238294 239340 238300 239352
rect 237432 239312 238300 239340
rect 237432 239300 237438 239312
rect 238294 239300 238300 239312
rect 238352 239340 238358 239352
rect 238404 239340 238432 239856
rect 238524 239844 238530 239896
rect 238582 239844 238588 239896
rect 238708 239884 238714 239896
rect 238680 239844 238714 239884
rect 238766 239844 238772 239896
rect 238542 239760 238570 239844
rect 238478 239708 238484 239760
rect 238536 239720 238570 239760
rect 238536 239708 238542 239720
rect 238680 239692 238708 239844
rect 238818 239816 238846 239924
rect 238772 239788 238846 239816
rect 238956 239924 239266 239952
rect 238662 239640 238668 239692
rect 238720 239640 238726 239692
rect 238570 239572 238576 239624
rect 238628 239612 238634 239624
rect 238772 239612 238800 239788
rect 238628 239584 238800 239612
rect 238628 239572 238634 239584
rect 238956 239488 238984 239924
rect 239260 239912 239266 239924
rect 239318 239912 239324 239964
rect 239352 239912 239358 239964
rect 239410 239912 239416 239964
rect 239444 239912 239450 239964
rect 239502 239912 239508 239964
rect 239812 239952 239818 239964
rect 239784 239912 239818 239952
rect 239870 239912 239876 239964
rect 239996 239912 240002 239964
rect 240054 239912 240060 239964
rect 240180 239912 240186 239964
rect 240238 239912 240244 239964
rect 240456 239912 240462 239964
rect 240514 239912 240520 239964
rect 240732 239912 240738 239964
rect 240790 239912 240796 239964
rect 240916 239952 240922 239964
rect 240888 239912 240922 239952
rect 240974 239912 240980 239964
rect 241008 239912 241014 239964
rect 241066 239912 241072 239964
rect 241468 239952 241474 239964
rect 241210 239924 241474 239952
rect 239076 239884 239082 239896
rect 239048 239844 239082 239884
rect 239134 239844 239140 239896
rect 239048 239612 239076 239844
rect 239214 239776 239220 239828
rect 239272 239776 239278 239828
rect 239462 239816 239490 239912
rect 239324 239788 239490 239816
rect 239232 239692 239260 239776
rect 239324 239760 239352 239788
rect 239306 239708 239312 239760
rect 239364 239708 239370 239760
rect 239214 239640 239220 239692
rect 239272 239640 239278 239692
rect 239582 239612 239588 239624
rect 239048 239584 239588 239612
rect 239582 239572 239588 239584
rect 239640 239572 239646 239624
rect 238938 239436 238944 239488
rect 238996 239436 239002 239488
rect 239306 239436 239312 239488
rect 239364 239476 239370 239488
rect 239784 239476 239812 239912
rect 240014 239692 240042 239912
rect 240198 239748 240226 239912
rect 240640 239844 240646 239896
rect 240698 239844 240704 239896
rect 240318 239748 240324 239760
rect 240198 239720 240324 239748
rect 240318 239708 240324 239720
rect 240376 239708 240382 239760
rect 240658 239692 240686 239844
rect 240750 239760 240778 239912
rect 240888 239760 240916 239912
rect 241026 239828 241054 239912
rect 240962 239776 240968 239828
rect 241020 239788 241054 239828
rect 241020 239776 241026 239788
rect 240750 239720 240784 239760
rect 240778 239708 240784 239720
rect 240836 239708 240842 239760
rect 240870 239708 240876 239760
rect 240928 239708 240934 239760
rect 241210 239692 241238 239924
rect 241468 239912 241474 239924
rect 241526 239912 241532 239964
rect 241560 239912 241566 239964
rect 241618 239912 241624 239964
rect 241652 239912 241658 239964
rect 241710 239912 241716 239964
rect 241744 239912 241750 239964
rect 241802 239912 241808 239964
rect 241928 239912 241934 239964
rect 241986 239912 241992 239964
rect 242296 239912 242302 239964
rect 242354 239912 242360 239964
rect 242388 239912 242394 239964
rect 242446 239912 242452 239964
rect 242480 239912 242486 239964
rect 242538 239912 242544 239964
rect 242848 239952 242854 239964
rect 242820 239912 242854 239952
rect 242906 239912 242912 239964
rect 243032 239912 243038 239964
rect 243090 239912 243096 239964
rect 243308 239912 243314 239964
rect 243366 239912 243372 239964
rect 243492 239912 243498 239964
rect 243550 239912 243556 239964
rect 244136 239912 244142 239964
rect 244194 239912 244200 239964
rect 244412 239952 244418 239964
rect 244292 239924 244418 239952
rect 241284 239844 241290 239896
rect 241342 239844 241348 239896
rect 241578 239884 241606 239912
rect 241532 239856 241606 239884
rect 241302 239748 241330 239844
rect 241302 239720 241376 239748
rect 240014 239652 240048 239692
rect 240042 239640 240048 239652
rect 240100 239640 240106 239692
rect 240658 239652 240692 239692
rect 240686 239640 240692 239652
rect 240744 239640 240750 239692
rect 241210 239652 241244 239692
rect 241238 239640 241244 239652
rect 241296 239640 241302 239692
rect 239364 239448 239812 239476
rect 239364 239436 239370 239448
rect 240594 239436 240600 239488
rect 240652 239476 240658 239488
rect 241348 239476 241376 239720
rect 241532 239692 241560 239856
rect 241670 239692 241698 239912
rect 241762 239760 241790 239912
rect 241762 239720 241796 239760
rect 241790 239708 241796 239720
rect 241848 239708 241854 239760
rect 241514 239640 241520 239692
rect 241572 239640 241578 239692
rect 241606 239640 241612 239692
rect 241664 239652 241698 239692
rect 241664 239640 241670 239652
rect 241946 239556 241974 239912
rect 242314 239612 242342 239912
rect 242176 239584 242342 239612
rect 241946 239516 241980 239556
rect 241974 239504 241980 239516
rect 242032 239504 242038 239556
rect 240652 239448 241376 239476
rect 240652 239436 240658 239448
rect 238754 239368 238760 239420
rect 238812 239408 238818 239420
rect 242176 239408 242204 239584
rect 242406 239556 242434 239912
rect 242342 239504 242348 239556
rect 242400 239516 242434 239556
rect 242400 239504 242406 239516
rect 242498 239488 242526 239912
rect 242820 239556 242848 239912
rect 243050 239680 243078 239912
rect 243170 239680 243176 239692
rect 243050 239652 243176 239680
rect 243170 239640 243176 239652
rect 243228 239640 243234 239692
rect 243326 239624 243354 239912
rect 243262 239572 243268 239624
rect 243320 239584 243354 239624
rect 243320 239572 243326 239584
rect 242802 239504 242808 239556
rect 242860 239504 242866 239556
rect 242894 239504 242900 239556
rect 242952 239544 242958 239556
rect 243510 239544 243538 239912
rect 243676 239844 243682 239896
rect 243734 239844 243740 239896
rect 243694 239760 243722 239844
rect 244154 239816 244182 239912
rect 243630 239708 243636 239760
rect 243688 239720 243722 239760
rect 244016 239788 244182 239816
rect 243688 239708 243694 239720
rect 242952 239516 243538 239544
rect 242952 239504 242958 239516
rect 244016 239488 244044 239788
rect 244292 239748 244320 239924
rect 244412 239912 244418 239924
rect 244470 239912 244476 239964
rect 244596 239952 244602 239964
rect 244568 239912 244602 239952
rect 244654 239912 244660 239964
rect 244688 239912 244694 239964
rect 244746 239912 244752 239964
rect 244780 239912 244786 239964
rect 244838 239912 244844 239964
rect 245056 239912 245062 239964
rect 245114 239912 245120 239964
rect 244568 239760 244596 239912
rect 244706 239884 244734 239912
rect 245074 239884 245102 239912
rect 244660 239856 244734 239884
rect 244844 239856 245102 239884
rect 244200 239720 244320 239748
rect 242434 239436 242440 239488
rect 242492 239448 242526 239488
rect 242492 239436 242498 239448
rect 243998 239436 244004 239488
rect 244056 239436 244062 239488
rect 238812 239380 242204 239408
rect 238812 239368 238818 239380
rect 242710 239368 242716 239420
rect 242768 239408 242774 239420
rect 242986 239408 242992 239420
rect 242768 239380 242992 239408
rect 242768 239368 242774 239380
rect 242986 239368 242992 239380
rect 243044 239368 243050 239420
rect 238352 239312 238432 239340
rect 238352 239300 238358 239312
rect 238662 239300 238668 239352
rect 238720 239340 238726 239352
rect 239030 239340 239036 239352
rect 238720 239312 239036 239340
rect 238720 239300 238726 239312
rect 239030 239300 239036 239312
rect 239088 239300 239094 239352
rect 241514 239340 241520 239352
rect 240520 239312 241520 239340
rect 218974 239232 218980 239284
rect 219032 239272 219038 239284
rect 240520 239272 240548 239312
rect 241514 239300 241520 239312
rect 241572 239300 241578 239352
rect 243262 239300 243268 239352
rect 243320 239340 243326 239352
rect 244200 239340 244228 239720
rect 244550 239708 244556 239760
rect 244608 239708 244614 239760
rect 244660 239692 244688 239856
rect 244734 239776 244740 239828
rect 244792 239816 244798 239828
rect 244844 239816 244872 239856
rect 244964 239816 244970 239828
rect 244792 239788 244872 239816
rect 244792 239776 244798 239788
rect 244936 239776 244970 239816
rect 245022 239776 245028 239828
rect 244936 239692 244964 239776
rect 245166 239748 245194 239992
rect 245994 239964 246022 240060
rect 248340 240020 248368 241080
rect 269206 241068 269212 241080
rect 269264 241068 269270 241120
rect 272242 241040 272248 241052
rect 256896 241012 272248 241040
rect 251146 240196 253704 240224
rect 246316 239992 248368 240020
rect 248938 239992 250530 240020
rect 245332 239912 245338 239964
rect 245390 239912 245396 239964
rect 245424 239912 245430 239964
rect 245482 239912 245488 239964
rect 245700 239912 245706 239964
rect 245758 239912 245764 239964
rect 245976 239912 245982 239964
rect 246034 239912 246040 239964
rect 246160 239912 246166 239964
rect 246218 239912 246224 239964
rect 245028 239720 245194 239748
rect 244642 239640 244648 239692
rect 244700 239640 244706 239692
rect 244918 239640 244924 239692
rect 244976 239640 244982 239692
rect 245028 239544 245056 239720
rect 245350 239624 245378 239912
rect 245286 239572 245292 239624
rect 245344 239584 245378 239624
rect 245442 239624 245470 239912
rect 245718 239760 245746 239912
rect 245792 239844 245798 239896
rect 245850 239884 245856 239896
rect 245850 239844 245884 239884
rect 245856 239760 245884 239844
rect 246178 239760 246206 239912
rect 245718 239720 245752 239760
rect 245746 239708 245752 239720
rect 245804 239708 245810 239760
rect 245838 239708 245844 239760
rect 245896 239708 245902 239760
rect 246114 239708 246120 239760
rect 246172 239720 246206 239760
rect 246172 239708 246178 239720
rect 246316 239692 246344 239992
rect 246620 239912 246626 239964
rect 246678 239912 246684 239964
rect 246712 239912 246718 239964
rect 246770 239912 246776 239964
rect 247356 239912 247362 239964
rect 247414 239912 247420 239964
rect 247724 239912 247730 239964
rect 247782 239912 247788 239964
rect 247816 239912 247822 239964
rect 247874 239912 247880 239964
rect 247908 239912 247914 239964
rect 247966 239912 247972 239964
rect 248276 239912 248282 239964
rect 248334 239912 248340 239964
rect 248460 239912 248466 239964
rect 248518 239952 248524 239964
rect 248518 239924 248644 239952
rect 248518 239912 248524 239924
rect 246436 239844 246442 239896
rect 246494 239844 246500 239896
rect 246454 239760 246482 239844
rect 246390 239708 246396 239760
rect 246448 239720 246482 239760
rect 246448 239708 246454 239720
rect 246298 239640 246304 239692
rect 246356 239640 246362 239692
rect 245442 239584 245476 239624
rect 245344 239572 245350 239584
rect 245470 239572 245476 239584
rect 245528 239572 245534 239624
rect 245378 239544 245384 239556
rect 245028 239516 245384 239544
rect 245120 239352 245148 239516
rect 245378 239504 245384 239516
rect 245436 239504 245442 239556
rect 246482 239504 246488 239556
rect 246540 239544 246546 239556
rect 246638 239544 246666 239912
rect 246540 239516 246666 239544
rect 246540 239504 246546 239516
rect 246390 239436 246396 239488
rect 246448 239476 246454 239488
rect 246730 239476 246758 239912
rect 246448 239448 246758 239476
rect 246448 239436 246454 239448
rect 246942 239368 246948 239420
rect 247000 239408 247006 239420
rect 247374 239408 247402 239912
rect 247632 239844 247638 239896
rect 247690 239844 247696 239896
rect 247650 239680 247678 239844
rect 247512 239652 247678 239680
rect 247512 239556 247540 239652
rect 247742 239556 247770 239912
rect 247494 239504 247500 239556
rect 247552 239504 247558 239556
rect 247678 239504 247684 239556
rect 247736 239516 247770 239556
rect 247834 239556 247862 239912
rect 247926 239760 247954 239912
rect 248000 239844 248006 239896
rect 248058 239844 248064 239896
rect 248092 239844 248098 239896
rect 248150 239844 248156 239896
rect 247908 239708 247914 239760
rect 247966 239708 247972 239760
rect 248018 239624 248046 239844
rect 248110 239692 248138 239844
rect 248294 239692 248322 239912
rect 248616 239692 248644 239924
rect 248828 239912 248834 239964
rect 248886 239912 248892 239964
rect 248846 239816 248874 239912
rect 248938 239896 248966 239992
rect 249196 239912 249202 239964
rect 249254 239952 249260 239964
rect 249254 239912 249288 239952
rect 249380 239912 249386 239964
rect 249438 239952 249444 239964
rect 249438 239912 249472 239952
rect 249932 239912 249938 239964
rect 249990 239912 249996 239964
rect 248920 239844 248926 239896
rect 248978 239844 248984 239896
rect 249012 239844 249018 239896
rect 249070 239884 249076 239896
rect 249070 239856 249196 239884
rect 249070 239844 249076 239856
rect 248846 239788 249104 239816
rect 249076 239760 249104 239788
rect 249058 239708 249064 239760
rect 249116 239708 249122 239760
rect 248110 239652 248144 239692
rect 248138 239640 248144 239652
rect 248196 239640 248202 239692
rect 248294 239652 248328 239692
rect 248322 239640 248328 239652
rect 248380 239640 248386 239692
rect 248598 239640 248604 239692
rect 248656 239640 248662 239692
rect 248874 239640 248880 239692
rect 248932 239640 248938 239692
rect 248966 239640 248972 239692
rect 249024 239680 249030 239692
rect 249168 239680 249196 239856
rect 249024 239652 249196 239680
rect 249024 239640 249030 239652
rect 247954 239572 247960 239624
rect 248012 239584 248046 239624
rect 248892 239612 248920 239640
rect 249260 239612 249288 239912
rect 249334 239640 249340 239692
rect 249392 239640 249398 239692
rect 248892 239584 249288 239612
rect 248012 239572 248018 239584
rect 249352 239556 249380 239640
rect 249444 239612 249472 239912
rect 249564 239844 249570 239896
rect 249622 239844 249628 239896
rect 249656 239844 249662 239896
rect 249714 239884 249720 239896
rect 249714 239844 249748 239884
rect 249840 239844 249846 239896
rect 249898 239844 249904 239896
rect 249582 239748 249610 239844
rect 249582 239720 249656 239748
rect 249444 239584 249518 239612
rect 247834 239516 247868 239556
rect 247736 239504 247742 239516
rect 247862 239504 247868 239516
rect 247920 239504 247926 239556
rect 249334 239504 249340 239556
rect 249392 239504 249398 239556
rect 248690 239436 248696 239488
rect 248748 239476 248754 239488
rect 249490 239476 249518 239584
rect 249628 239544 249656 239720
rect 249720 239612 249748 239844
rect 249858 239816 249886 239844
rect 249812 239788 249886 239816
rect 249812 239760 249840 239788
rect 249950 239760 249978 239912
rect 249794 239708 249800 239760
rect 249852 239708 249858 239760
rect 249886 239708 249892 239760
rect 249944 239720 249978 239760
rect 249944 239708 249950 239720
rect 249720 239584 249840 239612
rect 249702 239544 249708 239556
rect 249628 239516 249708 239544
rect 249702 239504 249708 239516
rect 249760 239504 249766 239556
rect 248748 239448 249518 239476
rect 248748 239436 248754 239448
rect 249610 239436 249616 239488
rect 249668 239476 249674 239488
rect 249812 239476 249840 239584
rect 250502 239556 250530 239992
rect 250576 239912 250582 239964
rect 250634 239912 250640 239964
rect 250668 239912 250674 239964
rect 250726 239952 250732 239964
rect 251146 239952 251174 240196
rect 253676 240020 253704 240196
rect 251514 239992 252186 240020
rect 251514 239964 251542 239992
rect 250726 239924 251174 239952
rect 250726 239912 250732 239924
rect 251220 239912 251226 239964
rect 251278 239912 251284 239964
rect 251312 239912 251318 239964
rect 251370 239912 251376 239964
rect 251404 239912 251410 239964
rect 251462 239912 251468 239964
rect 251496 239912 251502 239964
rect 251554 239912 251560 239964
rect 251680 239912 251686 239964
rect 251738 239912 251744 239964
rect 251772 239912 251778 239964
rect 251830 239912 251836 239964
rect 251864 239912 251870 239964
rect 251922 239952 251928 239964
rect 251922 239912 251956 239952
rect 250594 239748 250622 239912
rect 251036 239844 251042 239896
rect 251094 239844 251100 239896
rect 250714 239748 250720 239760
rect 250594 239720 250720 239748
rect 250714 239708 250720 239720
rect 250772 239708 250778 239760
rect 251054 239624 251082 239844
rect 251238 239680 251266 239912
rect 250990 239572 250996 239624
rect 251048 239584 251082 239624
rect 251192 239652 251266 239680
rect 251048 239572 251054 239584
rect 250502 239516 250536 239556
rect 250530 239504 250536 239516
rect 250588 239504 250594 239556
rect 251192 239488 251220 239652
rect 251330 239624 251358 239912
rect 251266 239572 251272 239624
rect 251324 239584 251358 239624
rect 251324 239572 251330 239584
rect 249668 239448 249840 239476
rect 249668 239436 249674 239448
rect 251174 239436 251180 239488
rect 251232 239436 251238 239488
rect 247000 239380 247402 239408
rect 247000 239368 247006 239380
rect 248782 239368 248788 239420
rect 248840 239408 248846 239420
rect 249058 239408 249064 239420
rect 248840 239380 249064 239408
rect 248840 239368 248846 239380
rect 249058 239368 249064 239380
rect 249116 239368 249122 239420
rect 249242 239368 249248 239420
rect 249300 239408 249306 239420
rect 250162 239408 250168 239420
rect 249300 239380 250168 239408
rect 249300 239368 249306 239380
rect 250162 239368 250168 239380
rect 250220 239368 250226 239420
rect 250806 239368 250812 239420
rect 250864 239408 250870 239420
rect 251422 239408 251450 239912
rect 251698 239884 251726 239912
rect 251652 239856 251726 239884
rect 251542 239708 251548 239760
rect 251600 239748 251606 239760
rect 251652 239748 251680 239856
rect 251790 239828 251818 239912
rect 251726 239776 251732 239828
rect 251784 239788 251818 239828
rect 251784 239776 251790 239788
rect 251818 239748 251824 239760
rect 251600 239720 251824 239748
rect 251600 239708 251606 239720
rect 251818 239708 251824 239720
rect 251876 239708 251882 239760
rect 251928 239624 251956 239912
rect 252048 239884 252054 239896
rect 252020 239844 252054 239884
rect 252106 239844 252112 239896
rect 251910 239572 251916 239624
rect 251968 239572 251974 239624
rect 251634 239504 251640 239556
rect 251692 239544 251698 239556
rect 251818 239544 251824 239556
rect 251692 239516 251824 239544
rect 251692 239504 251698 239516
rect 251818 239504 251824 239516
rect 251876 239504 251882 239556
rect 252020 239488 252048 239844
rect 252002 239436 252008 239488
rect 252060 239436 252066 239488
rect 252158 239476 252186 239992
rect 252894 239992 253612 240020
rect 253676 239992 254716 240020
rect 252894 239964 252922 239992
rect 252232 239912 252238 239964
rect 252290 239952 252296 239964
rect 252290 239924 252600 239952
rect 252290 239912 252296 239924
rect 252416 239844 252422 239896
rect 252474 239844 252480 239896
rect 252434 239760 252462 239844
rect 252370 239708 252376 239760
rect 252428 239720 252462 239760
rect 252428 239708 252434 239720
rect 252572 239556 252600 239924
rect 252692 239912 252698 239964
rect 252750 239912 252756 239964
rect 252876 239912 252882 239964
rect 252934 239912 252940 239964
rect 252968 239912 252974 239964
rect 253026 239912 253032 239964
rect 253244 239912 253250 239964
rect 253302 239912 253308 239964
rect 253584 239952 253612 239992
rect 253888 239952 253894 239964
rect 253584 239924 253796 239952
rect 252710 239884 252738 239912
rect 252710 239856 252876 239884
rect 252848 239692 252876 239856
rect 252830 239640 252836 239692
rect 252888 239640 252894 239692
rect 252738 239572 252744 239624
rect 252796 239612 252802 239624
rect 252986 239612 253014 239912
rect 252796 239584 253014 239612
rect 252796 239572 252802 239584
rect 252554 239504 252560 239556
rect 252612 239504 252618 239556
rect 252922 239476 252928 239488
rect 252158 239448 252928 239476
rect 252922 239436 252928 239448
rect 252980 239436 252986 239488
rect 250864 239380 251450 239408
rect 250864 239368 250870 239380
rect 243320 239312 244228 239340
rect 243320 239300 243326 239312
rect 245102 239300 245108 239352
rect 245160 239300 245166 239352
rect 247034 239300 247040 239352
rect 247092 239340 247098 239352
rect 251542 239340 251548 239352
rect 247092 239312 251548 239340
rect 247092 239300 247098 239312
rect 251542 239300 251548 239312
rect 251600 239300 251606 239352
rect 252554 239300 252560 239352
rect 252612 239340 252618 239352
rect 253262 239340 253290 239912
rect 253520 239844 253526 239896
rect 253578 239844 253584 239896
rect 253612 239844 253618 239896
rect 253670 239844 253676 239896
rect 253538 239760 253566 239844
rect 253630 239816 253658 239844
rect 253630 239788 253704 239816
rect 253538 239720 253572 239760
rect 253566 239708 253572 239720
rect 253624 239708 253630 239760
rect 253382 239572 253388 239624
rect 253440 239612 253446 239624
rect 253676 239612 253704 239788
rect 253440 239584 253704 239612
rect 253440 239572 253446 239584
rect 252612 239312 253290 239340
rect 253768 239340 253796 239924
rect 253860 239912 253894 239952
rect 253946 239912 253952 239964
rect 254256 239912 254262 239964
rect 254314 239912 254320 239964
rect 254532 239952 254538 239964
rect 254412 239924 254538 239952
rect 253860 239556 253888 239912
rect 254164 239844 254170 239896
rect 254222 239844 254228 239896
rect 253842 239504 253848 239556
rect 253900 239504 253906 239556
rect 254182 239476 254210 239844
rect 254274 239544 254302 239912
rect 254412 239760 254440 239924
rect 254532 239912 254538 239924
rect 254590 239912 254596 239964
rect 254394 239708 254400 239760
rect 254452 239708 254458 239760
rect 254688 239692 254716 239992
rect 256896 239964 256924 241012
rect 272242 241000 272248 241012
rect 272300 241000 272306 241052
rect 273438 241000 273444 241052
rect 273496 241040 273502 241052
rect 274450 241040 274456 241052
rect 273496 241012 274456 241040
rect 273496 241000 273502 241012
rect 274450 241000 274456 241012
rect 274508 241000 274514 241052
rect 267550 240932 267556 240984
rect 267608 240972 267614 240984
rect 270678 240972 270684 240984
rect 267608 240944 270684 240972
rect 267608 240932 267614 240944
rect 270678 240932 270684 240944
rect 270736 240932 270742 240984
rect 283006 240932 283012 240984
rect 283064 240972 283070 240984
rect 308398 240972 308404 240984
rect 283064 240944 308404 240972
rect 283064 240932 283070 240944
rect 308398 240932 308404 240944
rect 308456 240932 308462 240984
rect 267458 240864 267464 240916
rect 267516 240904 267522 240916
rect 267734 240904 267740 240916
rect 267516 240876 267740 240904
rect 267516 240864 267522 240876
rect 267734 240864 267740 240876
rect 267792 240864 267798 240916
rect 271598 240904 271604 240916
rect 268948 240876 271604 240904
rect 268838 240836 268844 240848
rect 259564 240808 268844 240836
rect 259564 240496 259592 240808
rect 268838 240796 268844 240808
rect 268896 240796 268902 240848
rect 268948 240768 268976 240876
rect 271598 240864 271604 240876
rect 271656 240864 271662 240916
rect 278130 240864 278136 240916
rect 278188 240904 278194 240916
rect 306098 240904 306104 240916
rect 278188 240876 306104 240904
rect 278188 240864 278194 240876
rect 306098 240864 306104 240876
rect 306156 240864 306162 240916
rect 269482 240836 269488 240848
rect 257770 240468 259592 240496
rect 261450 240740 268976 240768
rect 269040 240808 269488 240836
rect 257770 240020 257798 240468
rect 259702 240060 260788 240088
rect 257770 239992 258074 240020
rect 257770 239964 257798 239992
rect 255176 239952 255182 239964
rect 254918 239924 255182 239952
rect 254670 239640 254676 239692
rect 254728 239640 254734 239692
rect 254274 239516 254440 239544
rect 254302 239476 254308 239488
rect 254182 239448 254308 239476
rect 254302 239436 254308 239448
rect 254360 239436 254366 239488
rect 254026 239368 254032 239420
rect 254084 239408 254090 239420
rect 254412 239408 254440 239516
rect 254084 239380 254440 239408
rect 254084 239368 254090 239380
rect 254918 239352 254946 239924
rect 255176 239912 255182 239924
rect 255234 239912 255240 239964
rect 255452 239912 255458 239964
rect 255510 239912 255516 239964
rect 255820 239952 255826 239964
rect 255792 239912 255826 239952
rect 255878 239912 255884 239964
rect 256372 239912 256378 239964
rect 256430 239912 256436 239964
rect 256648 239912 256654 239964
rect 256706 239912 256712 239964
rect 256740 239912 256746 239964
rect 256798 239912 256804 239964
rect 256832 239912 256838 239964
rect 256890 239924 256924 239964
rect 256890 239912 256896 239924
rect 257108 239912 257114 239964
rect 257166 239912 257172 239964
rect 257476 239912 257482 239964
rect 257534 239912 257540 239964
rect 257752 239912 257758 239964
rect 257810 239912 257816 239964
rect 257936 239952 257942 239964
rect 257908 239912 257942 239952
rect 257994 239912 258000 239964
rect 258046 239952 258074 239992
rect 258414 239992 259638 240020
rect 258414 239964 258442 239992
rect 258046 239924 258212 239952
rect 254992 239844 254998 239896
rect 255050 239844 255056 239896
rect 255010 239612 255038 239844
rect 255130 239776 255136 239828
rect 255188 239776 255194 239828
rect 255148 239680 255176 239776
rect 255470 239748 255498 239912
rect 255636 239844 255642 239896
rect 255694 239884 255700 239896
rect 255694 239844 255728 239884
rect 255470 239720 255636 239748
rect 255608 239692 255636 239720
rect 255700 239692 255728 239844
rect 255148 239652 255544 239680
rect 255314 239612 255320 239624
rect 255010 239584 255320 239612
rect 255314 239572 255320 239584
rect 255372 239572 255378 239624
rect 253842 239340 253848 239352
rect 253768 239312 253848 239340
rect 252612 239300 252618 239312
rect 253842 239300 253848 239312
rect 253900 239300 253906 239352
rect 254918 239312 254952 239352
rect 254946 239300 254952 239312
rect 255004 239300 255010 239352
rect 255516 239340 255544 239652
rect 255590 239640 255596 239692
rect 255648 239640 255654 239692
rect 255682 239640 255688 239692
rect 255740 239640 255746 239692
rect 255792 239544 255820 239912
rect 256004 239844 256010 239896
rect 256062 239844 256068 239896
rect 256022 239760 256050 239844
rect 256022 239720 256056 239760
rect 256050 239708 256056 239720
rect 256108 239708 256114 239760
rect 255958 239640 255964 239692
rect 256016 239680 256022 239692
rect 256390 239680 256418 239912
rect 256666 239828 256694 239912
rect 256758 239884 256786 239912
rect 256758 239856 256832 239884
rect 256804 239828 256832 239856
rect 257016 239844 257022 239896
rect 257074 239844 257080 239896
rect 256666 239788 256700 239828
rect 256694 239776 256700 239788
rect 256752 239776 256758 239828
rect 256786 239776 256792 239828
rect 256844 239776 256850 239828
rect 257034 239680 257062 239844
rect 256016 239652 256418 239680
rect 256804 239652 257062 239680
rect 256016 239640 256022 239652
rect 256234 239544 256240 239556
rect 255792 239516 256240 239544
rect 256234 239504 256240 239516
rect 256292 239504 256298 239556
rect 256804 239488 256832 239652
rect 257126 239624 257154 239912
rect 257384 239844 257390 239896
rect 257442 239844 257448 239896
rect 257402 239692 257430 239844
rect 257494 239748 257522 239912
rect 257908 239760 257936 239912
rect 258028 239884 258034 239896
rect 258000 239844 258034 239884
rect 258086 239844 258092 239896
rect 257494 239720 257660 239748
rect 257632 239692 257660 239720
rect 257890 239708 257896 239760
rect 257948 239708 257954 239760
rect 257402 239652 257436 239692
rect 257430 239640 257436 239652
rect 257488 239640 257494 239692
rect 257614 239640 257620 239692
rect 257672 239640 257678 239692
rect 257062 239572 257068 239624
rect 257120 239584 257154 239624
rect 257120 239572 257126 239584
rect 257246 239572 257252 239624
rect 257304 239612 257310 239624
rect 258000 239612 258028 239844
rect 258184 239624 258212 239924
rect 258396 239912 258402 239964
rect 258454 239912 258460 239964
rect 258764 239912 258770 239964
rect 258822 239912 258828 239964
rect 258856 239912 258862 239964
rect 258914 239912 258920 239964
rect 259132 239912 259138 239964
rect 259190 239912 259196 239964
rect 258304 239844 258310 239896
rect 258362 239884 258368 239896
rect 258580 239884 258586 239896
rect 258362 239844 258396 239884
rect 257304 239584 258028 239612
rect 257304 239572 257310 239584
rect 258166 239572 258172 239624
rect 258224 239572 258230 239624
rect 257706 239504 257712 239556
rect 257764 239544 257770 239556
rect 257982 239544 257988 239556
rect 257764 239516 257988 239544
rect 257764 239504 257770 239516
rect 257982 239504 257988 239516
rect 258040 239504 258046 239556
rect 258368 239488 258396 239844
rect 258552 239844 258586 239884
rect 258638 239844 258644 239896
rect 258672 239844 258678 239896
rect 258730 239844 258736 239896
rect 258552 239692 258580 239844
rect 258690 239816 258718 239844
rect 258644 239788 258718 239816
rect 258534 239640 258540 239692
rect 258592 239640 258598 239692
rect 258644 239612 258672 239788
rect 258782 239760 258810 239912
rect 258718 239708 258724 239760
rect 258776 239720 258810 239760
rect 258776 239708 258782 239720
rect 258718 239612 258724 239624
rect 258644 239584 258724 239612
rect 258718 239572 258724 239584
rect 258776 239572 258782 239624
rect 258874 239612 258902 239912
rect 259040 239844 259046 239896
rect 259098 239844 259104 239896
rect 259058 239760 259086 239844
rect 258994 239708 259000 239760
rect 259052 239720 259086 239760
rect 259052 239708 259058 239720
rect 259150 239680 259178 239912
rect 259408 239884 259414 239896
rect 259380 239844 259414 239884
rect 259466 239844 259472 239896
rect 259500 239844 259506 239896
rect 259558 239844 259564 239896
rect 259610 239884 259638 239992
rect 259702 239964 259730 240060
rect 259886 239992 260282 240020
rect 259886 239964 259914 239992
rect 259684 239912 259690 239964
rect 259742 239912 259748 239964
rect 259868 239912 259874 239964
rect 259926 239912 259932 239964
rect 259960 239912 259966 239964
rect 260018 239912 260024 239964
rect 260144 239912 260150 239964
rect 260202 239912 260208 239964
rect 259610 239856 259684 239884
rect 259380 239748 259408 239844
rect 259518 239816 259546 239844
rect 259518 239788 259592 239816
rect 259454 239748 259460 239760
rect 259380 239720 259460 239748
rect 259454 239708 259460 239720
rect 259512 239708 259518 239760
rect 259150 239652 259408 239680
rect 259380 239624 259408 239652
rect 259564 239624 259592 239788
rect 259086 239612 259092 239624
rect 258874 239584 259092 239612
rect 259086 239572 259092 239584
rect 259144 239572 259150 239624
rect 259362 239572 259368 239624
rect 259420 239572 259426 239624
rect 259546 239572 259552 239624
rect 259604 239572 259610 239624
rect 256786 239436 256792 239488
rect 256844 239436 256850 239488
rect 258350 239436 258356 239488
rect 258408 239436 258414 239488
rect 259656 239476 259684 239856
rect 259978 239816 260006 239912
rect 259840 239788 260006 239816
rect 259840 239544 259868 239788
rect 260162 239748 260190 239912
rect 259932 239720 260190 239748
rect 259932 239612 259960 239720
rect 260006 239640 260012 239692
rect 260064 239680 260070 239692
rect 260254 239680 260282 239992
rect 260420 239912 260426 239964
rect 260478 239912 260484 239964
rect 260438 239760 260466 239912
rect 260604 239844 260610 239896
rect 260662 239844 260668 239896
rect 260438 239720 260472 239760
rect 260466 239708 260472 239720
rect 260524 239708 260530 239760
rect 260064 239652 260282 239680
rect 260622 239680 260650 239844
rect 260622 239652 260696 239680
rect 260064 239640 260070 239652
rect 260668 239624 260696 239652
rect 259932 239584 260512 239612
rect 260006 239544 260012 239556
rect 259840 239516 260012 239544
rect 260006 239504 260012 239516
rect 260064 239504 260070 239556
rect 260282 239476 260288 239488
rect 258460 239448 260288 239476
rect 258460 239420 258488 239448
rect 260282 239436 260288 239448
rect 260340 239436 260346 239488
rect 258442 239368 258448 239420
rect 258500 239368 258506 239420
rect 259638 239368 259644 239420
rect 259696 239408 259702 239420
rect 260484 239408 260512 239584
rect 260650 239572 260656 239624
rect 260708 239572 260714 239624
rect 260760 239544 260788 240060
rect 260880 239912 260886 239964
rect 260938 239912 260944 239964
rect 261156 239912 261162 239964
rect 261214 239912 261220 239964
rect 261248 239912 261254 239964
rect 261306 239952 261312 239964
rect 261450 239952 261478 240740
rect 269040 240700 269068 240808
rect 269482 240796 269488 240808
rect 269540 240796 269546 240848
rect 271138 240796 271144 240848
rect 271196 240836 271202 240848
rect 287698 240836 287704 240848
rect 271196 240808 287704 240836
rect 271196 240796 271202 240808
rect 287698 240796 287704 240808
rect 287756 240796 287762 240848
rect 287974 240796 287980 240848
rect 288032 240836 288038 240848
rect 312538 240836 312544 240848
rect 288032 240808 312544 240836
rect 288032 240796 288038 240808
rect 312538 240796 312544 240808
rect 312596 240796 312602 240848
rect 269206 240728 269212 240780
rect 269264 240768 269270 240780
rect 299198 240768 299204 240780
rect 269264 240740 299204 240768
rect 269264 240728 269270 240740
rect 299198 240728 299204 240740
rect 299256 240728 299262 240780
rect 261306 239924 261478 239952
rect 261542 240672 269068 240700
rect 261306 239912 261312 239924
rect 260898 239612 260926 239912
rect 261018 239640 261024 239692
rect 261076 239680 261082 239692
rect 261174 239680 261202 239912
rect 261076 239652 261202 239680
rect 261076 239640 261082 239652
rect 261294 239612 261300 239624
rect 260898 239584 261300 239612
rect 261294 239572 261300 239584
rect 261352 239572 261358 239624
rect 261542 239544 261570 240672
rect 269114 240660 269120 240712
rect 269172 240700 269178 240712
rect 274726 240700 274732 240712
rect 269172 240672 274732 240700
rect 269172 240660 269178 240672
rect 274726 240660 274732 240672
rect 274784 240660 274790 240712
rect 269574 240632 269580 240644
rect 262002 240604 269580 240632
rect 262002 239964 262030 240604
rect 269574 240592 269580 240604
rect 269632 240592 269638 240644
rect 267918 240564 267924 240576
rect 266234 240536 267924 240564
rect 266234 240496 266262 240536
rect 267918 240524 267924 240536
rect 267976 240524 267982 240576
rect 269206 240524 269212 240576
rect 269264 240564 269270 240576
rect 278774 240564 278780 240576
rect 269264 240536 278780 240564
rect 269264 240524 269270 240536
rect 278774 240524 278780 240536
rect 278832 240564 278838 240576
rect 278958 240564 278964 240576
rect 278832 240536 278964 240564
rect 278832 240524 278838 240536
rect 278958 240524 278964 240536
rect 279016 240524 279022 240576
rect 262830 240468 266262 240496
rect 261800 239912 261806 239964
rect 261858 239952 261864 239964
rect 261858 239912 261892 239952
rect 261984 239912 261990 239964
rect 262042 239912 262048 239964
rect 262168 239912 262174 239964
rect 262226 239952 262232 239964
rect 262226 239924 262490 239952
rect 262226 239912 262232 239924
rect 261616 239844 261622 239896
rect 261674 239884 261680 239896
rect 261674 239844 261708 239884
rect 261680 239624 261708 239844
rect 261864 239692 261892 239912
rect 262352 239844 262358 239896
rect 262410 239844 262416 239896
rect 262370 239760 262398 239844
rect 262306 239708 262312 239760
rect 262364 239720 262398 239760
rect 262364 239708 262370 239720
rect 261846 239640 261852 239692
rect 261904 239640 261910 239692
rect 261662 239572 261668 239624
rect 261720 239572 261726 239624
rect 262462 239556 262490 239924
rect 262720 239912 262726 239964
rect 262778 239952 262784 239964
rect 262830 239952 262858 240468
rect 270126 240456 270132 240508
rect 270184 240496 270190 240508
rect 287790 240496 287796 240508
rect 270184 240468 287796 240496
rect 270184 240456 270190 240468
rect 287790 240456 287796 240468
rect 287848 240496 287854 240508
rect 287974 240496 287980 240508
rect 287848 240468 287980 240496
rect 287848 240456 287854 240468
rect 287974 240456 287980 240468
rect 288032 240456 288038 240508
rect 268286 240428 268292 240440
rect 262922 240400 268292 240428
rect 262922 239964 262950 240400
rect 268286 240388 268292 240400
rect 268344 240388 268350 240440
rect 268194 240360 268200 240372
rect 264532 240332 268200 240360
rect 264532 240020 264560 240332
rect 268194 240320 268200 240332
rect 268252 240320 268258 240372
rect 268838 240320 268844 240372
rect 268896 240360 268902 240372
rect 283006 240360 283012 240372
rect 268896 240332 283012 240360
rect 268896 240320 268902 240332
rect 283006 240320 283012 240332
rect 283064 240320 283070 240372
rect 263014 239992 263640 240020
rect 263014 239964 263042 239992
rect 262778 239924 262858 239952
rect 262778 239912 262784 239924
rect 262904 239912 262910 239964
rect 262962 239912 262968 239964
rect 262996 239912 263002 239964
rect 263054 239912 263060 239964
rect 263088 239912 263094 239964
rect 263146 239912 263152 239964
rect 263272 239952 263278 239964
rect 263244 239912 263278 239952
rect 263330 239912 263336 239964
rect 263456 239912 263462 239964
rect 263514 239912 263520 239964
rect 262536 239844 262542 239896
rect 262594 239844 262600 239896
rect 262922 239884 262950 239912
rect 262922 239856 262996 239884
rect 262554 239612 262582 239844
rect 262968 239828 262996 239856
rect 263106 239828 263134 239912
rect 262950 239776 262956 239828
rect 263008 239776 263014 239828
rect 263042 239776 263048 239828
rect 263100 239788 263134 239828
rect 263100 239776 263106 239788
rect 263244 239748 263272 239912
rect 263474 239760 263502 239912
rect 263152 239720 263272 239748
rect 263152 239692 263180 239720
rect 263410 239708 263416 239760
rect 263468 239720 263502 239760
rect 263468 239708 263474 239720
rect 263612 239692 263640 239992
rect 264026 239992 264560 240020
rect 264026 239964 264054 239992
rect 263732 239912 263738 239964
rect 263790 239912 263796 239964
rect 264008 239912 264014 239964
rect 264066 239912 264072 239964
rect 264376 239952 264382 239964
rect 264164 239924 264382 239952
rect 263750 239692 263778 239912
rect 263824 239844 263830 239896
rect 263882 239844 263888 239896
rect 263842 239760 263870 239844
rect 263842 239720 263876 239760
rect 263870 239708 263876 239720
rect 263928 239708 263934 239760
rect 263134 239640 263140 239692
rect 263192 239640 263198 239692
rect 263594 239640 263600 239692
rect 263652 239640 263658 239692
rect 263750 239652 263784 239692
rect 263778 239640 263784 239652
rect 263836 239640 263842 239692
rect 264164 239624 264192 239924
rect 264376 239912 264382 239924
rect 264434 239912 264440 239964
rect 264532 239624 264560 239992
rect 265590 240264 267872 240292
rect 265590 239964 265618 240264
rect 267844 240224 267872 240264
rect 267918 240252 267924 240304
rect 267976 240292 267982 240304
rect 288434 240292 288440 240304
rect 267976 240264 288440 240292
rect 267976 240252 267982 240264
rect 288434 240252 288440 240264
rect 288492 240252 288498 240304
rect 270126 240224 270132 240236
rect 267844 240196 270132 240224
rect 270126 240184 270132 240196
rect 270184 240184 270190 240236
rect 270678 240184 270684 240236
rect 270736 240224 270742 240236
rect 278130 240224 278136 240236
rect 270736 240196 278136 240224
rect 270736 240184 270742 240196
rect 278130 240184 278136 240196
rect 278188 240184 278194 240236
rect 269482 240156 269488 240168
rect 266740 240128 269488 240156
rect 266740 240020 266768 240128
rect 269482 240116 269488 240128
rect 269540 240116 269546 240168
rect 267550 240048 267556 240100
rect 267608 240088 267614 240100
rect 268194 240088 268200 240100
rect 267608 240060 268200 240088
rect 267608 240048 267614 240060
rect 268194 240048 268200 240060
rect 268252 240048 268258 240100
rect 285766 240048 285772 240100
rect 285824 240088 285830 240100
rect 286778 240088 286784 240100
rect 285824 240060 286784 240088
rect 285824 240048 285830 240060
rect 286778 240048 286784 240060
rect 286836 240048 286842 240100
rect 265682 239992 266768 240020
rect 265682 239964 265710 239992
rect 264836 239952 264842 239964
rect 264808 239912 264842 239952
rect 264894 239912 264900 239964
rect 264928 239912 264934 239964
rect 264986 239952 264992 239964
rect 264986 239912 265020 239952
rect 265572 239912 265578 239964
rect 265630 239912 265636 239964
rect 265664 239912 265670 239964
rect 265722 239912 265728 239964
rect 266768 239912 266774 239964
rect 266826 239952 266832 239964
rect 266826 239924 266998 239952
rect 266826 239912 266832 239924
rect 264808 239692 264836 239912
rect 264790 239640 264796 239692
rect 264848 239640 264854 239692
rect 264054 239612 264060 239624
rect 262554 239584 264060 239612
rect 264054 239572 264060 239584
rect 264112 239572 264118 239624
rect 264146 239572 264152 239624
rect 264204 239572 264210 239624
rect 264514 239572 264520 239624
rect 264572 239572 264578 239624
rect 264992 239612 265020 239912
rect 265112 239844 265118 239896
rect 265170 239844 265176 239896
rect 265480 239844 265486 239896
rect 265538 239884 265544 239896
rect 265538 239856 265756 239884
rect 265538 239844 265544 239856
rect 265130 239816 265158 239844
rect 265618 239816 265624 239828
rect 265130 239788 265624 239816
rect 265618 239776 265624 239788
rect 265676 239776 265682 239828
rect 265526 239708 265532 239760
rect 265584 239748 265590 239760
rect 265728 239748 265756 239856
rect 266032 239844 266038 239896
rect 266090 239844 266096 239896
rect 266216 239844 266222 239896
rect 266274 239884 266280 239896
rect 266274 239856 266768 239884
rect 266274 239844 266280 239856
rect 265584 239720 265756 239748
rect 265584 239708 265590 239720
rect 265434 239640 265440 239692
rect 265492 239680 265498 239692
rect 266050 239680 266078 239844
rect 265492 239652 266078 239680
rect 265492 239640 265498 239652
rect 265894 239612 265900 239624
rect 264992 239584 265900 239612
rect 265894 239572 265900 239584
rect 265952 239572 265958 239624
rect 262122 239544 262128 239556
rect 260760 239516 261340 239544
rect 261542 239516 262128 239544
rect 261018 239436 261024 239488
rect 261076 239476 261082 239488
rect 261202 239476 261208 239488
rect 261076 239448 261208 239476
rect 261076 239436 261082 239448
rect 261202 239436 261208 239448
rect 261260 239436 261266 239488
rect 261312 239476 261340 239516
rect 262122 239504 262128 239516
rect 262180 239504 262186 239556
rect 262462 239516 262496 239556
rect 262490 239504 262496 239516
rect 262548 239544 262554 239556
rect 266740 239544 266768 239856
rect 266970 239680 266998 239924
rect 267044 239912 267050 239964
rect 267102 239912 267108 239964
rect 267228 239912 267234 239964
rect 267286 239952 267292 239964
rect 268102 239952 268108 239964
rect 267286 239924 268108 239952
rect 267286 239912 267292 239924
rect 268102 239912 268108 239924
rect 268160 239912 268166 239964
rect 267062 239760 267090 239912
rect 267734 239776 267740 239828
rect 267792 239816 267798 239828
rect 299106 239816 299112 239828
rect 267792 239788 299112 239816
rect 267792 239776 267798 239788
rect 299106 239776 299112 239788
rect 299164 239776 299170 239828
rect 267062 239720 267096 239760
rect 267090 239708 267096 239720
rect 267148 239708 267154 239760
rect 267182 239708 267188 239760
rect 267240 239748 267246 239760
rect 268470 239748 268476 239760
rect 267240 239720 268476 239748
rect 267240 239708 267246 239720
rect 268470 239708 268476 239720
rect 268528 239708 268534 239760
rect 271230 239708 271236 239760
rect 271288 239748 271294 239760
rect 293586 239748 293592 239760
rect 271288 239720 293592 239748
rect 271288 239708 271294 239720
rect 293586 239708 293592 239720
rect 293644 239708 293650 239760
rect 268010 239680 268016 239692
rect 266970 239652 268016 239680
rect 268010 239640 268016 239652
rect 268068 239640 268074 239692
rect 278682 239680 278688 239692
rect 271248 239652 278688 239680
rect 266952 239572 266958 239624
rect 267010 239612 267016 239624
rect 270862 239612 270868 239624
rect 267010 239584 270868 239612
rect 267010 239572 267016 239584
rect 270862 239572 270868 239584
rect 270920 239572 270926 239624
rect 269206 239544 269212 239556
rect 262548 239516 266676 239544
rect 266740 239516 269212 239544
rect 262548 239504 262554 239516
rect 262582 239476 262588 239488
rect 261312 239448 262588 239476
rect 262582 239436 262588 239448
rect 262640 239436 262646 239488
rect 266648 239476 266676 239516
rect 269206 239504 269212 239516
rect 269264 239504 269270 239556
rect 267182 239476 267188 239488
rect 263612 239448 266584 239476
rect 266648 239448 267188 239476
rect 263612 239420 263640 239448
rect 259696 239380 260512 239408
rect 259696 239368 259702 239380
rect 263134 239368 263140 239420
rect 263192 239408 263198 239420
rect 263594 239408 263600 239420
rect 263192 239380 263600 239408
rect 263192 239368 263198 239380
rect 263594 239368 263600 239380
rect 263652 239368 263658 239420
rect 264698 239368 264704 239420
rect 264756 239408 264762 239420
rect 265894 239408 265900 239420
rect 264756 239380 265900 239408
rect 264756 239368 264762 239380
rect 265894 239368 265900 239380
rect 265952 239368 265958 239420
rect 259730 239340 259736 239352
rect 255516 239312 259736 239340
rect 259730 239300 259736 239312
rect 259788 239300 259794 239352
rect 260282 239300 260288 239352
rect 260340 239340 260346 239352
rect 264882 239340 264888 239352
rect 260340 239312 264888 239340
rect 260340 239300 260346 239312
rect 264882 239300 264888 239312
rect 264940 239300 264946 239352
rect 266556 239340 266584 239448
rect 267182 239436 267188 239448
rect 267240 239436 267246 239488
rect 267274 239436 267280 239488
rect 267332 239476 267338 239488
rect 267734 239476 267740 239488
rect 267332 239448 267740 239476
rect 267332 239436 267338 239448
rect 267734 239436 267740 239448
rect 267792 239476 267798 239488
rect 268746 239476 268752 239488
rect 267792 239448 268752 239476
rect 267792 239436 267798 239448
rect 268746 239436 268752 239448
rect 268804 239436 268810 239488
rect 266630 239368 266636 239420
rect 266688 239408 266694 239420
rect 267550 239408 267556 239420
rect 266688 239380 267556 239408
rect 266688 239368 266694 239380
rect 267550 239368 267556 239380
rect 267608 239368 267614 239420
rect 269482 239368 269488 239420
rect 269540 239408 269546 239420
rect 271248 239408 271276 239652
rect 278682 239640 278688 239652
rect 278740 239640 278746 239692
rect 271506 239572 271512 239624
rect 271564 239612 271570 239624
rect 297818 239612 297824 239624
rect 271564 239584 297824 239612
rect 271564 239572 271570 239584
rect 297818 239572 297824 239584
rect 297876 239572 297882 239624
rect 273254 239504 273260 239556
rect 273312 239544 273318 239556
rect 311250 239544 311256 239556
rect 273312 239516 311256 239544
rect 273312 239504 273318 239516
rect 311250 239504 311256 239516
rect 311308 239504 311314 239556
rect 271598 239436 271604 239488
rect 271656 239476 271662 239488
rect 320818 239476 320824 239488
rect 271656 239448 320824 239476
rect 271656 239436 271662 239448
rect 320818 239436 320824 239448
rect 320876 239436 320882 239488
rect 269540 239380 271276 239408
rect 269540 239368 269546 239380
rect 274266 239368 274272 239420
rect 274324 239408 274330 239420
rect 293862 239408 293868 239420
rect 274324 239380 293868 239408
rect 274324 239368 274330 239380
rect 293862 239368 293868 239380
rect 293920 239408 293926 239420
rect 527174 239408 527180 239420
rect 293920 239380 527180 239408
rect 293920 239368 293926 239380
rect 527174 239368 527180 239380
rect 527232 239368 527238 239420
rect 269942 239340 269948 239352
rect 266556 239312 269948 239340
rect 269942 239300 269948 239312
rect 270000 239300 270006 239352
rect 270678 239300 270684 239352
rect 270736 239340 270742 239352
rect 285766 239340 285772 239352
rect 270736 239312 285772 239340
rect 270736 239300 270742 239312
rect 285766 239300 285772 239312
rect 285824 239300 285830 239352
rect 219032 239244 240548 239272
rect 219032 239232 219038 239244
rect 241422 239232 241428 239284
rect 241480 239272 241486 239284
rect 269390 239272 269396 239284
rect 241480 239244 269396 239272
rect 241480 239232 241486 239244
rect 269390 239232 269396 239244
rect 269448 239232 269454 239284
rect 214742 239164 214748 239216
rect 214800 239204 214806 239216
rect 221090 239204 221096 239216
rect 214800 239176 221096 239204
rect 214800 239164 214806 239176
rect 221090 239164 221096 239176
rect 221148 239204 221154 239216
rect 223390 239204 223396 239216
rect 221148 239176 223396 239204
rect 221148 239164 221154 239176
rect 223390 239164 223396 239176
rect 223448 239164 223454 239216
rect 223482 239164 223488 239216
rect 223540 239204 223546 239216
rect 223850 239204 223856 239216
rect 223540 239176 223856 239204
rect 223540 239164 223546 239176
rect 223850 239164 223856 239176
rect 223908 239164 223914 239216
rect 224954 239164 224960 239216
rect 225012 239204 225018 239216
rect 225690 239204 225696 239216
rect 225012 239176 225696 239204
rect 225012 239164 225018 239176
rect 225690 239164 225696 239176
rect 225748 239164 225754 239216
rect 227898 239164 227904 239216
rect 227956 239204 227962 239216
rect 228174 239204 228180 239216
rect 227956 239176 228180 239204
rect 227956 239164 227962 239176
rect 228174 239164 228180 239176
rect 228232 239164 228238 239216
rect 233418 239164 233424 239216
rect 233476 239204 233482 239216
rect 241146 239204 241152 239216
rect 233476 239176 241152 239204
rect 233476 239164 233482 239176
rect 241146 239164 241152 239176
rect 241204 239164 241210 239216
rect 245654 239164 245660 239216
rect 245712 239204 245718 239216
rect 270034 239204 270040 239216
rect 245712 239176 270040 239204
rect 245712 239164 245718 239176
rect 270034 239164 270040 239176
rect 270092 239164 270098 239216
rect 215754 239096 215760 239148
rect 215812 239136 215818 239148
rect 225966 239136 225972 239148
rect 215812 239108 225972 239136
rect 215812 239096 215818 239108
rect 225966 239096 225972 239108
rect 226024 239096 226030 239148
rect 236178 239136 236184 239148
rect 229020 239108 236184 239136
rect 221182 239028 221188 239080
rect 221240 239068 221246 239080
rect 223114 239068 223120 239080
rect 221240 239040 223120 239068
rect 221240 239028 221246 239040
rect 223114 239028 223120 239040
rect 223172 239028 223178 239080
rect 228082 239028 228088 239080
rect 228140 239068 228146 239080
rect 228818 239068 228824 239080
rect 228140 239040 228824 239068
rect 228140 239028 228146 239040
rect 228818 239028 228824 239040
rect 228876 239028 228882 239080
rect 211982 238960 211988 239012
rect 212040 239000 212046 239012
rect 212258 239000 212264 239012
rect 212040 238972 212264 239000
rect 212040 238960 212046 238972
rect 212258 238960 212264 238972
rect 212316 238960 212322 239012
rect 213270 238960 213276 239012
rect 213328 239000 213334 239012
rect 229020 239000 229048 239108
rect 236178 239096 236184 239108
rect 236236 239136 236242 239148
rect 236914 239136 236920 239148
rect 236236 239108 236920 239136
rect 236236 239096 236242 239108
rect 236914 239096 236920 239108
rect 236972 239096 236978 239148
rect 237834 239096 237840 239148
rect 237892 239136 237898 239148
rect 238110 239136 238116 239148
rect 237892 239108 238116 239136
rect 237892 239096 237898 239108
rect 238110 239096 238116 239108
rect 238168 239096 238174 239148
rect 238570 239096 238576 239148
rect 238628 239136 238634 239148
rect 238628 239108 240732 239136
rect 238628 239096 238634 239108
rect 229830 239028 229836 239080
rect 229888 239068 229894 239080
rect 240704 239068 240732 239108
rect 242250 239096 242256 239148
rect 242308 239136 242314 239148
rect 242526 239136 242532 239148
rect 242308 239108 242532 239136
rect 242308 239096 242314 239108
rect 242526 239096 242532 239108
rect 242584 239096 242590 239148
rect 246298 239136 246304 239148
rect 242636 239108 246304 239136
rect 242636 239068 242664 239108
rect 246298 239096 246304 239108
rect 246356 239096 246362 239148
rect 247770 239096 247776 239148
rect 247828 239136 247834 239148
rect 269850 239136 269856 239148
rect 247828 239108 269856 239136
rect 247828 239096 247834 239108
rect 269850 239096 269856 239108
rect 269908 239096 269914 239148
rect 229888 239040 240640 239068
rect 240704 239040 242664 239068
rect 229888 239028 229894 239040
rect 213328 238972 229048 239000
rect 213328 238960 213334 238972
rect 229462 238960 229468 239012
rect 229520 239000 229526 239012
rect 229520 238972 239812 239000
rect 229520 238960 229526 238972
rect 154298 238892 154304 238944
rect 154356 238932 154362 238944
rect 223758 238932 223764 238944
rect 154356 238904 223764 238932
rect 154356 238892 154362 238904
rect 223758 238892 223764 238904
rect 223816 238892 223822 238944
rect 223850 238892 223856 238944
rect 223908 238932 223914 238944
rect 227714 238932 227720 238944
rect 223908 238904 227720 238932
rect 223908 238892 223914 238904
rect 227714 238892 227720 238904
rect 227772 238892 227778 238944
rect 227990 238892 227996 238944
rect 228048 238932 228054 238944
rect 229480 238932 229508 238960
rect 228048 238904 229508 238932
rect 228048 238892 228054 238904
rect 231118 238892 231124 238944
rect 231176 238932 231182 238944
rect 231578 238932 231584 238944
rect 231176 238904 231584 238932
rect 231176 238892 231182 238904
rect 231578 238892 231584 238904
rect 231636 238892 231642 238944
rect 235534 238892 235540 238944
rect 235592 238932 235598 238944
rect 235592 238904 239720 238932
rect 235592 238892 235598 238904
rect 215938 238824 215944 238876
rect 215996 238864 216002 238876
rect 238478 238864 238484 238876
rect 215996 238836 238484 238864
rect 215996 238824 216002 238836
rect 238478 238824 238484 238836
rect 238536 238824 238542 238876
rect 151538 238756 151544 238808
rect 151596 238796 151602 238808
rect 221274 238796 221280 238808
rect 151596 238768 221280 238796
rect 151596 238756 151602 238768
rect 221274 238756 221280 238768
rect 221332 238756 221338 238808
rect 221458 238756 221464 238808
rect 221516 238796 221522 238808
rect 223850 238796 223856 238808
rect 221516 238768 223856 238796
rect 221516 238756 221522 238768
rect 223850 238756 223856 238768
rect 223908 238756 223914 238808
rect 232314 238796 232320 238808
rect 225708 238768 232320 238796
rect 218974 238688 218980 238740
rect 219032 238728 219038 238740
rect 219434 238728 219440 238740
rect 219032 238700 219440 238728
rect 219032 238688 219038 238700
rect 219434 238688 219440 238700
rect 219492 238688 219498 238740
rect 191650 238620 191656 238672
rect 191708 238660 191714 238672
rect 222378 238660 222384 238672
rect 191708 238632 222384 238660
rect 191708 238620 191714 238632
rect 222378 238620 222384 238632
rect 222436 238620 222442 238672
rect 223114 238620 223120 238672
rect 223172 238660 223178 238672
rect 225708 238660 225736 238768
rect 232314 238756 232320 238768
rect 232372 238756 232378 238808
rect 232406 238756 232412 238808
rect 232464 238796 232470 238808
rect 239030 238796 239036 238808
rect 232464 238768 239036 238796
rect 232464 238756 232470 238768
rect 239030 238756 239036 238768
rect 239088 238756 239094 238808
rect 226426 238688 226432 238740
rect 226484 238728 226490 238740
rect 235534 238728 235540 238740
rect 226484 238700 235540 238728
rect 226484 238688 226490 238700
rect 235534 238688 235540 238700
rect 235592 238688 235598 238740
rect 235994 238688 236000 238740
rect 236052 238728 236058 238740
rect 236052 238700 236500 238728
rect 236052 238688 236058 238700
rect 223172 238632 225736 238660
rect 223172 238620 223178 238632
rect 225966 238620 225972 238672
rect 226024 238660 226030 238672
rect 233510 238660 233516 238672
rect 226024 238632 233516 238660
rect 226024 238620 226030 238632
rect 233510 238620 233516 238632
rect 233568 238620 233574 238672
rect 233786 238620 233792 238672
rect 233844 238660 233850 238672
rect 234430 238660 234436 238672
rect 233844 238632 234436 238660
rect 233844 238620 233850 238632
rect 234430 238620 234436 238632
rect 234488 238620 234494 238672
rect 234614 238620 234620 238672
rect 234672 238660 234678 238672
rect 236362 238660 236368 238672
rect 234672 238632 236368 238660
rect 234672 238620 234678 238632
rect 236362 238620 236368 238632
rect 236420 238620 236426 238672
rect 236472 238660 236500 238700
rect 237834 238688 237840 238740
rect 237892 238728 237898 238740
rect 238018 238728 238024 238740
rect 237892 238700 238024 238728
rect 237892 238688 237898 238700
rect 238018 238688 238024 238700
rect 238076 238728 238082 238740
rect 239692 238728 239720 238904
rect 239784 238796 239812 238972
rect 240612 238864 240640 239040
rect 242894 239028 242900 239080
rect 242952 239068 242958 239080
rect 297634 239068 297640 239080
rect 242952 239040 297640 239068
rect 242952 239028 242958 239040
rect 297634 239028 297640 239040
rect 297692 239028 297698 239080
rect 242526 238960 242532 239012
rect 242584 239000 242590 239012
rect 297542 239000 297548 239012
rect 242584 238972 297548 239000
rect 242584 238960 242590 238972
rect 297542 238960 297548 238972
rect 297600 238960 297606 239012
rect 241146 238892 241152 238944
rect 241204 238932 241210 238944
rect 289354 238932 289360 238944
rect 241204 238904 289360 238932
rect 241204 238892 241210 238904
rect 289354 238892 289360 238904
rect 289412 238892 289418 238944
rect 247770 238864 247776 238876
rect 240612 238836 247776 238864
rect 247770 238824 247776 238836
rect 247828 238824 247834 238876
rect 250162 238824 250168 238876
rect 250220 238864 250226 238876
rect 255130 238864 255136 238876
rect 250220 238836 255136 238864
rect 250220 238824 250226 238836
rect 255130 238824 255136 238836
rect 255188 238824 255194 238876
rect 255682 238824 255688 238876
rect 255740 238864 255746 238876
rect 255958 238864 255964 238876
rect 255740 238836 255964 238864
rect 255740 238824 255746 238836
rect 255958 238824 255964 238836
rect 256016 238824 256022 238876
rect 257522 238824 257528 238876
rect 257580 238864 257586 238876
rect 258074 238864 258080 238876
rect 257580 238836 258080 238864
rect 257580 238824 257586 238836
rect 258074 238824 258080 238836
rect 258132 238824 258138 238876
rect 261110 238824 261116 238876
rect 261168 238864 261174 238876
rect 261386 238864 261392 238876
rect 261168 238836 261392 238864
rect 261168 238824 261174 238836
rect 261386 238824 261392 238836
rect 261444 238824 261450 238876
rect 273254 238864 273260 238876
rect 261496 238836 273260 238864
rect 246850 238796 246856 238808
rect 239784 238768 246856 238796
rect 246850 238756 246856 238768
rect 246908 238756 246914 238808
rect 248966 238756 248972 238808
rect 249024 238796 249030 238808
rect 249150 238796 249156 238808
rect 249024 238768 249156 238796
rect 249024 238756 249030 238768
rect 249150 238756 249156 238768
rect 249208 238756 249214 238808
rect 260558 238796 260564 238808
rect 250364 238768 260564 238796
rect 241422 238728 241428 238740
rect 238076 238700 239352 238728
rect 239692 238700 241428 238728
rect 238076 238688 238082 238700
rect 239324 238660 239352 238700
rect 241422 238688 241428 238700
rect 241480 238688 241486 238740
rect 242894 238660 242900 238672
rect 236472 238632 239260 238660
rect 239324 238632 242900 238660
rect 207658 238552 207664 238604
rect 207716 238592 207722 238604
rect 232130 238592 232136 238604
rect 207716 238564 232136 238592
rect 207716 238552 207722 238564
rect 232130 238552 232136 238564
rect 232188 238552 232194 238604
rect 232314 238552 232320 238604
rect 232372 238592 232378 238604
rect 235258 238592 235264 238604
rect 232372 238564 235264 238592
rect 232372 238552 232378 238564
rect 235258 238552 235264 238564
rect 235316 238552 235322 238604
rect 235534 238552 235540 238604
rect 235592 238592 235598 238604
rect 238846 238592 238852 238604
rect 235592 238564 238852 238592
rect 235592 238552 235598 238564
rect 238846 238552 238852 238564
rect 238904 238552 238910 238604
rect 239232 238592 239260 238632
rect 242894 238620 242900 238632
rect 242952 238620 242958 238672
rect 250364 238660 250392 238768
rect 260558 238756 260564 238768
rect 260616 238756 260622 238808
rect 261496 238796 261524 238836
rect 273254 238824 273260 238836
rect 273312 238824 273318 238876
rect 261220 238768 261524 238796
rect 251726 238688 251732 238740
rect 251784 238728 251790 238740
rect 256510 238728 256516 238740
rect 251784 238700 256516 238728
rect 251784 238688 251790 238700
rect 256510 238688 256516 238700
rect 256568 238688 256574 238740
rect 258166 238688 258172 238740
rect 258224 238728 258230 238740
rect 258810 238728 258816 238740
rect 258224 238700 258816 238728
rect 258224 238688 258230 238700
rect 258810 238688 258816 238700
rect 258868 238688 258874 238740
rect 243096 238632 250392 238660
rect 243096 238592 243124 238632
rect 252922 238620 252928 238672
rect 252980 238660 252986 238672
rect 261220 238660 261248 238768
rect 261570 238756 261576 238808
rect 261628 238796 261634 238808
rect 266354 238796 266360 238808
rect 261628 238768 266360 238796
rect 261628 238756 261634 238768
rect 266354 238756 266360 238768
rect 266412 238756 266418 238808
rect 266538 238756 266544 238808
rect 266596 238796 266602 238808
rect 267826 238796 267832 238808
rect 266596 238768 267832 238796
rect 266596 238756 266602 238768
rect 267826 238756 267832 238768
rect 267884 238756 267890 238808
rect 295242 238756 295248 238808
rect 295300 238796 295306 238808
rect 488534 238796 488540 238808
rect 295300 238768 488540 238796
rect 295300 238756 295306 238768
rect 488534 238756 488540 238768
rect 488592 238756 488598 238808
rect 261294 238688 261300 238740
rect 261352 238728 261358 238740
rect 262674 238728 262680 238740
rect 261352 238700 262680 238728
rect 261352 238688 261358 238700
rect 262674 238688 262680 238700
rect 262732 238688 262738 238740
rect 263686 238688 263692 238740
rect 263744 238728 263750 238740
rect 266630 238728 266636 238740
rect 263744 238700 266636 238728
rect 263744 238688 263750 238700
rect 266630 238688 266636 238700
rect 266688 238688 266694 238740
rect 267274 238688 267280 238740
rect 267332 238728 267338 238740
rect 271506 238728 271512 238740
rect 267332 238700 271512 238728
rect 267332 238688 267338 238700
rect 271506 238688 271512 238700
rect 271564 238688 271570 238740
rect 270678 238660 270684 238672
rect 252980 238632 261248 238660
rect 263888 238632 270684 238660
rect 252980 238620 252986 238632
rect 239232 238564 243124 238592
rect 246666 238552 246672 238604
rect 246724 238592 246730 238604
rect 255222 238592 255228 238604
rect 246724 238564 255228 238592
rect 246724 238552 246730 238564
rect 255222 238552 255228 238564
rect 255280 238552 255286 238604
rect 257154 238552 257160 238604
rect 257212 238592 257218 238604
rect 257982 238592 257988 238604
rect 257212 238564 257988 238592
rect 257212 238552 257218 238564
rect 257982 238552 257988 238564
rect 258040 238552 258046 238604
rect 259730 238552 259736 238604
rect 259788 238592 259794 238604
rect 263888 238592 263916 238632
rect 270678 238620 270684 238632
rect 270736 238620 270742 238672
rect 259788 238564 263916 238592
rect 259788 238552 259794 238564
rect 263962 238552 263968 238604
rect 264020 238592 264026 238604
rect 264974 238592 264980 238604
rect 264020 238564 264980 238592
rect 264020 238552 264026 238564
rect 264974 238552 264980 238564
rect 265032 238552 265038 238604
rect 265066 238552 265072 238604
rect 265124 238592 265130 238604
rect 278130 238592 278136 238604
rect 265124 238564 278136 238592
rect 265124 238552 265130 238564
rect 278130 238552 278136 238564
rect 278188 238592 278194 238604
rect 278188 238564 282914 238592
rect 278188 238552 278194 238564
rect 209038 238484 209044 238536
rect 209096 238524 209102 238536
rect 221366 238524 221372 238536
rect 209096 238496 221372 238524
rect 209096 238484 209102 238496
rect 221366 238484 221372 238496
rect 221424 238484 221430 238536
rect 224862 238484 224868 238536
rect 224920 238524 224926 238536
rect 226978 238524 226984 238536
rect 224920 238496 226984 238524
rect 224920 238484 224926 238496
rect 226978 238484 226984 238496
rect 227036 238484 227042 238536
rect 240778 238524 240784 238536
rect 230768 238496 240784 238524
rect 209130 238416 209136 238468
rect 209188 238456 209194 238468
rect 229278 238456 229284 238468
rect 209188 238428 229284 238456
rect 209188 238416 209194 238428
rect 229278 238416 229284 238428
rect 229336 238416 229342 238468
rect 193766 238348 193772 238400
rect 193824 238388 193830 238400
rect 224310 238388 224316 238400
rect 193824 238360 224316 238388
rect 193824 238348 193830 238360
rect 224310 238348 224316 238360
rect 224368 238348 224374 238400
rect 230768 238388 230796 238496
rect 240778 238484 240784 238496
rect 240836 238484 240842 238536
rect 241514 238484 241520 238536
rect 241572 238524 241578 238536
rect 245654 238524 245660 238536
rect 241572 238496 245660 238524
rect 241572 238484 241578 238496
rect 245654 238484 245660 238496
rect 245712 238484 245718 238536
rect 246850 238484 246856 238536
rect 246908 238524 246914 238536
rect 250162 238524 250168 238536
rect 246908 238496 250168 238524
rect 246908 238484 246914 238496
rect 250162 238484 250168 238496
rect 250220 238484 250226 238536
rect 250990 238484 250996 238536
rect 251048 238524 251054 238536
rect 251174 238524 251180 238536
rect 251048 238496 251180 238524
rect 251048 238484 251054 238496
rect 251174 238484 251180 238496
rect 251232 238484 251238 238536
rect 255130 238484 255136 238536
rect 255188 238524 255194 238536
rect 256694 238524 256700 238536
rect 255188 238496 256700 238524
rect 255188 238484 255194 238496
rect 256694 238484 256700 238496
rect 256752 238484 256758 238536
rect 259546 238484 259552 238536
rect 259604 238524 259610 238536
rect 269114 238524 269120 238536
rect 259604 238496 269120 238524
rect 259604 238484 259610 238496
rect 269114 238484 269120 238496
rect 269172 238484 269178 238536
rect 282886 238524 282914 238564
rect 296254 238524 296260 238536
rect 282886 238496 296260 238524
rect 296254 238484 296260 238496
rect 296312 238484 296318 238536
rect 230842 238416 230848 238468
rect 230900 238456 230906 238468
rect 268562 238456 268568 238468
rect 230900 238428 244504 238456
rect 230900 238416 230906 238428
rect 225432 238360 230796 238388
rect 161106 238280 161112 238332
rect 161164 238320 161170 238332
rect 210602 238320 210608 238332
rect 161164 238292 210608 238320
rect 161164 238280 161170 238292
rect 210602 238280 210608 238292
rect 210660 238280 210666 238332
rect 219710 238280 219716 238332
rect 219768 238320 219774 238332
rect 220538 238320 220544 238332
rect 219768 238292 220544 238320
rect 219768 238280 219774 238292
rect 220538 238280 220544 238292
rect 220596 238280 220602 238332
rect 222746 238280 222752 238332
rect 222804 238320 222810 238332
rect 225432 238320 225460 238360
rect 232590 238348 232596 238400
rect 232648 238388 232654 238400
rect 236638 238388 236644 238400
rect 232648 238360 236644 238388
rect 232648 238348 232654 238360
rect 236638 238348 236644 238360
rect 236696 238348 236702 238400
rect 239030 238348 239036 238400
rect 239088 238388 239094 238400
rect 241514 238388 241520 238400
rect 239088 238360 241520 238388
rect 239088 238348 239094 238360
rect 241514 238348 241520 238360
rect 241572 238348 241578 238400
rect 222804 238292 225460 238320
rect 222804 238280 222810 238292
rect 227898 238280 227904 238332
rect 227956 238320 227962 238332
rect 228082 238320 228088 238332
rect 227956 238292 228088 238320
rect 227956 238280 227962 238292
rect 228082 238280 228088 238292
rect 228140 238280 228146 238332
rect 228910 238280 228916 238332
rect 228968 238320 228974 238332
rect 240502 238320 240508 238332
rect 228968 238292 240508 238320
rect 228968 238280 228974 238292
rect 240502 238280 240508 238292
rect 240560 238280 240566 238332
rect 243722 238280 243728 238332
rect 243780 238280 243786 238332
rect 244476 238320 244504 238428
rect 248248 238428 268568 238456
rect 248248 238320 248276 238428
rect 268562 238416 268568 238428
rect 268620 238416 268626 238468
rect 273530 238416 273536 238468
rect 273588 238456 273594 238468
rect 295242 238456 295248 238468
rect 273588 238428 295248 238456
rect 273588 238416 273594 238428
rect 295242 238416 295248 238428
rect 295300 238416 295306 238468
rect 261570 238388 261576 238400
rect 244476 238292 248276 238320
rect 248340 238360 261576 238388
rect 192478 238212 192484 238264
rect 192536 238252 192542 238264
rect 219894 238252 219900 238264
rect 192536 238224 219900 238252
rect 192536 238212 192542 238224
rect 219894 238212 219900 238224
rect 219952 238212 219958 238264
rect 222930 238212 222936 238264
rect 222988 238252 222994 238264
rect 230382 238252 230388 238264
rect 222988 238224 230388 238252
rect 222988 238212 222994 238224
rect 230382 238212 230388 238224
rect 230440 238212 230446 238264
rect 231762 238252 231768 238264
rect 231504 238224 231768 238252
rect 210234 238144 210240 238196
rect 210292 238184 210298 238196
rect 231504 238184 231532 238224
rect 231762 238212 231768 238224
rect 231820 238212 231826 238264
rect 234890 238212 234896 238264
rect 234948 238252 234954 238264
rect 237650 238252 237656 238264
rect 234948 238224 237656 238252
rect 234948 238212 234954 238224
rect 237650 238212 237656 238224
rect 237708 238212 237714 238264
rect 243740 238252 243768 238280
rect 248340 238252 248368 238360
rect 261570 238348 261576 238360
rect 261628 238348 261634 238400
rect 302970 238388 302976 238400
rect 263704 238360 302976 238388
rect 248874 238280 248880 238332
rect 248932 238320 248938 238332
rect 259730 238320 259736 238332
rect 248932 238292 259736 238320
rect 248932 238280 248938 238292
rect 259730 238280 259736 238292
rect 259788 238280 259794 238332
rect 262214 238280 262220 238332
rect 262272 238320 262278 238332
rect 263594 238320 263600 238332
rect 262272 238292 263600 238320
rect 262272 238280 262278 238292
rect 263594 238280 263600 238292
rect 263652 238280 263658 238332
rect 243740 238224 248368 238252
rect 255222 238212 255228 238264
rect 255280 238252 255286 238264
rect 263042 238252 263048 238264
rect 255280 238224 263048 238252
rect 255280 238212 255286 238224
rect 263042 238212 263048 238224
rect 263100 238212 263106 238264
rect 210292 238156 231532 238184
rect 210292 238144 210298 238156
rect 231578 238144 231584 238196
rect 231636 238184 231642 238196
rect 243722 238184 243728 238196
rect 231636 238156 243728 238184
rect 231636 238144 231642 238156
rect 243722 238144 243728 238156
rect 243780 238144 243786 238196
rect 259362 238144 259368 238196
rect 259420 238184 259426 238196
rect 263704 238184 263732 238360
rect 302970 238348 302976 238360
rect 303028 238348 303034 238400
rect 265066 238280 265072 238332
rect 265124 238320 265130 238332
rect 265434 238320 265440 238332
rect 265124 238292 265440 238320
rect 265124 238280 265130 238292
rect 265434 238280 265440 238292
rect 265492 238280 265498 238332
rect 266446 238280 266452 238332
rect 266504 238320 266510 238332
rect 266814 238320 266820 238332
rect 266504 238292 266820 238320
rect 266504 238280 266510 238292
rect 266814 238280 266820 238292
rect 266872 238280 266878 238332
rect 267458 238280 267464 238332
rect 267516 238320 267522 238332
rect 268194 238320 268200 238332
rect 267516 238292 268200 238320
rect 267516 238280 267522 238292
rect 268194 238280 268200 238292
rect 268252 238280 268258 238332
rect 268470 238280 268476 238332
rect 268528 238320 268534 238332
rect 310238 238320 310244 238332
rect 268528 238292 310244 238320
rect 268528 238280 268534 238292
rect 310238 238280 310244 238292
rect 310296 238280 310302 238332
rect 269114 238212 269120 238264
rect 269172 238252 269178 238264
rect 316954 238252 316960 238264
rect 269172 238224 316960 238252
rect 269172 238212 269178 238224
rect 316954 238212 316960 238224
rect 317012 238212 317018 238264
rect 259420 238156 263732 238184
rect 259420 238144 259426 238156
rect 264422 238144 264428 238196
rect 264480 238184 264486 238196
rect 265802 238184 265808 238196
rect 264480 238156 265808 238184
rect 264480 238144 264486 238156
rect 265802 238144 265808 238156
rect 265860 238144 265866 238196
rect 266998 238144 267004 238196
rect 267056 238184 267062 238196
rect 315390 238184 315396 238196
rect 267056 238156 315396 238184
rect 267056 238144 267062 238156
rect 315390 238144 315396 238156
rect 315448 238144 315454 238196
rect 161198 238076 161204 238128
rect 161256 238116 161262 238128
rect 212350 238116 212356 238128
rect 161256 238088 212356 238116
rect 161256 238076 161262 238088
rect 212350 238076 212356 238088
rect 212408 238076 212414 238128
rect 220538 238076 220544 238128
rect 220596 238116 220602 238128
rect 230658 238116 230664 238128
rect 220596 238088 230664 238116
rect 220596 238076 220602 238088
rect 230658 238076 230664 238088
rect 230716 238076 230722 238128
rect 231302 238076 231308 238128
rect 231360 238116 231366 238128
rect 231486 238116 231492 238128
rect 231360 238088 231492 238116
rect 231360 238076 231366 238088
rect 231486 238076 231492 238088
rect 231544 238116 231550 238128
rect 239306 238116 239312 238128
rect 231544 238088 239312 238116
rect 231544 238076 231550 238088
rect 239306 238076 239312 238088
rect 239364 238076 239370 238128
rect 239490 238076 239496 238128
rect 239548 238116 239554 238128
rect 248138 238116 248144 238128
rect 239548 238088 248144 238116
rect 239548 238076 239554 238088
rect 248138 238076 248144 238088
rect 248196 238076 248202 238128
rect 249334 238076 249340 238128
rect 249392 238116 249398 238128
rect 260282 238116 260288 238128
rect 249392 238088 260288 238116
rect 249392 238076 249398 238088
rect 260282 238076 260288 238088
rect 260340 238076 260346 238128
rect 260374 238076 260380 238128
rect 260432 238116 260438 238128
rect 266814 238116 266820 238128
rect 260432 238088 266820 238116
rect 260432 238076 260438 238088
rect 266814 238076 266820 238088
rect 266872 238076 266878 238128
rect 269758 238116 269764 238128
rect 268304 238088 269764 238116
rect 161290 238008 161296 238060
rect 161348 238048 161354 238060
rect 237742 238048 237748 238060
rect 161348 238020 237748 238048
rect 161348 238008 161354 238020
rect 237742 238008 237748 238020
rect 237800 238048 237806 238060
rect 242526 238048 242532 238060
rect 237800 238020 242532 238048
rect 237800 238008 237806 238020
rect 242526 238008 242532 238020
rect 242584 238008 242590 238060
rect 245470 238008 245476 238060
rect 245528 238048 245534 238060
rect 251726 238048 251732 238060
rect 245528 238020 251732 238048
rect 245528 238008 245534 238020
rect 251726 238008 251732 238020
rect 251784 238008 251790 238060
rect 255406 238008 255412 238060
rect 255464 238048 255470 238060
rect 268194 238048 268200 238060
rect 255464 238020 268200 238048
rect 255464 238008 255470 238020
rect 268194 238008 268200 238020
rect 268252 238008 268258 238060
rect 217962 237940 217968 237992
rect 218020 237980 218026 237992
rect 218882 237980 218888 237992
rect 218020 237952 218888 237980
rect 218020 237940 218026 237952
rect 218882 237940 218888 237952
rect 218940 237980 218946 237992
rect 223206 237980 223212 237992
rect 218940 237952 223212 237980
rect 218940 237940 218946 237952
rect 223206 237940 223212 237952
rect 223264 237940 223270 237992
rect 225598 237940 225604 237992
rect 225656 237980 225662 237992
rect 234430 237980 234436 237992
rect 225656 237952 234436 237980
rect 225656 237940 225662 237952
rect 234430 237940 234436 237952
rect 234488 237940 234494 237992
rect 235442 237940 235448 237992
rect 235500 237980 235506 237992
rect 236086 237980 236092 237992
rect 235500 237952 236092 237980
rect 235500 237940 235506 237952
rect 236086 237940 236092 237952
rect 236144 237940 236150 237992
rect 236638 237940 236644 237992
rect 236696 237980 236702 237992
rect 236696 237952 251404 237980
rect 236696 237940 236702 237952
rect 210602 237872 210608 237924
rect 210660 237912 210666 237924
rect 234614 237912 234620 237924
rect 210660 237884 234620 237912
rect 210660 237872 210666 237884
rect 234614 237872 234620 237884
rect 234672 237872 234678 237924
rect 237006 237872 237012 237924
rect 237064 237912 237070 237924
rect 237650 237912 237656 237924
rect 237064 237884 237656 237912
rect 237064 237872 237070 237884
rect 237650 237872 237656 237884
rect 237708 237872 237714 237924
rect 238018 237872 238024 237924
rect 238076 237912 238082 237924
rect 240226 237912 240232 237924
rect 238076 237884 240232 237912
rect 238076 237872 238082 237884
rect 240226 237872 240232 237884
rect 240284 237872 240290 237924
rect 240502 237872 240508 237924
rect 240560 237912 240566 237924
rect 249058 237912 249064 237924
rect 240560 237884 249064 237912
rect 240560 237872 240566 237884
rect 249058 237872 249064 237884
rect 249116 237872 249122 237924
rect 251376 237912 251404 237952
rect 251450 237940 251456 237992
rect 251508 237980 251514 237992
rect 252830 237980 252836 237992
rect 251508 237952 252836 237980
rect 251508 237940 251514 237952
rect 252830 237940 252836 237952
rect 252888 237940 252894 237992
rect 254670 237940 254676 237992
rect 254728 237980 254734 237992
rect 261294 237980 261300 237992
rect 254728 237952 261300 237980
rect 254728 237940 254734 237952
rect 261294 237940 261300 237952
rect 261352 237940 261358 237992
rect 266722 237940 266728 237992
rect 266780 237980 266786 237992
rect 268304 237980 268332 238088
rect 269758 238076 269764 238088
rect 269816 238076 269822 238128
rect 269850 238076 269856 238128
rect 269908 238116 269914 238128
rect 318334 238116 318340 238128
rect 269908 238088 318340 238116
rect 269908 238076 269914 238088
rect 318334 238076 318340 238088
rect 318392 238076 318398 238128
rect 268654 238008 268660 238060
rect 268712 238048 268718 238060
rect 338390 238048 338396 238060
rect 268712 238020 338396 238048
rect 268712 238008 268718 238020
rect 338390 238008 338396 238020
rect 338448 238008 338454 238060
rect 266780 237952 268332 237980
rect 266780 237940 266786 237952
rect 268378 237940 268384 237992
rect 268436 237980 268442 237992
rect 273530 237980 273536 237992
rect 268436 237952 273536 237980
rect 268436 237940 268442 237952
rect 273530 237940 273536 237952
rect 273588 237940 273594 237992
rect 258442 237912 258448 237924
rect 251376 237884 258448 237912
rect 258442 237872 258448 237884
rect 258500 237872 258506 237924
rect 263410 237872 263416 237924
rect 263468 237912 263474 237924
rect 274266 237912 274272 237924
rect 263468 237884 274272 237912
rect 263468 237872 263474 237884
rect 274266 237872 274272 237884
rect 274324 237872 274330 237924
rect 212350 237804 212356 237856
rect 212408 237844 212414 237856
rect 236270 237844 236276 237856
rect 212408 237816 236276 237844
rect 212408 237804 212414 237816
rect 236270 237804 236276 237816
rect 236328 237804 236334 237856
rect 239214 237804 239220 237856
rect 239272 237844 239278 237856
rect 239272 237816 244872 237844
rect 239272 237804 239278 237816
rect 208854 237736 208860 237788
rect 208912 237776 208918 237788
rect 226610 237776 226616 237788
rect 208912 237748 226616 237776
rect 208912 237736 208918 237748
rect 226610 237736 226616 237748
rect 226668 237736 226674 237788
rect 226702 237736 226708 237788
rect 226760 237776 226766 237788
rect 227070 237776 227076 237788
rect 226760 237748 227076 237776
rect 226760 237736 226766 237748
rect 227070 237736 227076 237748
rect 227128 237736 227134 237788
rect 227438 237736 227444 237788
rect 227496 237776 227502 237788
rect 236914 237776 236920 237788
rect 227496 237748 236920 237776
rect 227496 237736 227502 237748
rect 236914 237736 236920 237748
rect 236972 237776 236978 237788
rect 240226 237776 240232 237788
rect 236972 237748 240232 237776
rect 236972 237736 236978 237748
rect 240226 237736 240232 237748
rect 240284 237736 240290 237788
rect 244844 237776 244872 237816
rect 251450 237804 251456 237856
rect 251508 237844 251514 237856
rect 251634 237844 251640 237856
rect 251508 237816 251640 237844
rect 251508 237804 251514 237816
rect 251634 237804 251640 237816
rect 251692 237804 251698 237856
rect 261570 237804 261576 237856
rect 261628 237844 261634 237856
rect 268930 237844 268936 237856
rect 261628 237816 268936 237844
rect 261628 237804 261634 237816
rect 268930 237804 268936 237816
rect 268988 237804 268994 237856
rect 269022 237776 269028 237788
rect 244844 237748 269028 237776
rect 269022 237736 269028 237748
rect 269080 237736 269086 237788
rect 238386 237708 238392 237720
rect 225800 237680 238392 237708
rect 161934 237464 161940 237516
rect 161992 237504 161998 237516
rect 225414 237504 225420 237516
rect 161992 237476 225420 237504
rect 161992 237464 161998 237476
rect 225414 237464 225420 237476
rect 225472 237464 225478 237516
rect 161382 237396 161388 237448
rect 161440 237436 161446 237448
rect 225800 237436 225828 237680
rect 238386 237668 238392 237680
rect 238444 237668 238450 237720
rect 238726 237680 239352 237708
rect 232130 237600 232136 237652
rect 232188 237640 232194 237652
rect 238726 237640 238754 237680
rect 232188 237612 238754 237640
rect 239324 237640 239352 237680
rect 240134 237668 240140 237720
rect 240192 237708 240198 237720
rect 241698 237708 241704 237720
rect 240192 237680 241704 237708
rect 240192 237668 240198 237680
rect 241698 237668 241704 237680
rect 241756 237668 241762 237720
rect 243722 237668 243728 237720
rect 243780 237708 243786 237720
rect 270402 237708 270408 237720
rect 243780 237680 270408 237708
rect 243780 237668 243786 237680
rect 270402 237668 270408 237680
rect 270460 237668 270466 237720
rect 261570 237640 261576 237652
rect 239324 237612 261576 237640
rect 232188 237600 232194 237612
rect 261570 237600 261576 237612
rect 261628 237600 261634 237652
rect 263686 237600 263692 237652
rect 263744 237640 263750 237652
rect 264698 237640 264704 237652
rect 263744 237612 264704 237640
rect 263744 237600 263750 237612
rect 264698 237600 264704 237612
rect 264756 237600 264762 237652
rect 265066 237600 265072 237652
rect 265124 237640 265130 237652
rect 265342 237640 265348 237652
rect 265124 237612 265348 237640
rect 265124 237600 265130 237612
rect 265342 237600 265348 237612
rect 265400 237600 265406 237652
rect 265526 237600 265532 237652
rect 265584 237640 265590 237652
rect 266170 237640 266176 237652
rect 265584 237612 266176 237640
rect 265584 237600 265590 237612
rect 266170 237600 266176 237612
rect 266228 237600 266234 237652
rect 226610 237532 226616 237584
rect 226668 237572 226674 237584
rect 226886 237572 226892 237584
rect 226668 237544 226892 237572
rect 226668 237532 226674 237544
rect 226886 237532 226892 237544
rect 226944 237532 226950 237584
rect 231670 237532 231676 237584
rect 231728 237572 231734 237584
rect 239214 237572 239220 237584
rect 231728 237544 239220 237572
rect 231728 237532 231734 237544
rect 239214 237532 239220 237544
rect 239272 237532 239278 237584
rect 239508 237544 256694 237572
rect 235994 237504 236000 237516
rect 161440 237408 225828 237436
rect 225892 237476 236000 237504
rect 161440 237396 161446 237408
rect 225414 237328 225420 237380
rect 225472 237368 225478 237380
rect 225892 237368 225920 237476
rect 235994 237464 236000 237476
rect 236052 237464 236058 237516
rect 239306 237464 239312 237516
rect 239364 237504 239370 237516
rect 239508 237504 239536 237544
rect 239364 237476 239536 237504
rect 256666 237504 256694 237544
rect 257798 237532 257804 237584
rect 257856 237572 257862 237584
rect 263502 237572 263508 237584
rect 257856 237544 263508 237572
rect 257856 237532 257862 237544
rect 263502 237532 263508 237544
rect 263560 237532 263566 237584
rect 264238 237532 264244 237584
rect 264296 237572 264302 237584
rect 272702 237572 272708 237584
rect 264296 237544 272708 237572
rect 264296 237532 264302 237544
rect 272702 237532 272708 237544
rect 272760 237532 272766 237584
rect 266722 237504 266728 237516
rect 256666 237476 266728 237504
rect 239364 237464 239370 237476
rect 266722 237464 266728 237476
rect 266780 237464 266786 237516
rect 266814 237464 266820 237516
rect 266872 237504 266878 237516
rect 266872 237476 276014 237504
rect 266872 237464 266878 237476
rect 229370 237396 229376 237448
rect 229428 237436 229434 237448
rect 230106 237436 230112 237448
rect 229428 237408 230112 237436
rect 229428 237396 229434 237408
rect 230106 237396 230112 237408
rect 230164 237396 230170 237448
rect 239030 237396 239036 237448
rect 239088 237436 239094 237448
rect 244182 237436 244188 237448
rect 239088 237408 244188 237436
rect 239088 237396 239094 237408
rect 244182 237396 244188 237408
rect 244240 237396 244246 237448
rect 253566 237396 253572 237448
rect 253624 237436 253630 237448
rect 254670 237436 254676 237448
rect 253624 237408 254676 237436
rect 253624 237396 253630 237408
rect 254670 237396 254676 237408
rect 254728 237396 254734 237448
rect 263704 237408 264652 237436
rect 225472 237340 225920 237368
rect 225472 237328 225478 237340
rect 229278 237328 229284 237380
rect 229336 237368 229342 237380
rect 230198 237368 230204 237380
rect 229336 237340 230204 237368
rect 229336 237328 229342 237340
rect 230198 237328 230204 237340
rect 230256 237328 230262 237380
rect 230750 237328 230756 237380
rect 230808 237368 230814 237380
rect 231762 237368 231768 237380
rect 230808 237340 231768 237368
rect 230808 237328 230814 237340
rect 231762 237328 231768 237340
rect 231820 237328 231826 237380
rect 239122 237368 239128 237380
rect 234816 237340 239128 237368
rect 215846 237260 215852 237312
rect 215904 237300 215910 237312
rect 220262 237300 220268 237312
rect 215904 237272 220268 237300
rect 215904 237260 215910 237272
rect 220262 237260 220268 237272
rect 220320 237300 220326 237312
rect 234816 237300 234844 237340
rect 239122 237328 239128 237340
rect 239180 237328 239186 237380
rect 258626 237328 258632 237380
rect 258684 237368 258690 237380
rect 259270 237368 259276 237380
rect 258684 237340 259276 237368
rect 258684 237328 258690 237340
rect 259270 237328 259276 237340
rect 259328 237328 259334 237380
rect 261018 237328 261024 237380
rect 261076 237368 261082 237380
rect 263704 237368 263732 237408
rect 261076 237340 263732 237368
rect 264624 237368 264652 237408
rect 264974 237396 264980 237448
rect 265032 237436 265038 237448
rect 275986 237436 276014 237476
rect 288526 237436 288532 237448
rect 265032 237408 267780 237436
rect 275986 237408 288532 237436
rect 265032 237396 265038 237408
rect 267274 237368 267280 237380
rect 264624 237340 267280 237368
rect 261076 237328 261082 237340
rect 267274 237328 267280 237340
rect 267332 237328 267338 237380
rect 267752 237368 267780 237408
rect 288526 237396 288532 237408
rect 288584 237436 288590 237448
rect 288986 237436 288992 237448
rect 288584 237408 288992 237436
rect 288584 237396 288590 237408
rect 288986 237396 288992 237408
rect 289044 237396 289050 237448
rect 299014 237396 299020 237448
rect 299072 237436 299078 237448
rect 301682 237436 301688 237448
rect 299072 237408 301688 237436
rect 299072 237396 299078 237408
rect 301682 237396 301688 237408
rect 301740 237396 301746 237448
rect 268838 237368 268844 237380
rect 267752 237340 268844 237368
rect 268838 237328 268844 237340
rect 268896 237368 268902 237380
rect 268896 237340 273254 237368
rect 268896 237328 268902 237340
rect 220320 237272 234844 237300
rect 220320 237260 220326 237272
rect 235350 237260 235356 237312
rect 235408 237300 235414 237312
rect 235718 237300 235724 237312
rect 235408 237272 235724 237300
rect 235408 237260 235414 237272
rect 235718 237260 235724 237272
rect 235776 237260 235782 237312
rect 243722 237260 243728 237312
rect 243780 237300 243786 237312
rect 243998 237300 244004 237312
rect 243780 237272 244004 237300
rect 243780 237260 243786 237272
rect 243998 237260 244004 237272
rect 244056 237260 244062 237312
rect 251174 237260 251180 237312
rect 251232 237300 251238 237312
rect 251450 237300 251456 237312
rect 251232 237272 251456 237300
rect 251232 237260 251238 237272
rect 251450 237260 251456 237272
rect 251508 237260 251514 237312
rect 253566 237260 253572 237312
rect 253624 237300 253630 237312
rect 268470 237300 268476 237312
rect 253624 237272 268476 237300
rect 253624 237260 253630 237272
rect 268470 237260 268476 237272
rect 268528 237260 268534 237312
rect 273226 237300 273254 237340
rect 275922 237328 275928 237380
rect 275980 237368 275986 237380
rect 276290 237368 276296 237380
rect 275980 237340 276296 237368
rect 275980 237328 275986 237340
rect 276290 237328 276296 237340
rect 276348 237328 276354 237380
rect 330110 237300 330116 237312
rect 273226 237272 330116 237300
rect 330110 237260 330116 237272
rect 330168 237260 330174 237312
rect 208394 237192 208400 237244
rect 208452 237232 208458 237244
rect 209222 237232 209228 237244
rect 208452 237204 209228 237232
rect 208452 237192 208458 237204
rect 209222 237192 209228 237204
rect 209280 237232 209286 237244
rect 226242 237232 226248 237244
rect 209280 237204 226248 237232
rect 209280 237192 209286 237204
rect 226242 237192 226248 237204
rect 226300 237192 226306 237244
rect 226518 237192 226524 237244
rect 226576 237232 226582 237244
rect 226794 237232 226800 237244
rect 226576 237204 226800 237232
rect 226576 237192 226582 237204
rect 226794 237192 226800 237204
rect 226852 237192 226858 237244
rect 234154 237192 234160 237244
rect 234212 237232 234218 237244
rect 234338 237232 234344 237244
rect 234212 237204 234344 237232
rect 234212 237192 234218 237204
rect 234338 237192 234344 237204
rect 234396 237192 234402 237244
rect 240594 237192 240600 237244
rect 240652 237232 240658 237244
rect 248414 237232 248420 237244
rect 240652 237204 248420 237232
rect 240652 237192 240658 237204
rect 248414 237192 248420 237204
rect 248472 237192 248478 237244
rect 256510 237192 256516 237244
rect 256568 237232 256574 237244
rect 286870 237232 286876 237244
rect 256568 237204 286876 237232
rect 256568 237192 256574 237204
rect 286870 237192 286876 237204
rect 286928 237192 286934 237244
rect 214466 237124 214472 237176
rect 214524 237164 214530 237176
rect 214524 237136 226334 237164
rect 214524 237124 214530 237136
rect 207842 237056 207848 237108
rect 207900 237096 207906 237108
rect 222562 237096 222568 237108
rect 207900 237068 222568 237096
rect 207900 237056 207906 237068
rect 222562 237056 222568 237068
rect 222620 237056 222626 237108
rect 226306 237096 226334 237136
rect 226978 237124 226984 237176
rect 227036 237164 227042 237176
rect 229094 237164 229100 237176
rect 227036 237136 229100 237164
rect 227036 237124 227042 237136
rect 229094 237124 229100 237136
rect 229152 237124 229158 237176
rect 243814 237124 243820 237176
rect 243872 237164 243878 237176
rect 275922 237164 275928 237176
rect 243872 237136 275928 237164
rect 243872 237124 243878 237136
rect 275922 237124 275928 237136
rect 275980 237124 275986 237176
rect 234706 237096 234712 237108
rect 226306 237068 234712 237096
rect 234706 237056 234712 237068
rect 234764 237056 234770 237108
rect 244366 237056 244372 237108
rect 244424 237096 244430 237108
rect 245102 237096 245108 237108
rect 244424 237068 245108 237096
rect 244424 237056 244430 237068
rect 245102 237056 245108 237068
rect 245160 237056 245166 237108
rect 247862 237056 247868 237108
rect 247920 237096 247926 237108
rect 248230 237096 248236 237108
rect 247920 237068 248236 237096
rect 247920 237056 247926 237068
rect 248230 237056 248236 237068
rect 248288 237056 248294 237108
rect 253566 237096 253572 237108
rect 251146 237068 253572 237096
rect 208026 236988 208032 237040
rect 208084 237028 208090 237040
rect 222470 237028 222476 237040
rect 208084 237000 222476 237028
rect 208084 236988 208090 237000
rect 222470 236988 222476 237000
rect 222528 236988 222534 237040
rect 222838 236988 222844 237040
rect 222896 237028 222902 237040
rect 230014 237028 230020 237040
rect 222896 237000 230020 237028
rect 222896 236988 222902 237000
rect 230014 236988 230020 237000
rect 230072 236988 230078 237040
rect 236178 236988 236184 237040
rect 236236 237028 236242 237040
rect 237466 237028 237472 237040
rect 236236 237000 237472 237028
rect 236236 236988 236242 237000
rect 237466 236988 237472 237000
rect 237524 236988 237530 237040
rect 244734 236988 244740 237040
rect 244792 237028 244798 237040
rect 244918 237028 244924 237040
rect 244792 237000 244924 237028
rect 244792 236988 244798 237000
rect 244918 236988 244924 237000
rect 244976 236988 244982 237040
rect 211798 236920 211804 236972
rect 211856 236960 211862 236972
rect 249242 236960 249248 236972
rect 211856 236932 249248 236960
rect 211856 236920 211862 236932
rect 249242 236920 249248 236932
rect 249300 236960 249306 236972
rect 251146 236960 251174 237068
rect 253566 237056 253572 237068
rect 253624 237056 253630 237108
rect 254394 237056 254400 237108
rect 254452 237096 254458 237108
rect 261018 237096 261024 237108
rect 254452 237068 261024 237096
rect 254452 237056 254458 237068
rect 261018 237056 261024 237068
rect 261076 237056 261082 237108
rect 262858 237056 262864 237108
rect 262916 237096 262922 237108
rect 289722 237096 289728 237108
rect 262916 237068 289728 237096
rect 262916 237056 262922 237068
rect 289722 237056 289728 237068
rect 289780 237056 289786 237108
rect 251542 236988 251548 237040
rect 251600 237028 251606 237040
rect 274818 237028 274824 237040
rect 251600 237000 274824 237028
rect 251600 236988 251606 237000
rect 274818 236988 274824 237000
rect 274876 237028 274882 237040
rect 275370 237028 275376 237040
rect 274876 237000 275376 237028
rect 274876 236988 274882 237000
rect 275370 236988 275376 237000
rect 275428 236988 275434 237040
rect 249300 236932 251174 236960
rect 249300 236920 249306 236932
rect 251726 236920 251732 236972
rect 251784 236960 251790 236972
rect 261018 236960 261024 236972
rect 251784 236932 261024 236960
rect 251784 236920 251790 236932
rect 261018 236920 261024 236932
rect 261076 236920 261082 236972
rect 262306 236920 262312 236972
rect 262364 236960 262370 236972
rect 284386 236960 284392 236972
rect 262364 236932 284392 236960
rect 262364 236920 262370 236932
rect 284386 236920 284392 236932
rect 284444 236960 284450 236972
rect 284754 236960 284760 236972
rect 284444 236932 284760 236960
rect 284444 236920 284450 236932
rect 284754 236920 284760 236932
rect 284812 236920 284818 236972
rect 213086 236852 213092 236904
rect 213144 236892 213150 236904
rect 254394 236892 254400 236904
rect 213144 236864 254400 236892
rect 213144 236852 213150 236864
rect 254394 236852 254400 236864
rect 254452 236852 254458 236904
rect 257338 236852 257344 236904
rect 257396 236892 257402 236904
rect 259270 236892 259276 236904
rect 257396 236864 259276 236892
rect 257396 236852 257402 236864
rect 259270 236852 259276 236864
rect 259328 236852 259334 236904
rect 262582 236852 262588 236904
rect 262640 236892 262646 236904
rect 274634 236892 274640 236904
rect 262640 236864 274640 236892
rect 262640 236852 262646 236864
rect 274634 236852 274640 236864
rect 274692 236892 274698 236904
rect 275646 236892 275652 236904
rect 274692 236864 275652 236892
rect 274692 236852 274698 236864
rect 275646 236852 275652 236864
rect 275704 236852 275710 236904
rect 197262 236784 197268 236836
rect 197320 236824 197326 236836
rect 255682 236824 255688 236836
rect 197320 236796 255688 236824
rect 197320 236784 197326 236796
rect 255682 236784 255688 236796
rect 255740 236784 255746 236836
rect 257706 236784 257712 236836
rect 257764 236824 257770 236836
rect 258258 236824 258264 236836
rect 257764 236796 258264 236824
rect 257764 236784 257770 236796
rect 258258 236784 258264 236796
rect 258316 236784 258322 236836
rect 261754 236784 261760 236836
rect 261812 236824 261818 236836
rect 266906 236824 266912 236836
rect 261812 236796 266912 236824
rect 261812 236784 261818 236796
rect 266906 236784 266912 236796
rect 266964 236784 266970 236836
rect 159910 236716 159916 236768
rect 159968 236756 159974 236768
rect 218882 236756 218888 236768
rect 159968 236728 218888 236756
rect 159968 236716 159974 236728
rect 218882 236716 218888 236728
rect 218940 236716 218946 236768
rect 218974 236716 218980 236768
rect 219032 236756 219038 236768
rect 238570 236756 238576 236768
rect 219032 236728 238576 236756
rect 219032 236716 219038 236728
rect 238570 236716 238576 236728
rect 238628 236716 238634 236768
rect 241698 236716 241704 236768
rect 241756 236756 241762 236768
rect 242250 236756 242256 236768
rect 241756 236728 242256 236756
rect 241756 236716 241762 236728
rect 242250 236716 242256 236728
rect 242308 236716 242314 236768
rect 244918 236716 244924 236768
rect 244976 236756 244982 236768
rect 245194 236756 245200 236768
rect 244976 236728 245200 236756
rect 244976 236716 244982 236728
rect 245194 236716 245200 236728
rect 245252 236716 245258 236768
rect 258276 236756 258304 236784
rect 268654 236756 268660 236768
rect 258276 236728 268660 236756
rect 268654 236716 268660 236728
rect 268712 236716 268718 236768
rect 269574 236716 269580 236768
rect 269632 236756 269638 236768
rect 295334 236756 295340 236768
rect 269632 236728 295340 236756
rect 269632 236716 269638 236728
rect 295334 236716 295340 236728
rect 295392 236716 295398 236768
rect 155586 236648 155592 236700
rect 155644 236688 155650 236700
rect 213822 236688 213828 236700
rect 155644 236660 213828 236688
rect 155644 236648 155650 236660
rect 213822 236648 213828 236660
rect 213880 236648 213886 236700
rect 220170 236648 220176 236700
rect 220228 236688 220234 236700
rect 257338 236688 257344 236700
rect 220228 236660 257344 236688
rect 220228 236648 220234 236660
rect 257338 236648 257344 236660
rect 257396 236648 257402 236700
rect 258258 236648 258264 236700
rect 258316 236688 258322 236700
rect 258902 236688 258908 236700
rect 258316 236660 258908 236688
rect 258316 236648 258322 236660
rect 258902 236648 258908 236660
rect 258960 236648 258966 236700
rect 265434 236648 265440 236700
rect 265492 236688 265498 236700
rect 287974 236688 287980 236700
rect 265492 236660 287980 236688
rect 265492 236648 265498 236660
rect 287974 236648 287980 236660
rect 288032 236688 288038 236700
rect 334986 236688 334992 236700
rect 288032 236660 334992 236688
rect 288032 236648 288038 236660
rect 334986 236648 334992 236660
rect 335044 236648 335050 236700
rect 209498 236580 209504 236632
rect 209556 236620 209562 236632
rect 227806 236620 227812 236632
rect 209556 236592 227812 236620
rect 209556 236580 209562 236592
rect 227806 236580 227812 236592
rect 227864 236620 227870 236632
rect 227990 236620 227996 236632
rect 227864 236592 227996 236620
rect 227864 236580 227870 236592
rect 227990 236580 227996 236592
rect 228048 236580 228054 236632
rect 229094 236580 229100 236632
rect 229152 236620 229158 236632
rect 231210 236620 231216 236632
rect 229152 236592 231216 236620
rect 229152 236580 229158 236592
rect 231210 236580 231216 236592
rect 231268 236580 231274 236632
rect 237466 236580 237472 236632
rect 237524 236620 237530 236632
rect 237742 236620 237748 236632
rect 237524 236592 237748 236620
rect 237524 236580 237530 236592
rect 237742 236580 237748 236592
rect 237800 236580 237806 236632
rect 242066 236580 242072 236632
rect 242124 236620 242130 236632
rect 242250 236620 242256 236632
rect 242124 236592 242256 236620
rect 242124 236580 242130 236592
rect 242250 236580 242256 236592
rect 242308 236580 242314 236632
rect 243998 236580 244004 236632
rect 244056 236620 244062 236632
rect 244642 236620 244648 236632
rect 244056 236592 244648 236620
rect 244056 236580 244062 236592
rect 244642 236580 244648 236592
rect 244700 236580 244706 236632
rect 247954 236580 247960 236632
rect 248012 236620 248018 236632
rect 248322 236620 248328 236632
rect 248012 236592 248328 236620
rect 248012 236580 248018 236592
rect 248322 236580 248328 236592
rect 248380 236580 248386 236632
rect 248966 236580 248972 236632
rect 249024 236620 249030 236632
rect 249702 236620 249708 236632
rect 249024 236592 249708 236620
rect 249024 236580 249030 236592
rect 249702 236580 249708 236592
rect 249760 236580 249766 236632
rect 252830 236580 252836 236632
rect 252888 236620 252894 236632
rect 265526 236620 265532 236632
rect 252888 236592 265532 236620
rect 252888 236580 252894 236592
rect 265526 236580 265532 236592
rect 265584 236580 265590 236632
rect 213822 236512 213828 236564
rect 213880 236552 213886 236564
rect 213880 236524 224632 236552
rect 213880 236512 213886 236524
rect 223942 236444 223948 236496
rect 224000 236484 224006 236496
rect 224310 236484 224316 236496
rect 224000 236456 224316 236484
rect 224000 236444 224006 236456
rect 224310 236444 224316 236456
rect 224368 236444 224374 236496
rect 224604 236484 224632 236524
rect 224678 236512 224684 236564
rect 224736 236552 224742 236564
rect 224862 236552 224868 236564
rect 224736 236524 224868 236552
rect 224736 236512 224742 236524
rect 224862 236512 224868 236524
rect 224920 236512 224926 236564
rect 230750 236512 230756 236564
rect 230808 236552 230814 236564
rect 230934 236552 230940 236564
rect 230808 236524 230940 236552
rect 230808 236512 230814 236524
rect 230934 236512 230940 236524
rect 230992 236512 230998 236564
rect 241882 236512 241888 236564
rect 241940 236552 241946 236564
rect 242434 236552 242440 236564
rect 241940 236524 242440 236552
rect 241940 236512 241946 236524
rect 242434 236512 242440 236524
rect 242492 236512 242498 236564
rect 253474 236512 253480 236564
rect 253532 236552 253538 236564
rect 262766 236552 262772 236564
rect 253532 236524 262772 236552
rect 253532 236512 253538 236524
rect 262766 236512 262772 236524
rect 262824 236512 262830 236564
rect 269850 236552 269856 236564
rect 266740 236524 269856 236552
rect 226058 236484 226064 236496
rect 224604 236456 226064 236484
rect 226058 236444 226064 236456
rect 226116 236444 226122 236496
rect 258442 236444 258448 236496
rect 258500 236484 258506 236496
rect 266740 236484 266768 236524
rect 269850 236512 269856 236524
rect 269908 236512 269914 236564
rect 258500 236456 266768 236484
rect 258500 236444 258506 236456
rect 223758 236376 223764 236428
rect 223816 236416 223822 236428
rect 226334 236416 226340 236428
rect 223816 236388 226340 236416
rect 223816 236376 223822 236388
rect 226334 236376 226340 236388
rect 226392 236376 226398 236428
rect 238202 236376 238208 236428
rect 238260 236416 238266 236428
rect 247862 236416 247868 236428
rect 238260 236388 247868 236416
rect 238260 236376 238266 236388
rect 247862 236376 247868 236388
rect 247920 236416 247926 236428
rect 327718 236416 327724 236428
rect 247920 236388 327724 236416
rect 247920 236376 247926 236388
rect 327718 236376 327724 236388
rect 327776 236376 327782 236428
rect 265894 236308 265900 236360
rect 265952 236348 265958 236360
rect 266814 236348 266820 236360
rect 265952 236320 266820 236348
rect 265952 236308 265958 236320
rect 266814 236308 266820 236320
rect 266872 236308 266878 236360
rect 245102 236240 245108 236292
rect 245160 236280 245166 236292
rect 245562 236280 245568 236292
rect 245160 236252 245568 236280
rect 245160 236240 245166 236252
rect 245562 236240 245568 236252
rect 245620 236240 245626 236292
rect 261018 236240 261024 236292
rect 261076 236280 261082 236292
rect 261846 236280 261852 236292
rect 261076 236252 261852 236280
rect 261076 236240 261082 236252
rect 261846 236240 261852 236252
rect 261904 236240 261910 236292
rect 214466 236172 214472 236224
rect 214524 236212 214530 236224
rect 215018 236212 215024 236224
rect 214524 236184 215024 236212
rect 214524 236172 214530 236184
rect 215018 236172 215024 236184
rect 215076 236172 215082 236224
rect 226426 236104 226432 236156
rect 226484 236144 226490 236156
rect 227622 236144 227628 236156
rect 226484 236116 227628 236144
rect 226484 236104 226490 236116
rect 227622 236104 227628 236116
rect 227680 236104 227686 236156
rect 261478 236104 261484 236156
rect 261536 236144 261542 236156
rect 276198 236144 276204 236156
rect 261536 236116 276204 236144
rect 261536 236104 261542 236116
rect 276198 236104 276204 236116
rect 276256 236104 276262 236156
rect 261202 236036 261208 236088
rect 261260 236076 261266 236088
rect 267274 236076 267280 236088
rect 261260 236048 267280 236076
rect 261260 236036 261266 236048
rect 267274 236036 267280 236048
rect 267332 236036 267338 236088
rect 207750 235968 207756 236020
rect 207808 236008 207814 236020
rect 208026 236008 208032 236020
rect 207808 235980 208032 236008
rect 207808 235968 207814 235980
rect 208026 235968 208032 235980
rect 208084 235968 208090 236020
rect 217686 235968 217692 236020
rect 217744 236008 217750 236020
rect 244642 236008 244648 236020
rect 217744 235980 244648 236008
rect 217744 235968 217750 235980
rect 244642 235968 244648 235980
rect 244700 235968 244706 236020
rect 255314 235968 255320 236020
rect 255372 236008 255378 236020
rect 255682 236008 255688 236020
rect 255372 235980 255688 236008
rect 255372 235968 255378 235980
rect 255682 235968 255688 235980
rect 255740 235968 255746 236020
rect 285582 235968 285588 236020
rect 285640 236008 285646 236020
rect 286870 236008 286876 236020
rect 285640 235980 286876 236008
rect 285640 235968 285646 235980
rect 286870 235968 286876 235980
rect 286928 235968 286934 236020
rect 289354 235968 289360 236020
rect 289412 236008 289418 236020
rect 289722 236008 289728 236020
rect 289412 235980 289728 236008
rect 289412 235968 289418 235980
rect 289722 235968 289728 235980
rect 289780 235968 289786 236020
rect 210878 235900 210884 235952
rect 210936 235940 210942 235952
rect 210936 235912 215294 235940
rect 210936 235900 210942 235912
rect 215266 235872 215294 235912
rect 217318 235900 217324 235952
rect 217376 235940 217382 235952
rect 219158 235940 219164 235952
rect 217376 235912 219164 235940
rect 217376 235900 217382 235912
rect 219158 235900 219164 235912
rect 219216 235900 219222 235952
rect 221826 235900 221832 235952
rect 221884 235940 221890 235952
rect 222010 235940 222016 235952
rect 221884 235912 222016 235940
rect 221884 235900 221890 235912
rect 222010 235900 222016 235912
rect 222068 235900 222074 235952
rect 233418 235900 233424 235952
rect 233476 235940 233482 235952
rect 233694 235940 233700 235952
rect 233476 235912 233700 235940
rect 233476 235900 233482 235912
rect 233694 235900 233700 235912
rect 233752 235900 233758 235952
rect 233878 235900 233884 235952
rect 233936 235940 233942 235952
rect 237466 235940 237472 235952
rect 233936 235912 237472 235940
rect 233936 235900 233942 235912
rect 237466 235900 237472 235912
rect 237524 235900 237530 235952
rect 253106 235900 253112 235952
rect 253164 235940 253170 235952
rect 253658 235940 253664 235952
rect 253164 235912 253664 235940
rect 253164 235900 253170 235912
rect 253658 235900 253664 235912
rect 253716 235900 253722 235952
rect 274542 235900 274548 235952
rect 274600 235940 274606 235952
rect 330018 235940 330024 235952
rect 274600 235912 330024 235940
rect 274600 235900 274606 235912
rect 330018 235900 330024 235912
rect 330076 235900 330082 235952
rect 223758 235872 223764 235884
rect 215266 235844 223764 235872
rect 223758 235832 223764 235844
rect 223816 235832 223822 235884
rect 259822 235832 259828 235884
rect 259880 235872 259886 235884
rect 268286 235872 268292 235884
rect 259880 235844 268292 235872
rect 259880 235832 259886 235844
rect 268286 235832 268292 235844
rect 268344 235832 268350 235884
rect 285674 235832 285680 235884
rect 285732 235872 285738 235884
rect 286962 235872 286968 235884
rect 285732 235844 286968 235872
rect 285732 235832 285738 235844
rect 286962 235832 286968 235844
rect 287020 235872 287026 235884
rect 287698 235872 287704 235884
rect 287020 235844 287704 235872
rect 287020 235832 287026 235844
rect 287698 235832 287704 235844
rect 287756 235832 287762 235884
rect 240226 235764 240232 235816
rect 240284 235804 240290 235816
rect 276014 235804 276020 235816
rect 240284 235776 276020 235804
rect 240284 235764 240290 235776
rect 276014 235764 276020 235776
rect 276072 235764 276078 235816
rect 223850 235696 223856 235748
rect 223908 235736 223914 235748
rect 224494 235736 224500 235748
rect 223908 235708 224500 235736
rect 223908 235696 223914 235708
rect 224494 235696 224500 235708
rect 224552 235696 224558 235748
rect 226150 235696 226156 235748
rect 226208 235736 226214 235748
rect 226518 235736 226524 235748
rect 226208 235708 226524 235736
rect 226208 235696 226214 235708
rect 226518 235696 226524 235708
rect 226576 235696 226582 235748
rect 244918 235696 244924 235748
rect 244976 235736 244982 235748
rect 291102 235736 291108 235748
rect 244976 235708 291108 235736
rect 244976 235696 244982 235708
rect 291102 235696 291108 235708
rect 291160 235696 291166 235748
rect 235994 235628 236000 235680
rect 236052 235668 236058 235680
rect 279970 235668 279976 235680
rect 236052 235640 279976 235668
rect 236052 235628 236058 235640
rect 279970 235628 279976 235640
rect 280028 235628 280034 235680
rect 220998 235560 221004 235612
rect 221056 235600 221062 235612
rect 233050 235600 233056 235612
rect 221056 235572 233056 235600
rect 221056 235560 221062 235572
rect 233050 235560 233056 235572
rect 233108 235560 233114 235612
rect 244734 235560 244740 235612
rect 244792 235600 244798 235612
rect 285674 235600 285680 235612
rect 244792 235572 285680 235600
rect 244792 235560 244798 235572
rect 285674 235560 285680 235572
rect 285732 235560 285738 235612
rect 222010 235492 222016 235544
rect 222068 235532 222074 235544
rect 230474 235532 230480 235544
rect 222068 235504 230480 235532
rect 222068 235492 222074 235504
rect 230474 235492 230480 235504
rect 230532 235492 230538 235544
rect 232866 235492 232872 235544
rect 232924 235532 232930 235544
rect 234614 235532 234620 235544
rect 232924 235504 234620 235532
rect 232924 235492 232930 235504
rect 234614 235492 234620 235504
rect 234672 235492 234678 235544
rect 242802 235492 242808 235544
rect 242860 235532 242866 235544
rect 283558 235532 283564 235544
rect 242860 235504 283564 235532
rect 242860 235492 242866 235504
rect 283558 235492 283564 235504
rect 283616 235492 283622 235544
rect 216030 235424 216036 235476
rect 216088 235464 216094 235476
rect 236546 235464 236552 235476
rect 216088 235436 236552 235464
rect 216088 235424 216094 235436
rect 236546 235424 236552 235436
rect 236604 235424 236610 235476
rect 243814 235424 243820 235476
rect 243872 235464 243878 235476
rect 248598 235464 248604 235476
rect 243872 235436 248604 235464
rect 243872 235424 243878 235436
rect 248598 235424 248604 235436
rect 248656 235464 248662 235476
rect 269482 235464 269488 235476
rect 248656 235436 269488 235464
rect 248656 235424 248662 235436
rect 269482 235424 269488 235436
rect 269540 235424 269546 235476
rect 269574 235424 269580 235476
rect 269632 235464 269638 235476
rect 270126 235464 270132 235476
rect 269632 235436 270132 235464
rect 269632 235424 269638 235436
rect 270126 235424 270132 235436
rect 270184 235464 270190 235476
rect 282730 235464 282736 235476
rect 270184 235436 282736 235464
rect 270184 235424 270190 235436
rect 282730 235424 282736 235436
rect 282788 235424 282794 235476
rect 211062 235356 211068 235408
rect 211120 235396 211126 235408
rect 220998 235396 221004 235408
rect 211120 235368 221004 235396
rect 211120 235356 211126 235368
rect 220998 235356 221004 235368
rect 221056 235356 221062 235408
rect 239214 235356 239220 235408
rect 239272 235396 239278 235408
rect 239766 235396 239772 235408
rect 239272 235368 239772 235396
rect 239272 235356 239278 235368
rect 239766 235356 239772 235368
rect 239824 235356 239830 235408
rect 243170 235356 243176 235408
rect 243228 235396 243234 235408
rect 262858 235396 262864 235408
rect 243228 235368 262864 235396
rect 243228 235356 243234 235368
rect 262858 235356 262864 235368
rect 262916 235356 262922 235408
rect 268286 235356 268292 235408
rect 268344 235396 268350 235408
rect 270402 235396 270408 235408
rect 268344 235368 270408 235396
rect 268344 235356 268350 235368
rect 270402 235356 270408 235368
rect 270460 235396 270466 235408
rect 280890 235396 280896 235408
rect 270460 235368 280896 235396
rect 270460 235356 270466 235368
rect 280890 235356 280896 235368
rect 280948 235356 280954 235408
rect 218882 235288 218888 235340
rect 218940 235328 218946 235340
rect 244734 235328 244740 235340
rect 218940 235300 244740 235328
rect 218940 235288 218946 235300
rect 244734 235288 244740 235300
rect 244792 235288 244798 235340
rect 253474 235288 253480 235340
rect 253532 235328 253538 235340
rect 253842 235328 253848 235340
rect 253532 235300 253848 235328
rect 253532 235288 253538 235300
rect 253842 235288 253848 235300
rect 253900 235288 253906 235340
rect 262030 235288 262036 235340
rect 262088 235328 262094 235340
rect 277394 235328 277400 235340
rect 262088 235300 277400 235328
rect 262088 235288 262094 235300
rect 277394 235288 277400 235300
rect 277452 235288 277458 235340
rect 219250 235220 219256 235272
rect 219308 235260 219314 235272
rect 255590 235260 255596 235272
rect 219308 235232 255596 235260
rect 219308 235220 219314 235232
rect 255590 235220 255596 235232
rect 255648 235220 255654 235272
rect 263134 235220 263140 235272
rect 263192 235260 263198 235272
rect 282546 235260 282552 235272
rect 263192 235232 282552 235260
rect 263192 235220 263198 235232
rect 282546 235220 282552 235232
rect 282604 235260 282610 235272
rect 331398 235260 331404 235272
rect 282604 235232 331404 235260
rect 282604 235220 282610 235232
rect 331398 235220 331404 235232
rect 331456 235220 331462 235272
rect 239306 235152 239312 235204
rect 239364 235192 239370 235204
rect 240042 235192 240048 235204
rect 239364 235164 240048 235192
rect 239364 235152 239370 235164
rect 240042 235152 240048 235164
rect 240100 235152 240106 235204
rect 243078 235152 243084 235204
rect 243136 235192 243142 235204
rect 243538 235192 243544 235204
rect 243136 235164 243544 235192
rect 243136 235152 243142 235164
rect 243538 235152 243544 235164
rect 243596 235152 243602 235204
rect 252002 235152 252008 235204
rect 252060 235192 252066 235204
rect 265066 235192 265072 235204
rect 252060 235164 265072 235192
rect 252060 235152 252066 235164
rect 265066 235152 265072 235164
rect 265124 235152 265130 235204
rect 267274 235152 267280 235204
rect 267332 235192 267338 235204
rect 269758 235192 269764 235204
rect 267332 235164 269764 235192
rect 267332 235152 267338 235164
rect 269758 235152 269764 235164
rect 269816 235192 269822 235204
rect 278590 235192 278596 235204
rect 269816 235164 278596 235192
rect 269816 235152 269822 235164
rect 278590 235152 278596 235164
rect 278648 235152 278654 235204
rect 227070 235084 227076 235136
rect 227128 235124 227134 235136
rect 239398 235124 239404 235136
rect 227128 235096 239404 235124
rect 227128 235084 227134 235096
rect 239398 235084 239404 235096
rect 239456 235084 239462 235136
rect 254762 235084 254768 235136
rect 254820 235124 254826 235136
rect 269022 235124 269028 235136
rect 254820 235096 269028 235124
rect 254820 235084 254826 235096
rect 269022 235084 269028 235096
rect 269080 235084 269086 235136
rect 216306 235016 216312 235068
rect 216364 235056 216370 235068
rect 227438 235056 227444 235068
rect 216364 235028 227444 235056
rect 216364 235016 216370 235028
rect 227438 235016 227444 235028
rect 227496 235016 227502 235068
rect 240778 235016 240784 235068
rect 240836 235056 240842 235068
rect 300486 235056 300492 235068
rect 240836 235028 300492 235056
rect 240836 235016 240842 235028
rect 300486 235016 300492 235028
rect 300544 235016 300550 235068
rect 216214 234948 216220 235000
rect 216272 234988 216278 235000
rect 216272 234960 224954 234988
rect 216272 234948 216278 234960
rect 210602 234880 210608 234932
rect 210660 234920 210666 234932
rect 217226 234920 217232 234932
rect 210660 234892 217232 234920
rect 210660 234880 210666 234892
rect 217226 234880 217232 234892
rect 217284 234880 217290 234932
rect 224926 234852 224954 234960
rect 235258 234948 235264 235000
rect 235316 234988 235322 235000
rect 294966 234988 294972 235000
rect 235316 234960 294972 234988
rect 235316 234948 235322 234960
rect 294966 234948 294972 234960
rect 295024 234948 295030 235000
rect 254026 234880 254032 234932
rect 254084 234920 254090 234932
rect 255222 234920 255228 234932
rect 254084 234892 255228 234920
rect 254084 234880 254090 234892
rect 255222 234880 255228 234892
rect 255280 234880 255286 234932
rect 245562 234852 245568 234864
rect 224926 234824 245568 234852
rect 245562 234812 245568 234824
rect 245620 234852 245626 234864
rect 245838 234852 245844 234864
rect 245620 234824 245844 234852
rect 245620 234812 245626 234824
rect 245838 234812 245844 234824
rect 245896 234812 245902 234864
rect 213546 234744 213552 234796
rect 213604 234784 213610 234796
rect 246482 234784 246488 234796
rect 213604 234756 246488 234784
rect 213604 234744 213610 234756
rect 246482 234744 246488 234756
rect 246540 234784 246546 234796
rect 246850 234784 246856 234796
rect 246540 234756 246856 234784
rect 246540 234744 246546 234756
rect 246850 234744 246856 234756
rect 246908 234744 246914 234796
rect 210786 234676 210792 234728
rect 210844 234716 210850 234728
rect 210844 234688 215294 234716
rect 210844 234676 210850 234688
rect 215266 234648 215294 234688
rect 217226 234676 217232 234728
rect 217284 234716 217290 234728
rect 247310 234716 247316 234728
rect 217284 234688 247316 234716
rect 217284 234676 217290 234688
rect 247310 234676 247316 234688
rect 247368 234716 247374 234728
rect 247770 234716 247776 234728
rect 247368 234688 247776 234716
rect 247368 234676 247374 234688
rect 247770 234676 247776 234688
rect 247828 234676 247834 234728
rect 256786 234676 256792 234728
rect 256844 234716 256850 234728
rect 257890 234716 257896 234728
rect 256844 234688 257896 234716
rect 256844 234676 256850 234688
rect 257890 234676 257896 234688
rect 257948 234676 257954 234728
rect 258442 234648 258448 234660
rect 215266 234620 258448 234648
rect 258442 234608 258448 234620
rect 258500 234608 258506 234660
rect 291102 234608 291108 234660
rect 291160 234648 291166 234660
rect 291838 234648 291844 234660
rect 291160 234620 291844 234648
rect 291160 234608 291166 234620
rect 291838 234608 291844 234620
rect 291896 234608 291902 234660
rect 214742 234540 214748 234592
rect 214800 234580 214806 234592
rect 215202 234580 215208 234592
rect 214800 234552 215208 234580
rect 214800 234540 214806 234552
rect 215202 234540 215208 234552
rect 215260 234580 215266 234592
rect 240594 234580 240600 234592
rect 215260 234552 240600 234580
rect 215260 234540 215266 234552
rect 240594 234540 240600 234552
rect 240652 234540 240658 234592
rect 244642 234540 244648 234592
rect 244700 234580 244706 234592
rect 249150 234580 249156 234592
rect 244700 234552 249156 234580
rect 244700 234540 244706 234552
rect 249150 234540 249156 234552
rect 249208 234580 249214 234592
rect 257890 234580 257896 234592
rect 249208 234552 257896 234580
rect 249208 234540 249214 234552
rect 257890 234540 257896 234552
rect 257948 234540 257954 234592
rect 260098 234540 260104 234592
rect 260156 234580 260162 234592
rect 267642 234580 267648 234592
rect 260156 234552 267648 234580
rect 260156 234540 260162 234552
rect 267642 234540 267648 234552
rect 267700 234540 267706 234592
rect 272702 234540 272708 234592
rect 272760 234580 272766 234592
rect 273162 234580 273168 234592
rect 272760 234552 273168 234580
rect 272760 234540 272766 234552
rect 273162 234540 273168 234552
rect 273220 234580 273226 234592
rect 286502 234580 286508 234592
rect 273220 234552 286508 234580
rect 273220 234540 273226 234552
rect 286502 234540 286508 234552
rect 286560 234540 286566 234592
rect 243446 234472 243452 234524
rect 243504 234512 243510 234524
rect 303062 234512 303068 234524
rect 243504 234484 303068 234512
rect 243504 234472 243510 234484
rect 303062 234472 303068 234484
rect 303120 234472 303126 234524
rect 208486 234404 208492 234456
rect 208544 234444 208550 234456
rect 209314 234444 209320 234456
rect 208544 234416 209320 234444
rect 208544 234404 208550 234416
rect 209314 234404 209320 234416
rect 209372 234444 209378 234456
rect 239030 234444 239036 234456
rect 209372 234416 239036 234444
rect 209372 234404 209378 234416
rect 239030 234404 239036 234416
rect 239088 234404 239094 234456
rect 245746 234404 245752 234456
rect 245804 234444 245810 234456
rect 300394 234444 300400 234456
rect 245804 234416 300400 234444
rect 245804 234404 245810 234416
rect 300394 234404 300400 234416
rect 300452 234404 300458 234456
rect 202322 234336 202328 234388
rect 202380 234376 202386 234388
rect 202598 234376 202604 234388
rect 202380 234348 202604 234376
rect 202380 234336 202386 234348
rect 202598 234336 202604 234348
rect 202656 234376 202662 234388
rect 228174 234376 228180 234388
rect 202656 234348 228180 234376
rect 202656 234336 202662 234348
rect 228174 234336 228180 234348
rect 228232 234336 228238 234388
rect 237558 234336 237564 234388
rect 237616 234376 237622 234388
rect 282822 234376 282828 234388
rect 237616 234348 282828 234376
rect 237616 234336 237622 234348
rect 282822 234336 282828 234348
rect 282880 234336 282886 234388
rect 244274 234308 244280 234320
rect 215266 234280 244280 234308
rect 188890 234064 188896 234116
rect 188948 234104 188954 234116
rect 214742 234104 214748 234116
rect 188948 234076 214748 234104
rect 188948 234064 188954 234076
rect 214742 234064 214748 234076
rect 214800 234064 214806 234116
rect 184842 233996 184848 234048
rect 184900 234036 184906 234048
rect 211614 234036 211620 234048
rect 184900 234008 211620 234036
rect 184900 233996 184906 234008
rect 211614 233996 211620 234008
rect 211672 234036 211678 234048
rect 215266 234036 215294 234280
rect 244274 234268 244280 234280
rect 244332 234268 244338 234320
rect 250530 234268 250536 234320
rect 250588 234308 250594 234320
rect 258718 234308 258724 234320
rect 250588 234280 258724 234308
rect 250588 234268 250594 234280
rect 258718 234268 258724 234280
rect 258776 234268 258782 234320
rect 259270 234268 259276 234320
rect 259328 234308 259334 234320
rect 306006 234308 306012 234320
rect 259328 234280 306012 234308
rect 259328 234268 259334 234280
rect 306006 234268 306012 234280
rect 306064 234268 306070 234320
rect 235258 234200 235264 234252
rect 235316 234240 235322 234252
rect 235626 234240 235632 234252
rect 235316 234212 235632 234240
rect 235316 234200 235322 234212
rect 235626 234200 235632 234212
rect 235684 234240 235690 234252
rect 276474 234240 276480 234252
rect 235684 234212 276480 234240
rect 235684 234200 235690 234212
rect 276474 234200 276480 234212
rect 276532 234200 276538 234252
rect 235350 234132 235356 234184
rect 235408 234172 235414 234184
rect 275554 234172 275560 234184
rect 235408 234144 275560 234172
rect 235408 234132 235414 234144
rect 275554 234132 275560 234144
rect 275612 234132 275618 234184
rect 239122 234064 239128 234116
rect 239180 234104 239186 234116
rect 239674 234104 239680 234116
rect 239180 234076 239680 234104
rect 239180 234064 239186 234076
rect 239674 234064 239680 234076
rect 239732 234104 239738 234116
rect 279326 234104 279332 234116
rect 239732 234076 279332 234104
rect 239732 234064 239738 234076
rect 279326 234064 279332 234076
rect 279384 234064 279390 234116
rect 211672 234008 215294 234036
rect 211672 233996 211678 234008
rect 241238 233996 241244 234048
rect 241296 234036 241302 234048
rect 242342 234036 242348 234048
rect 241296 234008 242348 234036
rect 241296 233996 241302 234008
rect 242342 233996 242348 234008
rect 242400 234036 242406 234048
rect 280798 234036 280804 234048
rect 242400 234008 280804 234036
rect 242400 233996 242406 234008
rect 280798 233996 280804 234008
rect 280856 233996 280862 234048
rect 172330 233928 172336 233980
rect 172388 233968 172394 233980
rect 202598 233968 202604 233980
rect 172388 233940 202604 233968
rect 172388 233928 172394 233940
rect 202598 233928 202604 233940
rect 202656 233928 202662 233980
rect 235166 233928 235172 233980
rect 235224 233968 235230 233980
rect 235810 233968 235816 233980
rect 235224 233940 235816 233968
rect 235224 233928 235230 233940
rect 235810 233928 235816 233940
rect 235868 233928 235874 233980
rect 250898 233968 250904 233980
rect 241624 233940 250904 233968
rect 156966 233860 156972 233912
rect 157024 233900 157030 233912
rect 208394 233900 208400 233912
rect 157024 233872 208400 233900
rect 157024 233860 157030 233872
rect 208394 233860 208400 233872
rect 208452 233860 208458 233912
rect 211890 233860 211896 233912
rect 211948 233900 211954 233912
rect 212442 233900 212448 233912
rect 211948 233872 212448 233900
rect 211948 233860 211954 233872
rect 212442 233860 212448 233872
rect 212500 233860 212506 233912
rect 216398 233860 216404 233912
rect 216456 233900 216462 233912
rect 241624 233900 241652 233940
rect 250898 233928 250904 233940
rect 250956 233928 250962 233980
rect 258718 233928 258724 233980
rect 258776 233968 258782 233980
rect 284202 233968 284208 233980
rect 258776 233940 284208 233968
rect 258776 233928 258782 233940
rect 284202 233928 284208 233940
rect 284260 233928 284266 233980
rect 216456 233872 241652 233900
rect 216456 233860 216462 233872
rect 241698 233860 241704 233912
rect 241756 233900 241762 233912
rect 242710 233900 242716 233912
rect 241756 233872 242716 233900
rect 241756 233860 241762 233872
rect 242710 233860 242716 233872
rect 242768 233860 242774 233912
rect 243722 233860 243728 233912
rect 243780 233900 243786 233912
rect 278774 233900 278780 233912
rect 243780 233872 278780 233900
rect 243780 233860 243786 233872
rect 278774 233860 278780 233872
rect 278832 233900 278838 233912
rect 280062 233900 280068 233912
rect 278832 233872 280068 233900
rect 278832 233860 278838 233872
rect 280062 233860 280068 233872
rect 280120 233860 280126 233912
rect 212460 233832 212488 233860
rect 246390 233832 246396 233844
rect 212460 233804 246396 233832
rect 246390 233792 246396 233804
rect 246448 233792 246454 233844
rect 257890 233792 257896 233844
rect 257948 233832 257954 233844
rect 284018 233832 284024 233844
rect 257948 233804 284024 233832
rect 257948 233792 257954 233804
rect 284018 233792 284024 233804
rect 284076 233792 284082 233844
rect 232866 233724 232872 233776
rect 232924 233764 232930 233776
rect 233142 233764 233148 233776
rect 232924 233736 233148 233764
rect 232924 233724 232930 233736
rect 233142 233724 233148 233736
rect 233200 233724 233206 233776
rect 239950 233724 239956 233776
rect 240008 233764 240014 233776
rect 272886 233764 272892 233776
rect 240008 233736 253934 233764
rect 240008 233724 240014 233736
rect 218698 233656 218704 233708
rect 218756 233696 218762 233708
rect 251082 233696 251088 233708
rect 218756 233668 251088 233696
rect 218756 233656 218762 233668
rect 251082 233656 251088 233668
rect 251140 233656 251146 233708
rect 253906 233696 253934 233736
rect 260806 233736 272892 233764
rect 260806 233696 260834 233736
rect 272886 233724 272892 233736
rect 272944 233724 272950 233776
rect 253906 233668 260834 233696
rect 263778 233656 263784 233708
rect 263836 233696 263842 233708
rect 264698 233696 264704 233708
rect 263836 233668 264704 233696
rect 263836 233656 263842 233668
rect 264698 233656 264704 233668
rect 264756 233656 264762 233708
rect 267642 233656 267648 233708
rect 267700 233696 267706 233708
rect 270126 233696 270132 233708
rect 267700 233668 270132 233696
rect 267700 233656 267706 233668
rect 270126 233656 270132 233668
rect 270184 233696 270190 233708
rect 278498 233696 278504 233708
rect 270184 233668 278504 233696
rect 270184 233656 270190 233668
rect 278498 233656 278504 233668
rect 278556 233656 278562 233708
rect 298922 233628 298928 233640
rect 255286 233600 298928 233628
rect 253566 233452 253572 233504
rect 253624 233492 253630 233504
rect 253842 233492 253848 233504
rect 253624 233464 253848 233492
rect 253624 233452 253630 233464
rect 253842 233452 253848 233464
rect 253900 233452 253906 233504
rect 242986 233384 242992 233436
rect 243044 233424 243050 233436
rect 243630 233424 243636 233436
rect 243044 233396 243636 233424
rect 243044 233384 243050 233396
rect 243630 233384 243636 233396
rect 243688 233384 243694 233436
rect 239582 233316 239588 233368
rect 239640 233356 239646 233368
rect 255286 233356 255314 233600
rect 298922 233588 298928 233600
rect 298980 233588 298986 233640
rect 239640 233328 255314 233356
rect 239640 233316 239646 233328
rect 226518 233248 226524 233300
rect 226576 233288 226582 233300
rect 227346 233288 227352 233300
rect 226576 233260 227352 233288
rect 226576 233248 226582 233260
rect 227346 233248 227352 233260
rect 227404 233248 227410 233300
rect 245378 233248 245384 233300
rect 245436 233288 245442 233300
rect 245746 233288 245752 233300
rect 245436 233260 245752 233288
rect 245436 233248 245442 233260
rect 245746 233248 245752 233260
rect 245804 233248 245810 233300
rect 205634 233180 205640 233232
rect 205692 233220 205698 233232
rect 206554 233220 206560 233232
rect 205692 233192 206560 233220
rect 205692 233180 205698 233192
rect 206554 233180 206560 233192
rect 206612 233220 206618 233232
rect 229002 233220 229008 233232
rect 206612 233192 229008 233220
rect 206612 233180 206618 233192
rect 229002 233180 229008 233192
rect 229060 233180 229066 233232
rect 246114 233180 246120 233232
rect 246172 233220 246178 233232
rect 246666 233220 246672 233232
rect 246172 233192 246672 233220
rect 246172 233180 246178 233192
rect 246666 233180 246672 233192
rect 246724 233180 246730 233232
rect 253474 233180 253480 233232
rect 253532 233220 253538 233232
rect 253842 233220 253848 233232
rect 253532 233192 253848 233220
rect 253532 233180 253538 233192
rect 253842 233180 253848 233192
rect 253900 233180 253906 233232
rect 254026 233180 254032 233232
rect 254084 233220 254090 233232
rect 269666 233220 269672 233232
rect 254084 233192 269672 233220
rect 254084 233180 254090 233192
rect 269666 233180 269672 233192
rect 269724 233180 269730 233232
rect 270310 233180 270316 233232
rect 270368 233220 270374 233232
rect 270586 233220 270592 233232
rect 270368 233192 270592 233220
rect 270368 233180 270374 233192
rect 270586 233180 270592 233192
rect 270644 233180 270650 233232
rect 276382 233180 276388 233232
rect 276440 233220 276446 233232
rect 579614 233220 579620 233232
rect 276440 233192 579620 233220
rect 276440 233180 276446 233192
rect 579614 233180 579620 233192
rect 579672 233180 579678 233232
rect 251082 233112 251088 233164
rect 251140 233152 251146 233164
rect 309962 233152 309968 233164
rect 251140 233124 309968 233152
rect 251140 233112 251146 233124
rect 309962 233112 309968 233124
rect 310020 233112 310026 233164
rect 236730 233044 236736 233096
rect 236788 233084 236794 233096
rect 237006 233084 237012 233096
rect 236788 233056 237012 233084
rect 236788 233044 236794 233056
rect 237006 233044 237012 233056
rect 237064 233084 237070 233096
rect 295978 233084 295984 233096
rect 237064 233056 295984 233084
rect 237064 233044 237070 233056
rect 295978 233044 295984 233056
rect 296036 233044 296042 233096
rect 246206 232976 246212 233028
rect 246264 233016 246270 233028
rect 305730 233016 305736 233028
rect 246264 232988 305736 233016
rect 246264 232976 246270 232988
rect 305730 232976 305736 232988
rect 305788 232976 305794 233028
rect 249794 232908 249800 232960
rect 249852 232948 249858 232960
rect 253198 232948 253204 232960
rect 249852 232920 253204 232948
rect 249852 232908 249858 232920
rect 253198 232908 253204 232920
rect 253256 232908 253262 232960
rect 253842 232908 253848 232960
rect 253900 232948 253906 232960
rect 296346 232948 296352 232960
rect 253900 232920 296352 232948
rect 253900 232908 253906 232920
rect 296346 232908 296352 232920
rect 296404 232908 296410 232960
rect 236730 232840 236736 232892
rect 236788 232880 236794 232892
rect 277670 232880 277676 232892
rect 236788 232852 277676 232880
rect 236788 232840 236794 232852
rect 277670 232840 277676 232852
rect 277728 232840 277734 232892
rect 250162 232772 250168 232824
rect 250220 232812 250226 232824
rect 251082 232812 251088 232824
rect 250220 232784 251088 232812
rect 250220 232772 250226 232784
rect 251082 232772 251088 232784
rect 251140 232772 251146 232824
rect 253198 232772 253204 232824
rect 253256 232812 253262 232824
rect 286410 232812 286416 232824
rect 253256 232784 286416 232812
rect 253256 232772 253262 232784
rect 286410 232772 286416 232784
rect 286468 232772 286474 232824
rect 191742 232704 191748 232756
rect 191800 232744 191806 232756
rect 216398 232744 216404 232756
rect 191800 232716 216404 232744
rect 191800 232704 191806 232716
rect 216398 232704 216404 232716
rect 216456 232704 216462 232756
rect 240778 232704 240784 232756
rect 240836 232744 240842 232756
rect 240836 232716 273852 232744
rect 240836 232704 240842 232716
rect 194410 232636 194416 232688
rect 194468 232676 194474 232688
rect 221918 232676 221924 232688
rect 194468 232648 221924 232676
rect 194468 232636 194474 232648
rect 221918 232636 221924 232648
rect 221976 232636 221982 232688
rect 244182 232636 244188 232688
rect 244240 232676 244246 232688
rect 273714 232676 273720 232688
rect 244240 232648 273720 232676
rect 244240 232636 244246 232648
rect 273714 232636 273720 232648
rect 273772 232636 273778 232688
rect 273824 232676 273852 232716
rect 276014 232704 276020 232756
rect 276072 232744 276078 232756
rect 277026 232744 277032 232756
rect 276072 232716 277032 232744
rect 276072 232704 276078 232716
rect 277026 232704 277032 232716
rect 277084 232744 277090 232756
rect 279602 232744 279608 232756
rect 277084 232716 279608 232744
rect 277084 232704 277090 232716
rect 279602 232704 279608 232716
rect 279660 232704 279666 232756
rect 281534 232704 281540 232756
rect 281592 232744 281598 232756
rect 293402 232744 293408 232756
rect 281592 232716 293408 232744
rect 281592 232704 281598 232716
rect 293402 232704 293408 232716
rect 293460 232704 293466 232756
rect 276842 232676 276848 232688
rect 273824 232648 276848 232676
rect 276842 232636 276848 232648
rect 276900 232636 276906 232688
rect 283558 232636 283564 232688
rect 283616 232676 283622 232688
rect 329926 232676 329932 232688
rect 283616 232648 329932 232676
rect 283616 232636 283622 232648
rect 329926 232636 329932 232648
rect 329984 232636 329990 232688
rect 152826 232568 152832 232620
rect 152884 232608 152890 232620
rect 205634 232608 205640 232620
rect 152884 232580 205640 232608
rect 152884 232568 152890 232580
rect 205634 232568 205640 232580
rect 205692 232568 205698 232620
rect 228542 232568 228548 232620
rect 228600 232608 228606 232620
rect 231854 232608 231860 232620
rect 228600 232580 231860 232608
rect 228600 232568 228606 232580
rect 231854 232568 231860 232580
rect 231912 232568 231918 232620
rect 237282 232568 237288 232620
rect 237340 232608 237346 232620
rect 238938 232608 238944 232620
rect 237340 232580 238944 232608
rect 237340 232568 237346 232580
rect 238938 232568 238944 232580
rect 238996 232568 239002 232620
rect 252278 232568 252284 232620
rect 252336 232608 252342 232620
rect 279694 232608 279700 232620
rect 252336 232580 279700 232608
rect 252336 232568 252342 232580
rect 279694 232568 279700 232580
rect 279752 232608 279758 232620
rect 334066 232608 334072 232620
rect 279752 232580 334072 232608
rect 279752 232568 279758 232580
rect 334066 232568 334072 232580
rect 334124 232568 334130 232620
rect 161474 232500 161480 232552
rect 161532 232540 161538 232552
rect 191650 232540 191656 232552
rect 161532 232512 191656 232540
rect 161532 232500 161538 232512
rect 191650 232500 191656 232512
rect 191708 232500 191714 232552
rect 193122 232500 193128 232552
rect 193180 232540 193186 232552
rect 252462 232540 252468 232552
rect 193180 232512 252468 232540
rect 193180 232500 193186 232512
rect 252462 232500 252468 232512
rect 252520 232540 252526 232552
rect 254026 232540 254032 232552
rect 252520 232512 254032 232540
rect 252520 232500 252526 232512
rect 254026 232500 254032 232512
rect 254084 232500 254090 232552
rect 262766 232500 262772 232552
rect 262824 232540 262830 232552
rect 276014 232540 276020 232552
rect 262824 232512 276020 232540
rect 262824 232500 262830 232512
rect 276014 232500 276020 232512
rect 276072 232500 276078 232552
rect 280246 232500 280252 232552
rect 280304 232540 280310 232552
rect 337010 232540 337016 232552
rect 280304 232512 337016 232540
rect 280304 232500 280310 232512
rect 337010 232500 337016 232512
rect 337068 232500 337074 232552
rect 248046 232432 248052 232484
rect 248104 232472 248110 232484
rect 270034 232472 270040 232484
rect 248104 232444 270040 232472
rect 248104 232432 248110 232444
rect 270034 232432 270040 232444
rect 270092 232432 270098 232484
rect 270678 232432 270684 232484
rect 270736 232472 270742 232484
rect 270954 232472 270960 232484
rect 270736 232444 270960 232472
rect 270736 232432 270742 232444
rect 270954 232432 270960 232444
rect 271012 232432 271018 232484
rect 283558 232404 283564 232416
rect 270696 232376 283564 232404
rect 265066 232296 265072 232348
rect 265124 232336 265130 232348
rect 270696 232336 270724 232376
rect 283558 232364 283564 232376
rect 283616 232364 283622 232416
rect 265124 232308 270724 232336
rect 265124 232296 265130 232308
rect 236914 232228 236920 232280
rect 236972 232268 236978 232280
rect 237098 232268 237104 232280
rect 236972 232240 237104 232268
rect 236972 232228 236978 232240
rect 237098 232228 237104 232240
rect 237156 232268 237162 232280
rect 279510 232268 279516 232280
rect 237156 232240 279516 232268
rect 237156 232228 237162 232240
rect 279510 232228 279516 232240
rect 279568 232228 279574 232280
rect 270586 232160 270592 232212
rect 270644 232200 270650 232212
rect 271598 232200 271604 232212
rect 270644 232172 271604 232200
rect 270644 232160 270650 232172
rect 271598 232160 271604 232172
rect 271656 232160 271662 232212
rect 273622 232160 273628 232212
rect 273680 232200 273686 232212
rect 274266 232200 274272 232212
rect 273680 232172 274272 232200
rect 273680 232160 273686 232172
rect 274266 232160 274272 232172
rect 274324 232160 274330 232212
rect 270034 232092 270040 232144
rect 270092 232132 270098 232144
rect 275278 232132 275284 232144
rect 270092 232104 275284 232132
rect 270092 232092 270098 232104
rect 275278 232092 275284 232104
rect 275336 232092 275342 232144
rect 233694 232024 233700 232076
rect 233752 232064 233758 232076
rect 234246 232064 234252 232076
rect 233752 232036 234252 232064
rect 233752 232024 233758 232036
rect 234246 232024 234252 232036
rect 234304 232024 234310 232076
rect 241054 231956 241060 232008
rect 241112 231996 241118 232008
rect 241330 231996 241336 232008
rect 241112 231968 241336 231996
rect 241112 231956 241118 231968
rect 241330 231956 241336 231968
rect 241388 231956 241394 232008
rect 256878 231956 256884 232008
rect 256936 231996 256942 232008
rect 261570 231996 261576 232008
rect 256936 231968 261576 231996
rect 256936 231956 256942 231968
rect 261570 231956 261576 231968
rect 261628 231956 261634 232008
rect 195882 231820 195888 231872
rect 195940 231860 195946 231872
rect 252554 231860 252560 231872
rect 195940 231832 252560 231860
rect 195940 231820 195946 231832
rect 252554 231820 252560 231832
rect 252612 231820 252618 231872
rect 255590 231820 255596 231872
rect 255648 231860 255654 231872
rect 256602 231860 256608 231872
rect 255648 231832 256608 231860
rect 255648 231820 255654 231832
rect 256602 231820 256608 231832
rect 256660 231820 256666 231872
rect 256878 231820 256884 231872
rect 256936 231860 256942 231872
rect 258074 231860 258080 231872
rect 256936 231832 258080 231860
rect 256936 231820 256942 231832
rect 258074 231820 258080 231832
rect 258132 231820 258138 231872
rect 199010 231752 199016 231804
rect 199068 231792 199074 231804
rect 200022 231792 200028 231804
rect 199068 231764 200028 231792
rect 199068 231752 199074 231764
rect 200022 231752 200028 231764
rect 200080 231792 200086 231804
rect 228726 231792 228732 231804
rect 200080 231764 228732 231792
rect 200080 231752 200086 231764
rect 228726 231752 228732 231764
rect 228784 231752 228790 231804
rect 233418 231752 233424 231804
rect 233476 231792 233482 231804
rect 234062 231792 234068 231804
rect 233476 231764 234068 231792
rect 233476 231752 233482 231764
rect 234062 231752 234068 231764
rect 234120 231792 234126 231804
rect 234120 231764 238754 231792
rect 234120 231752 234126 231764
rect 238726 231724 238754 231764
rect 262858 231752 262864 231804
rect 262916 231792 262922 231804
rect 274910 231792 274916 231804
rect 262916 231764 274916 231792
rect 262916 231752 262922 231764
rect 274910 231752 274916 231764
rect 274968 231792 274974 231804
rect 275738 231792 275744 231804
rect 274968 231764 275744 231792
rect 274968 231752 274974 231764
rect 275738 231752 275744 231764
rect 275796 231752 275802 231804
rect 276106 231752 276112 231804
rect 276164 231792 276170 231804
rect 276934 231792 276940 231804
rect 276164 231764 276940 231792
rect 276164 231752 276170 231764
rect 276934 231752 276940 231764
rect 276992 231752 276998 231804
rect 293218 231724 293224 231736
rect 238726 231696 293224 231724
rect 293218 231684 293224 231696
rect 293276 231684 293282 231736
rect 250990 231616 250996 231668
rect 251048 231656 251054 231668
rect 301774 231656 301780 231668
rect 251048 231628 301780 231656
rect 251048 231616 251054 231628
rect 301774 231616 301780 231628
rect 301832 231616 301838 231668
rect 199838 231548 199844 231600
rect 199896 231588 199902 231600
rect 259362 231588 259368 231600
rect 199896 231560 259368 231588
rect 199896 231548 199902 231560
rect 259362 231548 259368 231560
rect 259420 231548 259426 231600
rect 247402 231480 247408 231532
rect 247460 231520 247466 231532
rect 296070 231520 296076 231532
rect 247460 231492 296076 231520
rect 247460 231480 247466 231492
rect 296070 231480 296076 231492
rect 296128 231480 296134 231532
rect 232038 231412 232044 231464
rect 232096 231452 232102 231464
rect 232406 231452 232412 231464
rect 232096 231424 232412 231452
rect 232096 231412 232102 231424
rect 232406 231412 232412 231424
rect 232464 231412 232470 231464
rect 244090 231412 244096 231464
rect 244148 231452 244154 231464
rect 275462 231452 275468 231464
rect 244148 231424 275468 231452
rect 244148 231412 244154 231424
rect 275462 231412 275468 231424
rect 275520 231412 275526 231464
rect 248966 231344 248972 231396
rect 249024 231384 249030 231396
rect 280246 231384 280252 231396
rect 249024 231356 280252 231384
rect 249024 231344 249030 231356
rect 280246 231344 280252 231356
rect 280304 231344 280310 231396
rect 253566 231276 253572 231328
rect 253624 231316 253630 231328
rect 283742 231316 283748 231328
rect 253624 231288 283748 231316
rect 253624 231276 253630 231288
rect 283742 231276 283748 231288
rect 283800 231276 283806 231328
rect 152734 231208 152740 231260
rect 152792 231248 152798 231260
rect 199010 231248 199016 231260
rect 152792 231220 199016 231248
rect 152792 231208 152798 231220
rect 199010 231208 199016 231220
rect 199068 231208 199074 231260
rect 248138 231208 248144 231260
rect 248196 231248 248202 231260
rect 276106 231248 276112 231260
rect 248196 231220 276112 231248
rect 248196 231208 248202 231220
rect 276106 231208 276112 231220
rect 276164 231208 276170 231260
rect 289722 231208 289728 231260
rect 289780 231248 289786 231260
rect 332778 231248 332784 231260
rect 289780 231220 332784 231248
rect 289780 231208 289786 231220
rect 332778 231208 332784 231220
rect 332836 231208 332842 231260
rect 256418 231140 256424 231192
rect 256476 231180 256482 231192
rect 290642 231180 290648 231192
rect 256476 231152 290648 231180
rect 256476 231140 256482 231152
rect 290642 231140 290648 231152
rect 290700 231180 290706 231192
rect 336918 231180 336924 231192
rect 290700 231152 336924 231180
rect 290700 231140 290706 231152
rect 336918 231140 336924 231152
rect 336976 231140 336982 231192
rect 196986 231072 196992 231124
rect 197044 231112 197050 231124
rect 256970 231112 256976 231124
rect 197044 231084 256976 231112
rect 197044 231072 197050 231084
rect 256970 231072 256976 231084
rect 257028 231072 257034 231124
rect 261570 231072 261576 231124
rect 261628 231112 261634 231124
rect 338298 231112 338304 231124
rect 261628 231084 338304 231112
rect 261628 231072 261634 231084
rect 338298 231072 338304 231084
rect 338356 231072 338362 231124
rect 260282 231004 260288 231056
rect 260340 231044 260346 231056
rect 281534 231044 281540 231056
rect 260340 231016 281540 231044
rect 260340 231004 260346 231016
rect 281534 231004 281540 231016
rect 281592 231004 281598 231056
rect 269022 230936 269028 230988
rect 269080 230976 269086 230988
rect 289170 230976 289176 230988
rect 269080 230948 289176 230976
rect 269080 230936 269086 230948
rect 289170 230936 289176 230948
rect 289228 230976 289234 230988
rect 289722 230976 289728 230988
rect 289228 230948 289728 230976
rect 289228 230936 289234 230948
rect 289722 230936 289728 230948
rect 289780 230936 289786 230988
rect 239398 230868 239404 230920
rect 239456 230908 239462 230920
rect 298646 230908 298652 230920
rect 239456 230880 298652 230908
rect 239456 230868 239462 230880
rect 298646 230868 298652 230880
rect 298704 230868 298710 230920
rect 252922 230800 252928 230852
rect 252980 230840 252986 230852
rect 312906 230840 312912 230852
rect 252980 230812 312912 230840
rect 252980 230800 252986 230812
rect 312906 230800 312912 230812
rect 312964 230800 312970 230852
rect 247402 230732 247408 230784
rect 247460 230772 247466 230784
rect 248138 230772 248144 230784
rect 247460 230744 248144 230772
rect 247460 230732 247466 230744
rect 248138 230732 248144 230744
rect 248196 230732 248202 230784
rect 255498 230732 255504 230784
rect 255556 230772 255562 230784
rect 256510 230772 256516 230784
rect 255556 230744 256516 230772
rect 255556 230732 255562 230744
rect 256510 230732 256516 230744
rect 256568 230732 256574 230784
rect 199930 230664 199936 230716
rect 199988 230704 199994 230716
rect 259454 230704 259460 230716
rect 199988 230676 259460 230704
rect 199988 230664 199994 230676
rect 259454 230664 259460 230676
rect 259512 230664 259518 230716
rect 197170 230596 197176 230648
rect 197228 230636 197234 230648
rect 255130 230636 255136 230648
rect 197228 230608 255136 230636
rect 197228 230596 197234 230608
rect 255130 230596 255136 230608
rect 255188 230596 255194 230648
rect 259270 230636 259276 230648
rect 255424 230608 259276 230636
rect 199746 230528 199752 230580
rect 199804 230568 199810 230580
rect 255424 230568 255452 230608
rect 259270 230596 259276 230608
rect 259328 230596 259334 230648
rect 199804 230540 255452 230568
rect 199804 230528 199810 230540
rect 198642 230460 198648 230512
rect 198700 230500 198706 230512
rect 257706 230500 257712 230512
rect 198700 230472 257712 230500
rect 198700 230460 198706 230472
rect 257706 230460 257712 230472
rect 257764 230460 257770 230512
rect 271414 230500 271420 230512
rect 271064 230472 271420 230500
rect 214742 230392 214748 230444
rect 214800 230432 214806 230444
rect 216122 230432 216128 230444
rect 214800 230404 216128 230432
rect 214800 230392 214806 230404
rect 216122 230392 216128 230404
rect 216180 230392 216186 230444
rect 232774 230392 232780 230444
rect 232832 230432 232838 230444
rect 233510 230432 233516 230444
rect 232832 230404 233516 230432
rect 232832 230392 232838 230404
rect 233510 230392 233516 230404
rect 233568 230392 233574 230444
rect 244274 230392 244280 230444
rect 244332 230432 244338 230444
rect 245102 230432 245108 230444
rect 244332 230404 245108 230432
rect 244332 230392 244338 230404
rect 245102 230392 245108 230404
rect 245160 230392 245166 230444
rect 249794 230392 249800 230444
rect 249852 230432 249858 230444
rect 250438 230432 250444 230444
rect 249852 230404 250444 230432
rect 249852 230392 249858 230404
rect 250438 230392 250444 230404
rect 250496 230432 250502 230444
rect 271064 230432 271092 230472
rect 271414 230460 271420 230472
rect 271472 230460 271478 230512
rect 250496 230404 271092 230432
rect 250496 230392 250502 230404
rect 271138 230392 271144 230444
rect 271196 230432 271202 230444
rect 273438 230432 273444 230444
rect 271196 230404 273444 230432
rect 271196 230392 271202 230404
rect 273438 230392 273444 230404
rect 273496 230392 273502 230444
rect 274450 230392 274456 230444
rect 274508 230432 274514 230444
rect 275462 230432 275468 230444
rect 274508 230404 275468 230432
rect 274508 230392 274514 230404
rect 275462 230392 275468 230404
rect 275520 230392 275526 230444
rect 301590 230364 301596 230376
rect 245120 230336 301596 230364
rect 244182 230256 244188 230308
rect 244240 230296 244246 230308
rect 244274 230296 244280 230308
rect 244240 230268 244280 230296
rect 244240 230256 244246 230268
rect 244274 230256 244280 230268
rect 244332 230256 244338 230308
rect 239398 230188 239404 230240
rect 239456 230228 239462 230240
rect 240042 230228 240048 230240
rect 239456 230200 240048 230228
rect 239456 230188 239462 230200
rect 240042 230188 240048 230200
rect 240100 230228 240106 230240
rect 245120 230228 245148 230336
rect 301590 230324 301596 230336
rect 301648 230324 301654 230376
rect 245194 230256 245200 230308
rect 245252 230296 245258 230308
rect 303614 230296 303620 230308
rect 245252 230268 303620 230296
rect 245252 230256 245258 230268
rect 303614 230256 303620 230268
rect 303672 230256 303678 230308
rect 304442 230228 304448 230240
rect 240100 230200 245148 230228
rect 247006 230200 304448 230228
rect 240100 230188 240106 230200
rect 247006 230172 247034 230200
rect 304442 230188 304448 230200
rect 304500 230188 304506 230240
rect 221826 230120 221832 230172
rect 221884 230160 221890 230172
rect 243722 230160 243728 230172
rect 221884 230132 243728 230160
rect 221884 230120 221890 230132
rect 243722 230120 243728 230132
rect 243780 230120 243786 230172
rect 246942 230120 246948 230172
rect 247000 230132 247034 230172
rect 247000 230120 247006 230132
rect 249334 230120 249340 230172
rect 249392 230160 249398 230172
rect 298830 230160 298836 230172
rect 249392 230132 298836 230160
rect 249392 230120 249398 230132
rect 298830 230120 298836 230132
rect 298888 230120 298894 230172
rect 233970 230052 233976 230104
rect 234028 230092 234034 230104
rect 240410 230092 240416 230104
rect 234028 230064 240416 230092
rect 234028 230052 234034 230064
rect 240410 230052 240416 230064
rect 240468 230092 240474 230104
rect 288342 230092 288348 230104
rect 240468 230064 288348 230092
rect 240468 230052 240474 230064
rect 288342 230052 288348 230064
rect 288400 230052 288406 230104
rect 215202 229984 215208 230036
rect 215260 230024 215266 230036
rect 240502 230024 240508 230036
rect 215260 229996 240508 230024
rect 215260 229984 215266 229996
rect 240502 229984 240508 229996
rect 240560 230024 240566 230036
rect 280982 230024 280988 230036
rect 240560 229996 280988 230024
rect 240560 229984 240566 229996
rect 280982 229984 280988 229996
rect 281040 229984 281046 230036
rect 212442 229916 212448 229968
rect 212500 229956 212506 229968
rect 239950 229956 239956 229968
rect 212500 229928 239956 229956
rect 212500 229916 212506 229928
rect 239950 229916 239956 229928
rect 240008 229916 240014 229968
rect 242618 229916 242624 229968
rect 242676 229956 242682 229968
rect 282270 229956 282276 229968
rect 242676 229928 282276 229956
rect 242676 229916 242682 229928
rect 282270 229916 282276 229928
rect 282328 229916 282334 229968
rect 212258 229848 212264 229900
rect 212316 229888 212322 229900
rect 239122 229888 239128 229900
rect 212316 229860 239128 229888
rect 212316 229848 212322 229860
rect 239122 229848 239128 229860
rect 239180 229848 239186 229900
rect 244826 229848 244832 229900
rect 244884 229888 244890 229900
rect 245194 229888 245200 229900
rect 244884 229860 245200 229888
rect 244884 229848 244890 229860
rect 245194 229848 245200 229860
rect 245252 229848 245258 229900
rect 246206 229848 246212 229900
rect 246264 229888 246270 229900
rect 246574 229888 246580 229900
rect 246264 229860 246580 229888
rect 246264 229848 246270 229860
rect 246574 229848 246580 229860
rect 246632 229888 246638 229900
rect 269298 229888 269304 229900
rect 246632 229860 269304 229888
rect 246632 229848 246638 229860
rect 269298 229848 269304 229860
rect 269356 229848 269362 229900
rect 269390 229848 269396 229900
rect 269448 229888 269454 229900
rect 276750 229888 276756 229900
rect 269448 229860 276756 229888
rect 269448 229848 269454 229860
rect 276750 229848 276756 229860
rect 276808 229848 276814 229900
rect 223574 229780 223580 229832
rect 223632 229820 223638 229832
rect 224862 229820 224868 229832
rect 223632 229792 224868 229820
rect 223632 229780 223638 229792
rect 224862 229780 224868 229792
rect 224920 229780 224926 229832
rect 233510 229780 233516 229832
rect 233568 229820 233574 229832
rect 278314 229820 278320 229832
rect 233568 229792 278320 229820
rect 233568 229780 233574 229792
rect 278314 229780 278320 229792
rect 278372 229780 278378 229832
rect 218698 229712 218704 229764
rect 218756 229752 218762 229764
rect 234890 229752 234896 229764
rect 218756 229724 234896 229752
rect 218756 229712 218762 229724
rect 234890 229712 234896 229724
rect 234948 229712 234954 229764
rect 238726 229724 241652 229752
rect 223758 229644 223764 229696
rect 223816 229684 223822 229696
rect 224034 229684 224040 229696
rect 223816 229656 224040 229684
rect 223816 229644 223822 229656
rect 224034 229644 224040 229656
rect 224092 229644 224098 229696
rect 228726 229644 228732 229696
rect 228784 229684 228790 229696
rect 238726 229684 238754 229724
rect 228784 229656 238754 229684
rect 241624 229684 241652 229724
rect 244642 229712 244648 229764
rect 244700 229752 244706 229764
rect 245470 229752 245476 229764
rect 244700 229724 245476 229752
rect 244700 229712 244706 229724
rect 245470 229712 245476 229724
rect 245528 229712 245534 229764
rect 246022 229712 246028 229764
rect 246080 229752 246086 229764
rect 246574 229752 246580 229764
rect 246080 229724 246580 229752
rect 246080 229712 246086 229724
rect 246574 229712 246580 229724
rect 246632 229712 246638 229764
rect 248414 229712 248420 229764
rect 248472 229752 248478 229764
rect 249518 229752 249524 229764
rect 248472 229724 249524 229752
rect 248472 229712 248478 229724
rect 249518 229712 249524 229724
rect 249576 229712 249582 229764
rect 251266 229712 251272 229764
rect 251324 229752 251330 229764
rect 252370 229752 252376 229764
rect 251324 229724 252376 229752
rect 251324 229712 251330 229724
rect 252370 229712 252376 229724
rect 252428 229712 252434 229764
rect 252554 229712 252560 229764
rect 252612 229752 252618 229764
rect 253750 229752 253756 229764
rect 252612 229724 253756 229752
rect 252612 229712 252618 229724
rect 253750 229712 253756 229724
rect 253808 229712 253814 229764
rect 254026 229712 254032 229764
rect 254084 229752 254090 229764
rect 254946 229752 254952 229764
rect 254084 229724 254952 229752
rect 254084 229712 254090 229724
rect 254946 229712 254952 229724
rect 255004 229712 255010 229764
rect 255498 229712 255504 229764
rect 255556 229752 255562 229764
rect 256326 229752 256332 229764
rect 255556 229724 256332 229752
rect 255556 229712 255562 229724
rect 256326 229712 256332 229724
rect 256384 229712 256390 229764
rect 265526 229712 265532 229764
rect 265584 229752 265590 229764
rect 285030 229752 285036 229764
rect 265584 229724 285036 229752
rect 265584 229712 265590 229724
rect 285030 229712 285036 229724
rect 285088 229752 285094 229764
rect 335446 229752 335452 229764
rect 285088 229724 335452 229752
rect 285088 229712 285094 229724
rect 335446 229712 335452 229724
rect 335504 229712 335510 229764
rect 249794 229684 249800 229696
rect 241624 229656 249800 229684
rect 228784 229644 228790 229656
rect 249794 229644 249800 229656
rect 249852 229644 249858 229696
rect 254302 229644 254308 229696
rect 254360 229684 254366 229696
rect 254578 229684 254584 229696
rect 254360 229656 254584 229684
rect 254360 229644 254366 229656
rect 254578 229644 254584 229656
rect 254636 229644 254642 229696
rect 269298 229644 269304 229696
rect 269356 229684 269362 229696
rect 272978 229684 272984 229696
rect 269356 229656 272984 229684
rect 269356 229644 269362 229656
rect 272978 229644 272984 229656
rect 273036 229644 273042 229696
rect 227162 229576 227168 229628
rect 227220 229616 227226 229628
rect 241514 229616 241520 229628
rect 227220 229588 241520 229616
rect 227220 229576 227226 229588
rect 241514 229576 241520 229588
rect 241572 229576 241578 229628
rect 241606 229576 241612 229628
rect 241664 229616 241670 229628
rect 242158 229616 242164 229628
rect 241664 229588 242164 229616
rect 241664 229576 241670 229588
rect 242158 229576 242164 229588
rect 242216 229576 242222 229628
rect 245470 229576 245476 229628
rect 245528 229616 245534 229628
rect 249334 229616 249340 229628
rect 245528 229588 249340 229616
rect 245528 229576 245534 229588
rect 249334 229576 249340 229588
rect 249392 229576 249398 229628
rect 253566 229576 253572 229628
rect 253624 229616 253630 229628
rect 253750 229616 253756 229628
rect 253624 229588 253756 229616
rect 253624 229576 253630 229588
rect 253750 229576 253756 229588
rect 253808 229576 253814 229628
rect 259822 229576 259828 229628
rect 259880 229616 259886 229628
rect 260834 229616 260840 229628
rect 259880 229588 260840 229616
rect 259880 229576 259886 229588
rect 260834 229576 260840 229588
rect 260892 229576 260898 229628
rect 223758 229508 223764 229560
rect 223816 229548 223822 229560
rect 224218 229548 224224 229560
rect 223816 229520 224224 229548
rect 223816 229508 223822 229520
rect 224218 229508 224224 229520
rect 224276 229508 224282 229560
rect 239582 229508 239588 229560
rect 239640 229548 239646 229560
rect 256142 229548 256148 229560
rect 239640 229520 256148 229548
rect 239640 229508 239646 229520
rect 256142 229508 256148 229520
rect 256200 229508 256206 229560
rect 222102 229440 222108 229492
rect 222160 229480 222166 229492
rect 302878 229480 302884 229492
rect 222160 229452 302884 229480
rect 222160 229440 222166 229452
rect 302878 229440 302884 229452
rect 302936 229440 302942 229492
rect 201218 229372 201224 229424
rect 201276 229412 201282 229424
rect 271966 229412 271972 229424
rect 201276 229384 271972 229412
rect 201276 229372 201282 229384
rect 271966 229372 271972 229384
rect 272024 229372 272030 229424
rect 241514 229304 241520 229356
rect 241572 229344 241578 229356
rect 248322 229344 248328 229356
rect 241572 229316 248328 229344
rect 241572 229304 241578 229316
rect 248322 229304 248328 229316
rect 248380 229304 248386 229356
rect 223298 229100 223304 229152
rect 223356 229140 223362 229152
rect 244182 229140 244188 229152
rect 223356 229112 244188 229140
rect 223356 229100 223362 229112
rect 244182 229100 244188 229112
rect 244240 229100 244246 229152
rect 208210 229032 208216 229084
rect 208268 229072 208274 229084
rect 226610 229072 226616 229084
rect 208268 229044 226616 229072
rect 208268 229032 208274 229044
rect 226610 229032 226616 229044
rect 226668 229032 226674 229084
rect 237282 229032 237288 229084
rect 237340 229072 237346 229084
rect 298738 229072 298744 229084
rect 237340 229044 298744 229072
rect 237340 229032 237346 229044
rect 298738 229032 298744 229044
rect 298796 229032 298802 229084
rect 161566 228964 161572 229016
rect 161624 229004 161630 229016
rect 207842 229004 207848 229016
rect 161624 228976 207848 229004
rect 161624 228964 161630 228976
rect 207842 228964 207848 228976
rect 207900 228964 207906 229016
rect 226058 229004 226064 229016
rect 209746 228976 226064 229004
rect 156690 228896 156696 228948
rect 156748 228936 156754 228948
rect 208118 228936 208124 228948
rect 156748 228908 208124 228936
rect 156748 228896 156754 228908
rect 208118 228896 208124 228908
rect 208176 228936 208182 228948
rect 209746 228936 209774 228976
rect 226058 228964 226064 228976
rect 226116 228964 226122 229016
rect 263778 228964 263784 229016
rect 263836 229004 263842 229016
rect 325142 229004 325148 229016
rect 263836 228976 325148 229004
rect 263836 228964 263842 228976
rect 325142 228964 325148 228976
rect 325200 228964 325206 229016
rect 208176 228908 209774 228936
rect 208176 228896 208182 228908
rect 210878 228896 210884 228948
rect 210936 228936 210942 228948
rect 237466 228936 237472 228948
rect 210936 228908 237472 228936
rect 210936 228896 210942 228908
rect 237466 228896 237472 228908
rect 237524 228896 237530 228948
rect 262306 228896 262312 228948
rect 262364 228936 262370 228948
rect 323670 228936 323676 228948
rect 262364 228908 323676 228936
rect 262364 228896 262370 228908
rect 323670 228896 323676 228908
rect 323728 228896 323734 228948
rect 156782 228828 156788 228880
rect 156840 228868 156846 228880
rect 208210 228868 208216 228880
rect 156840 228840 208216 228868
rect 156840 228828 156846 228840
rect 208210 228828 208216 228840
rect 208268 228828 208274 228880
rect 211062 228828 211068 228880
rect 211120 228868 211126 228880
rect 237282 228868 237288 228880
rect 211120 228840 237288 228868
rect 211120 228828 211126 228840
rect 237282 228828 237288 228840
rect 237340 228828 237346 228880
rect 264422 228828 264428 228880
rect 264480 228868 264486 228880
rect 264790 228868 264796 228880
rect 264480 228840 264796 228868
rect 264480 228828 264486 228840
rect 264790 228828 264796 228840
rect 264848 228868 264854 228880
rect 325050 228868 325056 228880
rect 264848 228840 325056 228868
rect 264848 228828 264854 228840
rect 325050 228828 325056 228840
rect 325108 228828 325114 228880
rect 156874 228760 156880 228812
rect 156932 228800 156938 228812
rect 210970 228800 210976 228812
rect 156932 228772 210976 228800
rect 156932 228760 156938 228772
rect 210970 228760 210976 228772
rect 211028 228760 211034 228812
rect 235534 228760 235540 228812
rect 235592 228800 235598 228812
rect 294414 228800 294420 228812
rect 235592 228772 294420 228800
rect 235592 228760 235598 228772
rect 294414 228760 294420 228772
rect 294472 228760 294478 228812
rect 159634 228692 159640 228744
rect 159692 228732 159698 228744
rect 214926 228732 214932 228744
rect 159692 228704 214932 228732
rect 159692 228692 159698 228704
rect 214926 228692 214932 228704
rect 214984 228692 214990 228744
rect 217778 228692 217784 228744
rect 217836 228732 217842 228744
rect 240778 228732 240784 228744
rect 217836 228704 240784 228732
rect 217836 228692 217842 228704
rect 240778 228692 240784 228704
rect 240836 228692 240842 228744
rect 264514 228692 264520 228744
rect 264572 228732 264578 228744
rect 323762 228732 323768 228744
rect 264572 228704 323768 228732
rect 264572 228692 264578 228704
rect 323762 228692 323768 228704
rect 323820 228692 323826 228744
rect 202322 228624 202328 228676
rect 202380 228664 202386 228676
rect 270494 228664 270500 228676
rect 202380 228636 270500 228664
rect 202380 228624 202386 228636
rect 270494 228624 270500 228636
rect 270552 228624 270558 228676
rect 200206 228556 200212 228608
rect 200264 228596 200270 228608
rect 270770 228596 270776 228608
rect 200264 228568 270776 228596
rect 200264 228556 200270 228568
rect 270770 228556 270776 228568
rect 270828 228556 270834 228608
rect 197906 228488 197912 228540
rect 197964 228528 197970 228540
rect 272150 228528 272156 228540
rect 197964 228500 272156 228528
rect 197964 228488 197970 228500
rect 272150 228488 272156 228500
rect 272208 228488 272214 228540
rect 159726 228420 159732 228472
rect 159784 228460 159790 228472
rect 234798 228460 234804 228472
rect 159784 228432 234804 228460
rect 159784 228420 159790 228432
rect 234798 228420 234804 228432
rect 234856 228420 234862 228472
rect 236546 228420 236552 228472
rect 236604 228460 236610 228472
rect 237650 228460 237656 228472
rect 236604 228432 237656 228460
rect 236604 228420 236610 228432
rect 237650 228420 237656 228432
rect 237708 228460 237714 228472
rect 297450 228460 297456 228472
rect 237708 228432 297456 228460
rect 237708 228420 237714 228432
rect 297450 228420 297456 228432
rect 297508 228420 297514 228472
rect 162026 228352 162032 228404
rect 162084 228392 162090 228404
rect 239674 228392 239680 228404
rect 162084 228364 239680 228392
rect 162084 228352 162090 228364
rect 239674 228352 239680 228364
rect 239732 228352 239738 228404
rect 260006 228352 260012 228404
rect 260064 228392 260070 228404
rect 319438 228392 319444 228404
rect 260064 228364 319444 228392
rect 260064 228352 260070 228364
rect 319438 228352 319444 228364
rect 319496 228352 319502 228404
rect 235166 228284 235172 228336
rect 235224 228324 235230 228336
rect 291930 228324 291936 228336
rect 235224 228296 291936 228324
rect 235224 228284 235230 228296
rect 291930 228284 291936 228296
rect 291988 228284 291994 228336
rect 236454 228216 236460 228268
rect 236512 228256 236518 228268
rect 288158 228256 288164 228268
rect 236512 228228 288164 228256
rect 236512 228216 236518 228228
rect 288158 228216 288164 228228
rect 288216 228216 288222 228268
rect 245010 228148 245016 228200
rect 245068 228188 245074 228200
rect 269298 228188 269304 228200
rect 245068 228160 269304 228188
rect 245068 228148 245074 228160
rect 269298 228148 269304 228160
rect 269356 228148 269362 228200
rect 227714 227808 227720 227860
rect 227772 227848 227778 227860
rect 228634 227848 228640 227860
rect 227772 227820 228640 227848
rect 227772 227808 227778 227820
rect 228634 227808 228640 227820
rect 228692 227808 228698 227860
rect 263778 227808 263784 227860
rect 263836 227848 263842 227860
rect 264238 227848 264244 227860
rect 263836 227820 264244 227848
rect 263836 227808 263842 227820
rect 264238 227808 264244 227820
rect 264296 227808 264302 227860
rect 235166 227740 235172 227792
rect 235224 227780 235230 227792
rect 235626 227780 235632 227792
rect 235224 227752 235632 227780
rect 235224 227740 235230 227752
rect 235626 227740 235632 227752
rect 235684 227740 235690 227792
rect 261754 227672 261760 227724
rect 261812 227712 261818 227724
rect 271322 227712 271328 227724
rect 261812 227684 271328 227712
rect 261812 227672 261818 227684
rect 271322 227672 271328 227684
rect 271380 227672 271386 227724
rect 238110 227604 238116 227656
rect 238168 227644 238174 227656
rect 260006 227644 260012 227656
rect 238168 227616 260012 227644
rect 238168 227604 238174 227616
rect 260006 227604 260012 227616
rect 260064 227604 260070 227656
rect 231118 227536 231124 227588
rect 231176 227576 231182 227588
rect 244458 227576 244464 227588
rect 231176 227548 244464 227576
rect 231176 227536 231182 227548
rect 244458 227536 244464 227548
rect 244516 227536 244522 227588
rect 252094 227536 252100 227588
rect 252152 227576 252158 227588
rect 312998 227576 313004 227588
rect 252152 227548 313004 227576
rect 252152 227536 252158 227548
rect 312998 227536 313004 227548
rect 313056 227536 313062 227588
rect 239674 227468 239680 227520
rect 239732 227508 239738 227520
rect 259914 227508 259920 227520
rect 239732 227480 259920 227508
rect 239732 227468 239738 227480
rect 259914 227468 259920 227480
rect 259972 227468 259978 227520
rect 260558 227468 260564 227520
rect 260616 227508 260622 227520
rect 321094 227508 321100 227520
rect 260616 227480 321100 227508
rect 260616 227468 260622 227480
rect 321094 227468 321100 227480
rect 321152 227468 321158 227520
rect 234154 227400 234160 227452
rect 234212 227440 234218 227452
rect 282638 227440 282644 227452
rect 234212 227412 282644 227440
rect 234212 227400 234218 227412
rect 282638 227400 282644 227412
rect 282696 227400 282702 227452
rect 228450 227332 228456 227384
rect 228508 227372 228514 227384
rect 248966 227372 248972 227384
rect 228508 227344 248972 227372
rect 228508 227332 228514 227344
rect 248966 227332 248972 227344
rect 249024 227332 249030 227384
rect 256694 227332 256700 227384
rect 256752 227372 256758 227384
rect 304350 227372 304356 227384
rect 256752 227344 304356 227372
rect 256752 227332 256758 227344
rect 304350 227332 304356 227344
rect 304408 227332 304414 227384
rect 238570 227264 238576 227316
rect 238628 227304 238634 227316
rect 262950 227304 262956 227316
rect 238628 227276 262956 227304
rect 238628 227264 238634 227276
rect 262950 227264 262956 227276
rect 263008 227264 263014 227316
rect 223206 227196 223212 227248
rect 223264 227236 223270 227248
rect 249334 227236 249340 227248
rect 223264 227208 249340 227236
rect 223264 227196 223270 227208
rect 249334 227196 249340 227208
rect 249392 227196 249398 227248
rect 258258 227196 258264 227248
rect 258316 227236 258322 227248
rect 292574 227236 292580 227248
rect 258316 227208 292580 227236
rect 258316 227196 258322 227208
rect 292574 227196 292580 227208
rect 292632 227196 292638 227248
rect 161658 227128 161664 227180
rect 161716 227168 161722 227180
rect 207750 227168 207756 227180
rect 161716 227140 207756 227168
rect 161716 227128 161722 227140
rect 207750 227128 207756 227140
rect 207808 227128 207814 227180
rect 223114 227128 223120 227180
rect 223172 227168 223178 227180
rect 237374 227168 237380 227180
rect 223172 227140 237380 227168
rect 223172 227128 223178 227140
rect 237374 227128 237380 227140
rect 237432 227128 237438 227180
rect 238478 227128 238484 227180
rect 238536 227168 238542 227180
rect 265158 227168 265164 227180
rect 238536 227140 265164 227168
rect 238536 227128 238542 227140
rect 265158 227128 265164 227140
rect 265216 227128 265222 227180
rect 291746 227128 291752 227180
rect 291804 227168 291810 227180
rect 292206 227168 292212 227180
rect 291804 227140 292212 227168
rect 291804 227128 291810 227140
rect 292206 227128 292212 227140
rect 292264 227168 292270 227180
rect 328546 227168 328552 227180
rect 292264 227140 328552 227168
rect 292264 227128 292270 227140
rect 328546 227128 328552 227140
rect 328604 227128 328610 227180
rect 161014 227060 161020 227112
rect 161072 227100 161078 227112
rect 236914 227100 236920 227112
rect 161072 227072 236920 227100
rect 161072 227060 161078 227072
rect 236914 227060 236920 227072
rect 236972 227060 236978 227112
rect 263502 227060 263508 227112
rect 263560 227100 263566 227112
rect 291930 227100 291936 227112
rect 263560 227072 291936 227100
rect 263560 227060 263566 227072
rect 291930 227060 291936 227072
rect 291988 227100 291994 227112
rect 335354 227100 335360 227112
rect 291988 227072 335360 227100
rect 291988 227060 291994 227072
rect 335354 227060 335360 227072
rect 335412 227060 335418 227112
rect 160922 226992 160928 227044
rect 160980 227032 160986 227044
rect 236546 227032 236552 227044
rect 160980 227004 236552 227032
rect 160980 226992 160986 227004
rect 236546 226992 236552 227004
rect 236604 226992 236610 227044
rect 257614 226992 257620 227044
rect 257672 227032 257678 227044
rect 291746 227032 291752 227044
rect 257672 227004 291752 227032
rect 257672 226992 257678 227004
rect 291746 226992 291752 227004
rect 291804 226992 291810 227044
rect 292574 226992 292580 227044
rect 292632 227032 292638 227044
rect 293218 227032 293224 227044
rect 292632 227004 293224 227032
rect 292632 226992 292638 227004
rect 293218 226992 293224 227004
rect 293276 227032 293282 227044
rect 338114 227032 338120 227044
rect 293276 227004 338120 227032
rect 293276 226992 293282 227004
rect 338114 226992 338120 227004
rect 338172 226992 338178 227044
rect 224402 226924 224408 226976
rect 224460 226964 224466 226976
rect 224586 226964 224592 226976
rect 224460 226936 224592 226964
rect 224460 226924 224466 226936
rect 224586 226924 224592 226936
rect 224644 226924 224650 226976
rect 239766 226924 239772 226976
rect 239824 226964 239830 226976
rect 259638 226964 259644 226976
rect 239824 226936 259644 226964
rect 239824 226924 239830 226936
rect 259638 226924 259644 226936
rect 259696 226924 259702 226976
rect 237006 226856 237012 226908
rect 237064 226896 237070 226908
rect 259730 226896 259736 226908
rect 237064 226868 259736 226896
rect 237064 226856 237070 226868
rect 259730 226856 259736 226868
rect 259788 226856 259794 226908
rect 260926 226896 260932 226908
rect 260024 226868 260932 226896
rect 240870 226788 240876 226840
rect 240928 226828 240934 226840
rect 260024 226828 260052 226868
rect 260926 226856 260932 226868
rect 260984 226896 260990 226908
rect 260984 226868 263594 226896
rect 260984 226856 260990 226868
rect 240928 226800 260052 226828
rect 263566 226828 263594 226868
rect 338206 226828 338212 226840
rect 263566 226800 338212 226828
rect 240928 226788 240934 226800
rect 338206 226788 338212 226800
rect 338264 226788 338270 226840
rect 248690 226720 248696 226772
rect 248748 226760 248754 226772
rect 249610 226760 249616 226772
rect 248748 226732 249616 226760
rect 248748 226720 248754 226732
rect 249610 226720 249616 226732
rect 249668 226720 249674 226772
rect 262398 226720 262404 226772
rect 262456 226760 262462 226772
rect 339586 226760 339592 226772
rect 262456 226732 339592 226760
rect 262456 226720 262462 226732
rect 339586 226720 339592 226732
rect 339644 226720 339650 226772
rect 270770 226312 270776 226364
rect 270828 226352 270834 226364
rect 271322 226352 271328 226364
rect 270828 226324 271328 226352
rect 270828 226312 270834 226324
rect 271322 226312 271328 226324
rect 271380 226312 271386 226364
rect 241882 226244 241888 226296
rect 241940 226284 241946 226296
rect 327350 226284 327356 226296
rect 241940 226256 327356 226284
rect 241940 226244 241946 226256
rect 327350 226244 327356 226256
rect 327408 226244 327414 226296
rect 239030 226176 239036 226228
rect 239088 226216 239094 226228
rect 239214 226216 239220 226228
rect 239088 226188 239220 226216
rect 239088 226176 239094 226188
rect 239214 226176 239220 226188
rect 239272 226216 239278 226228
rect 300210 226216 300216 226228
rect 239272 226188 300216 226216
rect 239272 226176 239278 226188
rect 300210 226176 300216 226188
rect 300268 226176 300274 226228
rect 246482 226108 246488 226160
rect 246540 226148 246546 226160
rect 246758 226148 246764 226160
rect 246540 226120 246764 226148
rect 246540 226108 246546 226120
rect 246758 226108 246764 226120
rect 246816 226108 246822 226160
rect 251818 226108 251824 226160
rect 251876 226148 251882 226160
rect 311342 226148 311348 226160
rect 251876 226120 311348 226148
rect 251876 226108 251882 226120
rect 311342 226108 311348 226120
rect 311400 226108 311406 226160
rect 246850 226040 246856 226092
rect 246908 226080 246914 226092
rect 305638 226080 305644 226092
rect 246908 226052 305644 226080
rect 246908 226040 246914 226052
rect 305638 226040 305644 226052
rect 305696 226040 305702 226092
rect 247770 225972 247776 226024
rect 247828 226012 247834 226024
rect 307018 226012 307024 226024
rect 247828 225984 307024 226012
rect 247828 225972 247834 225984
rect 307018 225972 307024 225984
rect 307076 225972 307082 226024
rect 243078 225904 243084 225956
rect 243136 225944 243142 225956
rect 301498 225944 301504 225956
rect 243136 225916 301504 225944
rect 243136 225904 243142 225916
rect 301498 225904 301504 225916
rect 301556 225904 301562 225956
rect 246114 225836 246120 225888
rect 246172 225876 246178 225888
rect 246850 225876 246856 225888
rect 246172 225848 246856 225876
rect 246172 225836 246178 225848
rect 246850 225836 246856 225848
rect 246908 225836 246914 225888
rect 259270 225836 259276 225888
rect 259328 225876 259334 225888
rect 314102 225876 314108 225888
rect 259328 225848 314108 225876
rect 259328 225836 259334 225848
rect 314102 225836 314108 225848
rect 314160 225836 314166 225888
rect 222010 225768 222016 225820
rect 222068 225808 222074 225820
rect 239030 225808 239036 225820
rect 222068 225780 239036 225808
rect 222068 225768 222074 225780
rect 239030 225768 239036 225780
rect 239088 225768 239094 225820
rect 245562 225768 245568 225820
rect 245620 225808 245626 225820
rect 299566 225808 299572 225820
rect 245620 225780 299572 225808
rect 245620 225768 245626 225780
rect 299566 225768 299572 225780
rect 299624 225808 299630 225820
rect 300578 225808 300584 225820
rect 299624 225780 300584 225808
rect 299624 225768 299630 225780
rect 300578 225768 300584 225780
rect 300636 225768 300642 225820
rect 163498 225700 163504 225752
rect 163556 225740 163562 225752
rect 232038 225740 232044 225752
rect 163556 225712 232044 225740
rect 163556 225700 163562 225712
rect 232038 225700 232044 225712
rect 232096 225700 232102 225752
rect 244182 225700 244188 225752
rect 244240 225740 244246 225752
rect 296714 225740 296720 225752
rect 244240 225712 296720 225740
rect 244240 225700 244246 225712
rect 296714 225700 296720 225712
rect 296772 225740 296778 225752
rect 297726 225740 297732 225752
rect 296772 225712 297732 225740
rect 296772 225700 296778 225712
rect 297726 225700 297732 225712
rect 297784 225700 297790 225752
rect 154206 225632 154212 225684
rect 154264 225672 154270 225684
rect 229922 225672 229928 225684
rect 154264 225644 229928 225672
rect 154264 225632 154270 225644
rect 229922 225632 229928 225644
rect 229980 225632 229986 225684
rect 246482 225632 246488 225684
rect 246540 225672 246546 225684
rect 305914 225672 305920 225684
rect 246540 225644 305920 225672
rect 246540 225632 246546 225644
rect 305914 225632 305920 225644
rect 305972 225632 305978 225684
rect 160830 225564 160836 225616
rect 160888 225604 160894 225616
rect 236454 225604 236460 225616
rect 160888 225576 236460 225604
rect 160888 225564 160894 225576
rect 236454 225564 236460 225576
rect 236512 225564 236518 225616
rect 260926 225564 260932 225616
rect 260984 225604 260990 225616
rect 327442 225604 327448 225616
rect 260984 225576 327448 225604
rect 260984 225564 260990 225576
rect 327442 225564 327448 225576
rect 327500 225564 327506 225616
rect 241790 225496 241796 225548
rect 241848 225536 241854 225548
rect 292390 225536 292396 225548
rect 241848 225508 292396 225536
rect 241848 225496 241854 225508
rect 292390 225496 292396 225508
rect 292448 225496 292454 225548
rect 241882 225428 241888 225480
rect 241940 225468 241946 225480
rect 242526 225468 242532 225480
rect 241940 225440 242532 225468
rect 241940 225428 241946 225440
rect 242526 225428 242532 225440
rect 242584 225428 242590 225480
rect 243078 225428 243084 225480
rect 243136 225468 243142 225480
rect 243538 225468 243544 225480
rect 243136 225440 243544 225468
rect 243136 225428 243142 225440
rect 243538 225428 243544 225440
rect 243596 225428 243602 225480
rect 289262 225468 289268 225480
rect 244246 225440 289268 225468
rect 242618 225360 242624 225412
rect 242676 225400 242682 225412
rect 244246 225400 244274 225440
rect 289262 225428 289268 225440
rect 289320 225428 289326 225480
rect 242676 225372 244274 225400
rect 242676 225360 242682 225372
rect 267090 225360 267096 225412
rect 267148 225400 267154 225412
rect 267366 225400 267372 225412
rect 267148 225372 267372 225400
rect 267148 225360 267154 225372
rect 267366 225360 267372 225372
rect 267424 225360 267430 225412
rect 241698 224952 241704 225004
rect 241756 224992 241762 225004
rect 242618 224992 242624 225004
rect 241756 224964 242624 224992
rect 241756 224952 241762 224964
rect 242618 224952 242624 224964
rect 242676 224952 242682 225004
rect 260190 224884 260196 224936
rect 260248 224924 260254 224936
rect 262398 224924 262404 224936
rect 260248 224896 262404 224924
rect 260248 224884 260254 224896
rect 262398 224884 262404 224896
rect 262456 224884 262462 224936
rect 263042 224884 263048 224936
rect 263100 224924 263106 224936
rect 273438 224924 273444 224936
rect 263100 224896 273444 224924
rect 263100 224884 263106 224896
rect 273438 224884 273444 224896
rect 273496 224924 273502 224936
rect 273898 224924 273904 224936
rect 273496 224896 273904 224924
rect 273496 224884 273502 224896
rect 273898 224884 273904 224896
rect 273956 224884 273962 224936
rect 310054 224856 310060 224868
rect 249444 224828 310060 224856
rect 249444 224800 249472 224828
rect 310054 224816 310060 224828
rect 310112 224816 310118 224868
rect 248690 224748 248696 224800
rect 248748 224788 248754 224800
rect 249426 224788 249432 224800
rect 248748 224760 249432 224788
rect 248748 224748 248754 224760
rect 249426 224748 249432 224760
rect 249484 224748 249490 224800
rect 252002 224748 252008 224800
rect 252060 224788 252066 224800
rect 252370 224788 252376 224800
rect 252060 224760 252376 224788
rect 252060 224748 252066 224760
rect 252370 224748 252376 224760
rect 252428 224788 252434 224800
rect 311526 224788 311532 224800
rect 252428 224760 311532 224788
rect 252428 224748 252434 224760
rect 311526 224748 311532 224760
rect 311584 224748 311590 224800
rect 232498 224680 232504 224732
rect 232556 224720 232562 224732
rect 292022 224720 292028 224732
rect 232556 224692 292028 224720
rect 232556 224680 232562 224692
rect 292022 224680 292028 224692
rect 292080 224680 292086 224732
rect 232682 224612 232688 224664
rect 232740 224652 232746 224664
rect 238294 224652 238300 224664
rect 232740 224624 238300 224652
rect 232740 224612 232746 224624
rect 238294 224612 238300 224624
rect 238352 224652 238358 224664
rect 297358 224652 297364 224664
rect 238352 224624 297364 224652
rect 238352 224612 238358 224624
rect 297358 224612 297364 224624
rect 297416 224612 297422 224664
rect 238386 224544 238392 224596
rect 238444 224584 238450 224596
rect 296162 224584 296168 224596
rect 238444 224556 296168 224584
rect 238444 224544 238450 224556
rect 296162 224544 296168 224556
rect 296220 224544 296226 224596
rect 240042 224476 240048 224528
rect 240100 224516 240106 224528
rect 294690 224516 294696 224528
rect 240100 224488 294696 224516
rect 240100 224476 240106 224488
rect 294690 224476 294696 224488
rect 294748 224476 294754 224528
rect 240778 224408 240784 224460
rect 240836 224448 240842 224460
rect 241422 224448 241428 224460
rect 240836 224420 241428 224448
rect 240836 224408 240842 224420
rect 241422 224408 241428 224420
rect 241480 224448 241486 224460
rect 288066 224448 288072 224460
rect 241480 224420 288072 224448
rect 241480 224408 241486 224420
rect 288066 224408 288072 224420
rect 288124 224408 288130 224460
rect 240962 224340 240968 224392
rect 241020 224380 241026 224392
rect 282362 224380 282368 224392
rect 241020 224352 282368 224380
rect 241020 224340 241026 224352
rect 282362 224340 282368 224352
rect 282420 224340 282426 224392
rect 233694 224272 233700 224324
rect 233752 224312 233758 224324
rect 273990 224312 273996 224324
rect 233752 224284 273996 224312
rect 233752 224272 233758 224284
rect 273990 224272 273996 224284
rect 274048 224272 274054 224324
rect 226242 224204 226248 224256
rect 226300 224244 226306 224256
rect 239306 224244 239312 224256
rect 226300 224216 239312 224244
rect 226300 224204 226306 224216
rect 239306 224204 239312 224216
rect 239364 224244 239370 224256
rect 240042 224244 240048 224256
rect 239364 224216 240048 224244
rect 239364 224204 239370 224216
rect 240042 224204 240048 224216
rect 240100 224204 240106 224256
rect 241054 224204 241060 224256
rect 241112 224244 241118 224256
rect 241514 224244 241520 224256
rect 241112 224216 241520 224244
rect 241112 224204 241118 224216
rect 241514 224204 241520 224216
rect 241572 224244 241578 224256
rect 283650 224244 283656 224256
rect 241572 224216 283656 224244
rect 241572 224204 241578 224216
rect 283650 224204 283656 224216
rect 283708 224204 283714 224256
rect 241606 224136 241612 224188
rect 241664 224176 241670 224188
rect 251266 224176 251272 224188
rect 241664 224148 251272 224176
rect 241664 224136 241670 224148
rect 251266 224136 251272 224148
rect 251324 224176 251330 224188
rect 286318 224176 286324 224188
rect 251324 224148 286324 224176
rect 251324 224136 251330 224148
rect 286318 224136 286324 224148
rect 286376 224136 286382 224188
rect 243722 224068 243728 224120
rect 243780 224108 243786 224120
rect 243998 224108 244004 224120
rect 243780 224080 244004 224108
rect 243780 224068 243786 224080
rect 243998 224068 244004 224080
rect 244056 224108 244062 224120
rect 277118 224108 277124 224120
rect 244056 224080 277124 224108
rect 244056 224068 244062 224080
rect 277118 224068 277124 224080
rect 277176 224068 277182 224120
rect 206922 224040 206928 224052
rect 206848 224012 206928 224040
rect 206848 223848 206876 224012
rect 206922 224000 206928 224012
rect 206980 224000 206986 224052
rect 229830 224000 229836 224052
rect 229888 224040 229894 224052
rect 237926 224040 237932 224052
rect 229888 224012 237932 224040
rect 229888 224000 229894 224012
rect 237926 224000 237932 224012
rect 237984 224040 237990 224052
rect 300854 224040 300860 224052
rect 237984 224012 300860 224040
rect 237984 224000 237990 224012
rect 300854 224000 300860 224012
rect 300912 224000 300918 224052
rect 265526 223932 265532 223984
rect 265584 223972 265590 223984
rect 265802 223972 265808 223984
rect 265584 223944 265808 223972
rect 265584 223932 265590 223944
rect 265802 223932 265808 223944
rect 265860 223932 265866 223984
rect 206830 223796 206836 223848
rect 206888 223796 206894 223848
rect 227346 223592 227352 223644
rect 227404 223632 227410 223644
rect 233694 223632 233700 223644
rect 227404 223604 233700 223632
rect 227404 223592 227410 223604
rect 233694 223592 233700 223604
rect 233752 223592 233758 223644
rect 258626 223592 258632 223644
rect 258684 223632 258690 223644
rect 264146 223632 264152 223644
rect 258684 223604 264152 223632
rect 258684 223592 258690 223604
rect 264146 223592 264152 223604
rect 264204 223592 264210 223644
rect 258810 223524 258816 223576
rect 258868 223564 258874 223576
rect 259178 223564 259184 223576
rect 258868 223536 259184 223564
rect 258868 223524 258874 223536
rect 259178 223524 259184 223536
rect 259236 223564 259242 223576
rect 319806 223564 319812 223576
rect 259236 223536 319812 223564
rect 259236 223524 259242 223536
rect 319806 223524 319812 223536
rect 319864 223524 319870 223576
rect 259362 223456 259368 223508
rect 259420 223496 259426 223508
rect 262950 223496 262956 223508
rect 259420 223468 262956 223496
rect 259420 223456 259426 223468
rect 262950 223456 262956 223468
rect 263008 223456 263014 223508
rect 264146 223456 264152 223508
rect 264204 223496 264210 223508
rect 319714 223496 319720 223508
rect 264204 223468 319720 223496
rect 264204 223456 264210 223468
rect 319714 223456 319720 223468
rect 319772 223456 319778 223508
rect 256878 223388 256884 223440
rect 256936 223428 256942 223440
rect 257338 223428 257344 223440
rect 256936 223400 257344 223428
rect 256936 223388 256942 223400
rect 257338 223388 257344 223400
rect 257396 223428 257402 223440
rect 318242 223428 318248 223440
rect 257396 223400 318248 223428
rect 257396 223388 257402 223400
rect 318242 223388 318248 223400
rect 318300 223388 318306 223440
rect 256786 223320 256792 223372
rect 256844 223360 256850 223372
rect 257430 223360 257436 223372
rect 256844 223332 257436 223360
rect 256844 223320 256850 223332
rect 257430 223320 257436 223332
rect 257488 223360 257494 223372
rect 318150 223360 318156 223372
rect 257488 223332 318156 223360
rect 257488 223320 257494 223332
rect 318150 223320 318156 223332
rect 318208 223320 318214 223372
rect 257706 223252 257712 223304
rect 257764 223292 257770 223304
rect 257764 223264 262904 223292
rect 257764 223252 257770 223264
rect 254210 223184 254216 223236
rect 254268 223224 254274 223236
rect 254854 223224 254860 223236
rect 254268 223196 254860 223224
rect 254268 223184 254274 223196
rect 254854 223184 254860 223196
rect 254912 223224 254918 223236
rect 262876 223224 262904 223264
rect 262950 223252 262956 223304
rect 263008 223292 263014 223304
rect 316678 223292 316684 223304
rect 263008 223264 316684 223292
rect 263008 223252 263014 223264
rect 316678 223252 316684 223264
rect 316736 223252 316742 223304
rect 316862 223224 316868 223236
rect 254912 223196 259500 223224
rect 262876 223196 316868 223224
rect 254912 223184 254918 223196
rect 255590 223116 255596 223168
rect 255648 223156 255654 223168
rect 256142 223156 256148 223168
rect 255648 223128 256148 223156
rect 255648 223116 255654 223128
rect 256142 223116 256148 223128
rect 256200 223156 256206 223168
rect 259362 223156 259368 223168
rect 256200 223128 259368 223156
rect 256200 223116 256206 223128
rect 259362 223116 259368 223128
rect 259420 223116 259426 223168
rect 259472 223156 259500 223196
rect 316862 223184 316868 223196
rect 316920 223184 316926 223236
rect 314286 223156 314292 223168
rect 259472 223128 314292 223156
rect 314286 223116 314292 223128
rect 314344 223116 314350 223168
rect 254302 223048 254308 223100
rect 254360 223088 254366 223100
rect 314194 223088 314200 223100
rect 254360 223060 314200 223088
rect 254360 223048 254366 223060
rect 314194 223048 314200 223060
rect 314252 223048 314258 223100
rect 289078 223020 289084 223032
rect 230032 222992 289084 223020
rect 230032 222964 230060 222992
rect 289078 222980 289084 222992
rect 289136 222980 289142 223032
rect 306466 223020 306472 223032
rect 296686 222992 306472 223020
rect 158622 222912 158628 222964
rect 158680 222952 158686 222964
rect 205634 222952 205640 222964
rect 158680 222924 205640 222952
rect 158680 222912 158686 222924
rect 205634 222912 205640 222924
rect 205692 222912 205698 222964
rect 229370 222912 229376 222964
rect 229428 222952 229434 222964
rect 230014 222952 230020 222964
rect 229428 222924 230020 222952
rect 229428 222912 229434 222924
rect 230014 222912 230020 222924
rect 230072 222912 230078 222964
rect 232774 222912 232780 222964
rect 232832 222952 232838 222964
rect 276658 222952 276664 222964
rect 232832 222924 276664 222952
rect 232832 222912 232838 222924
rect 276658 222912 276664 222924
rect 276716 222912 276722 222964
rect 162302 222844 162308 222896
rect 162360 222884 162366 222896
rect 237098 222884 237104 222896
rect 162360 222856 237104 222884
rect 162360 222844 162366 222856
rect 237098 222844 237104 222856
rect 237156 222844 237162 222896
rect 247494 222844 247500 222896
rect 247552 222884 247558 222896
rect 247770 222884 247776 222896
rect 247552 222856 247776 222884
rect 247552 222844 247558 222856
rect 247770 222844 247776 222856
rect 247828 222884 247834 222896
rect 296686 222884 296714 222992
rect 306466 222980 306472 222992
rect 306524 223020 306530 223032
rect 307110 223020 307116 223032
rect 306524 222992 307116 223020
rect 306524 222980 306530 222992
rect 307110 222980 307116 222992
rect 307168 222980 307174 223032
rect 247828 222856 296714 222884
rect 247828 222844 247834 222856
rect 253106 222776 253112 222828
rect 253164 222816 253170 222828
rect 271966 222816 271972 222828
rect 253164 222788 271972 222816
rect 253164 222776 253170 222788
rect 271966 222776 271972 222788
rect 272024 222816 272030 222828
rect 272518 222816 272524 222828
rect 272024 222788 272524 222816
rect 272024 222776 272030 222788
rect 272518 222776 272524 222788
rect 272576 222776 272582 222828
rect 262306 222708 262312 222760
rect 262364 222748 262370 222760
rect 262950 222748 262956 222760
rect 262364 222720 262956 222748
rect 262364 222708 262370 222720
rect 262950 222708 262956 222720
rect 263008 222708 263014 222760
rect 242986 222096 242992 222148
rect 243044 222136 243050 222148
rect 243630 222136 243636 222148
rect 243044 222108 243636 222136
rect 243044 222096 243050 222108
rect 243630 222096 243636 222108
rect 243688 222096 243694 222148
rect 248598 222096 248604 222148
rect 248656 222136 248662 222148
rect 249334 222136 249340 222148
rect 248656 222108 249340 222136
rect 248656 222096 248662 222108
rect 249334 222096 249340 222108
rect 249392 222096 249398 222148
rect 252738 222096 252744 222148
rect 252796 222136 252802 222148
rect 253198 222136 253204 222148
rect 252796 222108 253204 222136
rect 252796 222096 252802 222108
rect 253198 222096 253204 222108
rect 253256 222096 253262 222148
rect 254118 222096 254124 222148
rect 254176 222136 254182 222148
rect 254670 222136 254676 222148
rect 254176 222108 254676 222136
rect 254176 222096 254182 222108
rect 254670 222096 254676 222108
rect 254728 222096 254734 222148
rect 254946 222096 254952 222148
rect 255004 222136 255010 222148
rect 328454 222136 328460 222148
rect 255004 222108 328460 222136
rect 255004 222096 255010 222108
rect 328454 222096 328460 222108
rect 328512 222096 328518 222148
rect 252646 222028 252652 222080
rect 252704 222068 252710 222080
rect 253474 222068 253480 222080
rect 252704 222040 253480 222068
rect 252704 222028 252710 222040
rect 253474 222028 253480 222040
rect 253532 222028 253538 222080
rect 312814 222068 312820 222080
rect 254688 222040 312820 222068
rect 252186 221960 252192 222012
rect 252244 222000 252250 222012
rect 254688 222000 254716 222040
rect 312814 222028 312820 222040
rect 312872 222028 312878 222080
rect 252244 221972 254716 222000
rect 252244 221960 252250 221972
rect 254762 221960 254768 222012
rect 254820 222000 254826 222012
rect 315298 222000 315304 222012
rect 254820 221972 315304 222000
rect 254820 221960 254826 221972
rect 315298 221960 315304 221972
rect 315356 221960 315362 222012
rect 232590 221892 232596 221944
rect 232648 221932 232654 221944
rect 232648 221904 238754 221932
rect 232648 221892 232654 221904
rect 238726 221864 238754 221904
rect 253290 221892 253296 221944
rect 253348 221932 253354 221944
rect 254946 221932 254952 221944
rect 253348 221904 254952 221932
rect 253348 221892 253354 221904
rect 254946 221892 254952 221904
rect 255004 221892 255010 221944
rect 255498 221892 255504 221944
rect 255556 221932 255562 221944
rect 255958 221932 255964 221944
rect 255556 221904 255964 221932
rect 255556 221892 255562 221904
rect 255958 221892 255964 221904
rect 256016 221932 256022 221944
rect 316770 221932 316776 221944
rect 256016 221904 316776 221932
rect 256016 221892 256022 221904
rect 316770 221892 316776 221904
rect 316828 221892 316834 221944
rect 253934 221864 253940 221876
rect 238726 221836 253940 221864
rect 253934 221824 253940 221836
rect 253992 221824 253998 221876
rect 254670 221824 254676 221876
rect 254728 221864 254734 221876
rect 314378 221864 314384 221876
rect 254728 221836 314384 221864
rect 254728 221824 254734 221836
rect 314378 221824 314384 221836
rect 314436 221824 314442 221876
rect 253474 221756 253480 221808
rect 253532 221796 253538 221808
rect 312630 221796 312636 221808
rect 253532 221768 312636 221796
rect 253532 221756 253538 221768
rect 312630 221756 312636 221768
rect 312688 221756 312694 221808
rect 253198 221688 253204 221740
rect 253256 221728 253262 221740
rect 312722 221728 312728 221740
rect 253256 221700 312728 221728
rect 253256 221688 253262 221700
rect 312722 221688 312728 221700
rect 312780 221688 312786 221740
rect 243630 221620 243636 221672
rect 243688 221660 243694 221672
rect 287882 221660 287888 221672
rect 243688 221632 287888 221660
rect 243688 221620 243694 221632
rect 287882 221620 287888 221632
rect 287940 221620 287946 221672
rect 230750 221552 230756 221604
rect 230808 221592 230814 221604
rect 231486 221592 231492 221604
rect 230808 221564 231492 221592
rect 230808 221552 230814 221564
rect 231486 221552 231492 221564
rect 231544 221592 231550 221604
rect 271874 221592 271880 221604
rect 231544 221564 271880 221592
rect 231544 221552 231550 221564
rect 271874 221552 271880 221564
rect 271932 221552 271938 221604
rect 228634 221484 228640 221536
rect 228692 221524 228698 221536
rect 262214 221524 262220 221536
rect 228692 221496 262220 221524
rect 228692 221484 228698 221496
rect 262214 221484 262220 221496
rect 262272 221484 262278 221536
rect 162210 221416 162216 221468
rect 162268 221456 162274 221468
rect 236730 221456 236736 221468
rect 162268 221428 236736 221456
rect 162268 221416 162274 221428
rect 236730 221416 236736 221428
rect 236788 221416 236794 221468
rect 249334 221416 249340 221468
rect 249392 221456 249398 221468
rect 339494 221456 339500 221468
rect 249392 221428 339500 221456
rect 249392 221416 249398 221428
rect 339494 221416 339500 221428
rect 339552 221416 339558 221468
rect 254026 221348 254032 221400
rect 254084 221388 254090 221400
rect 254762 221388 254768 221400
rect 254084 221360 254768 221388
rect 254084 221348 254090 221360
rect 254762 221348 254768 221360
rect 254820 221348 254826 221400
rect 223942 220736 223948 220788
rect 224000 220776 224006 220788
rect 224310 220776 224316 220788
rect 224000 220748 224316 220776
rect 224000 220736 224006 220748
rect 224310 220736 224316 220748
rect 224368 220736 224374 220788
rect 227438 220736 227444 220788
rect 227496 220776 227502 220788
rect 288250 220776 288256 220788
rect 227496 220748 288256 220776
rect 227496 220736 227502 220748
rect 288250 220736 288256 220748
rect 288308 220736 288314 220788
rect 223850 220668 223856 220720
rect 223908 220708 223914 220720
rect 224494 220708 224500 220720
rect 223908 220680 224500 220708
rect 223908 220668 223914 220680
rect 224494 220668 224500 220680
rect 224552 220668 224558 220720
rect 284478 220708 284484 220720
rect 224926 220680 284484 220708
rect 224310 220600 224316 220652
rect 224368 220640 224374 220652
rect 224926 220640 224954 220680
rect 284478 220668 284484 220680
rect 284536 220668 284542 220720
rect 284294 220640 284300 220652
rect 224368 220612 224954 220640
rect 229756 220612 284300 220640
rect 224368 220600 224374 220612
rect 224494 220464 224500 220516
rect 224552 220504 224558 220516
rect 229756 220504 229784 220612
rect 284294 220600 284300 220612
rect 284352 220600 284358 220652
rect 286594 220572 286600 220584
rect 224552 220476 229784 220504
rect 229848 220544 286600 220572
rect 224552 220464 224558 220476
rect 226426 220396 226432 220448
rect 226484 220436 226490 220448
rect 227438 220436 227444 220448
rect 226484 220408 227444 220436
rect 226484 220396 226490 220408
rect 227438 220396 227444 220408
rect 227496 220396 227502 220448
rect 229848 220368 229876 220544
rect 286594 220532 286600 220544
rect 286652 220532 286658 220584
rect 283834 220504 283840 220516
rect 227272 220340 229876 220368
rect 229940 220476 283840 220504
rect 227272 220312 227300 220340
rect 226518 220260 226524 220312
rect 226576 220300 226582 220312
rect 227254 220300 227260 220312
rect 226576 220272 227260 220300
rect 226576 220260 226582 220272
rect 227254 220260 227260 220272
rect 227312 220260 227318 220312
rect 229278 220260 229284 220312
rect 229336 220300 229342 220312
rect 229940 220300 229968 220476
rect 283834 220464 283840 220476
rect 283892 220464 283898 220516
rect 275002 220436 275008 220448
rect 229336 220272 229968 220300
rect 234586 220408 275008 220436
rect 229336 220260 229342 220272
rect 225874 220192 225880 220244
rect 225932 220232 225938 220244
rect 234586 220232 234614 220408
rect 275002 220396 275008 220408
rect 275060 220396 275066 220448
rect 248506 220328 248512 220380
rect 248564 220368 248570 220380
rect 249150 220368 249156 220380
rect 248564 220340 249156 220368
rect 248564 220328 248570 220340
rect 249150 220328 249156 220340
rect 249208 220328 249214 220380
rect 225932 220204 234614 220232
rect 225932 220192 225938 220204
rect 158070 220056 158076 220108
rect 158128 220096 158134 220108
rect 229278 220096 229284 220108
rect 158128 220068 229284 220096
rect 158128 220056 158134 220068
rect 229278 220056 229284 220068
rect 229336 220056 229342 220108
rect 249150 220056 249156 220108
rect 249208 220096 249214 220108
rect 309778 220096 309784 220108
rect 249208 220068 309784 220096
rect 249208 220056 249214 220068
rect 309778 220056 309784 220068
rect 309836 220056 309842 220108
rect 229186 219376 229192 219428
rect 229244 219416 229250 219428
rect 229922 219416 229928 219428
rect 229244 219388 229928 219416
rect 229244 219376 229250 219388
rect 229922 219376 229928 219388
rect 229980 219376 229986 219428
rect 289446 219416 289452 219428
rect 230032 219388 289452 219416
rect 228910 219308 228916 219360
rect 228968 219348 228974 219360
rect 230032 219348 230060 219388
rect 289446 219376 289452 219388
rect 289504 219376 289510 219428
rect 228968 219320 230060 219348
rect 228968 219308 228974 219320
rect 230566 219308 230572 219360
rect 230624 219348 230630 219360
rect 231762 219348 231768 219360
rect 230624 219320 231768 219348
rect 230624 219308 230630 219320
rect 231762 219308 231768 219320
rect 231820 219348 231826 219360
rect 290458 219348 290464 219360
rect 231820 219320 290464 219348
rect 231820 219308 231826 219320
rect 290458 219308 290464 219320
rect 290516 219308 290522 219360
rect 246390 219240 246396 219292
rect 246448 219280 246454 219292
rect 249978 219280 249984 219292
rect 246448 219252 249984 219280
rect 246448 219240 246454 219252
rect 249978 219240 249984 219252
rect 250036 219280 250042 219292
rect 309870 219280 309876 219292
rect 250036 219252 309876 219280
rect 250036 219240 250042 219252
rect 309870 219240 309876 219252
rect 309928 219240 309934 219292
rect 256510 219172 256516 219224
rect 256568 219212 256574 219224
rect 314010 219212 314016 219224
rect 256568 219184 314016 219212
rect 256568 219172 256574 219184
rect 314010 219172 314016 219184
rect 314068 219172 314074 219224
rect 246758 219104 246764 219156
rect 246816 219144 246822 219156
rect 289538 219144 289544 219156
rect 246816 219116 289544 219144
rect 246816 219104 246822 219116
rect 289538 219104 289544 219116
rect 289596 219104 289602 219156
rect 229922 219036 229928 219088
rect 229980 219076 229986 219088
rect 273346 219076 273352 219088
rect 229980 219048 273352 219076
rect 229980 219036 229986 219048
rect 273346 219036 273352 219048
rect 273404 219036 273410 219088
rect 243906 218968 243912 219020
rect 243964 219008 243970 219020
rect 282178 219008 282184 219020
rect 243964 218980 282184 219008
rect 243964 218968 243970 218980
rect 282178 218968 282184 218980
rect 282236 218968 282242 219020
rect 152642 218764 152648 218816
rect 152700 218804 152706 218816
rect 228266 218804 228272 218816
rect 152700 218776 228272 218804
rect 152700 218764 152706 218776
rect 228266 218764 228272 218776
rect 228324 218804 228330 218816
rect 228910 218804 228916 218816
rect 228324 218776 228916 218804
rect 228324 218764 228330 218776
rect 228910 218764 228916 218776
rect 228968 218764 228974 218816
rect 160738 218696 160744 218748
rect 160796 218736 160802 218748
rect 237558 218736 237564 218748
rect 160796 218708 237564 218736
rect 160796 218696 160802 218708
rect 237558 218696 237564 218708
rect 237616 218696 237622 218748
rect 249518 218696 249524 218748
rect 249576 218736 249582 218748
rect 335354 218736 335360 218748
rect 249576 218708 335360 218736
rect 249576 218696 249582 218708
rect 335354 218696 335360 218708
rect 335412 218736 335418 218748
rect 335998 218736 336004 218748
rect 335412 218708 336004 218736
rect 335412 218696 335418 218708
rect 335998 218696 336004 218708
rect 336056 218696 336062 218748
rect 249242 218016 249248 218068
rect 249300 218056 249306 218068
rect 249518 218056 249524 218068
rect 249300 218028 249524 218056
rect 249300 218016 249306 218028
rect 249518 218016 249524 218028
rect 249576 218016 249582 218068
rect 204162 217948 204168 218000
rect 204220 217988 204226 218000
rect 225506 217988 225512 218000
rect 204220 217960 225512 217988
rect 204220 217948 204226 217960
rect 225506 217948 225512 217960
rect 225564 217948 225570 218000
rect 180150 217404 180156 217456
rect 180208 217444 180214 217456
rect 212902 217444 212908 217456
rect 180208 217416 212908 217444
rect 180208 217404 180214 217416
rect 212902 217404 212908 217416
rect 212960 217404 212966 217456
rect 303614 217404 303620 217456
rect 303672 217444 303678 217456
rect 304258 217444 304264 217456
rect 303672 217416 304264 217444
rect 303672 217404 303678 217416
rect 304258 217404 304264 217416
rect 304316 217404 304322 217456
rect 165338 217336 165344 217388
rect 165396 217376 165402 217388
rect 204162 217376 204168 217388
rect 165396 217348 204168 217376
rect 165396 217336 165402 217348
rect 204162 217336 204168 217348
rect 204220 217336 204226 217388
rect 166810 217268 166816 217320
rect 166868 217308 166874 217320
rect 226702 217308 226708 217320
rect 166868 217280 226708 217308
rect 166868 217268 166874 217280
rect 226702 217268 226708 217280
rect 226760 217268 226766 217320
rect 246574 217268 246580 217320
rect 246632 217308 246638 217320
rect 303614 217308 303620 217320
rect 246632 217280 303620 217308
rect 246632 217268 246638 217280
rect 303614 217268 303620 217280
rect 303672 217268 303678 217320
rect 205634 216588 205640 216640
rect 205692 216628 205698 216640
rect 206922 216628 206928 216640
rect 205692 216600 206928 216628
rect 205692 216588 205698 216600
rect 206922 216588 206928 216600
rect 206980 216628 206986 216640
rect 224678 216628 224684 216640
rect 206980 216600 224684 216628
rect 206980 216588 206986 216600
rect 224678 216588 224684 216600
rect 224736 216588 224742 216640
rect 188614 216044 188620 216096
rect 188672 216084 188678 216096
rect 212994 216084 213000 216096
rect 188672 216056 213000 216084
rect 188672 216044 188678 216056
rect 212994 216044 213000 216056
rect 213052 216044 213058 216096
rect 155402 215976 155408 216028
rect 155460 216016 155466 216028
rect 205634 216016 205640 216028
rect 155460 215988 205640 216016
rect 155460 215976 155466 215988
rect 205634 215976 205640 215988
rect 205692 215976 205698 216028
rect 161750 215908 161756 215960
rect 161808 215948 161814 215960
rect 223482 215948 223488 215960
rect 161808 215920 223488 215948
rect 161808 215908 161814 215920
rect 223482 215908 223488 215920
rect 223540 215908 223546 215960
rect 247126 215908 247132 215960
rect 247184 215948 247190 215960
rect 247862 215948 247868 215960
rect 247184 215920 247868 215948
rect 247184 215908 247190 215920
rect 247862 215908 247868 215920
rect 247920 215948 247926 215960
rect 317414 215948 317420 215960
rect 247920 215920 317420 215948
rect 247920 215908 247926 215920
rect 317414 215908 317420 215920
rect 317472 215908 317478 215960
rect 205634 215228 205640 215280
rect 205692 215268 205698 215280
rect 206830 215268 206836 215280
rect 205692 215240 206836 215268
rect 205692 215228 205698 215240
rect 206830 215228 206836 215240
rect 206888 215268 206894 215280
rect 227530 215268 227536 215280
rect 206888 215240 227536 215268
rect 206888 215228 206894 215240
rect 227530 215228 227536 215240
rect 227588 215228 227594 215280
rect 173894 214684 173900 214736
rect 173952 214724 173958 214736
rect 174722 214724 174728 214736
rect 173952 214696 174728 214724
rect 173952 214684 173958 214696
rect 174722 214684 174728 214696
rect 174780 214684 174786 214736
rect 176102 214684 176108 214736
rect 176160 214724 176166 214736
rect 210510 214724 210516 214736
rect 176160 214696 210516 214724
rect 176160 214684 176166 214696
rect 210510 214684 210516 214696
rect 210568 214684 210574 214736
rect 159358 214616 159364 214668
rect 159416 214656 159422 214668
rect 205634 214656 205640 214668
rect 159416 214628 205640 214656
rect 159416 214616 159422 214628
rect 205634 214616 205640 214628
rect 205692 214616 205698 214668
rect 3418 214548 3424 214600
rect 3476 214588 3482 214600
rect 200758 214588 200764 214600
rect 3476 214560 200764 214588
rect 3476 214548 3482 214560
rect 200758 214548 200764 214560
rect 200816 214548 200822 214600
rect 252554 214548 252560 214600
rect 252612 214588 252618 214600
rect 253566 214588 253572 214600
rect 252612 214560 253572 214588
rect 252612 214548 252618 214560
rect 253566 214548 253572 214560
rect 253624 214588 253630 214600
rect 313918 214588 313924 214600
rect 253624 214560 313924 214588
rect 253624 214548 253630 214560
rect 313918 214548 313924 214560
rect 313976 214548 313982 214600
rect 166994 214480 167000 214532
rect 167052 214520 167058 214532
rect 167730 214520 167736 214532
rect 167052 214492 167736 214520
rect 167052 214480 167058 214492
rect 167730 214480 167736 214492
rect 167788 214480 167794 214532
rect 168374 214480 168380 214532
rect 168432 214520 168438 214532
rect 168834 214520 168840 214532
rect 168432 214492 168840 214520
rect 168432 214480 168438 214492
rect 168834 214480 168840 214492
rect 168892 214480 168898 214532
rect 169754 214480 169760 214532
rect 169812 214520 169818 214532
rect 170306 214520 170312 214532
rect 169812 214492 170312 214520
rect 169812 214480 169818 214492
rect 170306 214480 170312 214492
rect 170364 214480 170370 214532
rect 171134 214480 171140 214532
rect 171192 214520 171198 214532
rect 172146 214520 172152 214532
rect 171192 214492 172152 214520
rect 171192 214480 171198 214492
rect 172146 214480 172152 214492
rect 172204 214480 172210 214532
rect 172514 214480 172520 214532
rect 172572 214520 172578 214532
rect 173250 214520 173256 214532
rect 172572 214492 173256 214520
rect 172572 214480 172578 214492
rect 173250 214480 173256 214492
rect 173308 214480 173314 214532
rect 173986 214480 173992 214532
rect 174044 214520 174050 214532
rect 174354 214520 174360 214532
rect 174044 214492 174360 214520
rect 174044 214480 174050 214492
rect 174354 214480 174360 214492
rect 174412 214480 174418 214532
rect 186406 214480 186412 214532
rect 186464 214520 186470 214532
rect 186866 214520 186872 214532
rect 186464 214492 186872 214520
rect 186464 214480 186470 214492
rect 186866 214480 186872 214492
rect 186924 214480 186930 214532
rect 187786 214480 187792 214532
rect 187844 214520 187850 214532
rect 188982 214520 188988 214532
rect 187844 214492 188988 214520
rect 187844 214480 187850 214492
rect 188982 214480 188988 214492
rect 189040 214480 189046 214532
rect 189074 214480 189080 214532
rect 189132 214520 189138 214532
rect 189810 214520 189816 214532
rect 189132 214492 189816 214520
rect 189132 214480 189138 214492
rect 189810 214480 189816 214492
rect 189868 214480 189874 214532
rect 190454 214480 190460 214532
rect 190512 214520 190518 214532
rect 190914 214520 190920 214532
rect 190512 214492 190920 214520
rect 190512 214480 190518 214492
rect 190914 214480 190920 214492
rect 190972 214480 190978 214532
rect 191926 214480 191932 214532
rect 191984 214520 191990 214532
rect 193030 214520 193036 214532
rect 191984 214492 193036 214520
rect 191984 214480 191990 214492
rect 193030 214480 193036 214492
rect 193088 214480 193094 214532
rect 193306 214480 193312 214532
rect 193364 214520 193370 214532
rect 193490 214520 193496 214532
rect 193364 214492 193496 214520
rect 193364 214480 193370 214492
rect 193490 214480 193496 214492
rect 193548 214480 193554 214532
rect 194594 214480 194600 214532
rect 194652 214520 194658 214532
rect 195330 214520 195336 214532
rect 194652 214492 195336 214520
rect 194652 214480 194658 214492
rect 195330 214480 195336 214492
rect 195388 214480 195394 214532
rect 186314 214412 186320 214464
rect 186372 214452 186378 214464
rect 187234 214452 187240 214464
rect 186372 214424 187240 214452
rect 186372 214412 186378 214424
rect 187234 214412 187240 214424
rect 187292 214412 187298 214464
rect 189166 214412 189172 214464
rect 189224 214452 189230 214464
rect 189442 214452 189448 214464
rect 189224 214424 189448 214452
rect 189224 214412 189230 214424
rect 189442 214412 189448 214424
rect 189500 214412 189506 214464
rect 190546 214412 190552 214464
rect 190604 214452 190610 214464
rect 190730 214452 190736 214464
rect 190604 214424 190736 214452
rect 190604 214412 190610 214424
rect 190730 214412 190736 214424
rect 190788 214412 190794 214464
rect 193214 214412 193220 214464
rect 193272 214452 193278 214464
rect 194502 214452 194508 214464
rect 193272 214424 194508 214452
rect 193272 214412 193278 214424
rect 194502 214412 194508 214424
rect 194560 214412 194566 214464
rect 194686 214412 194692 214464
rect 194744 214452 194750 214464
rect 194962 214452 194968 214464
rect 194744 214424 194968 214452
rect 194744 214412 194750 214424
rect 194962 214412 194968 214424
rect 195020 214412 195026 214464
rect 186406 214344 186412 214396
rect 186464 214384 186470 214396
rect 186682 214384 186688 214396
rect 186464 214356 186688 214384
rect 186464 214344 186470 214356
rect 186682 214344 186688 214356
rect 186740 214344 186746 214396
rect 201402 213868 201408 213920
rect 201460 213908 201466 213920
rect 223574 213908 223580 213920
rect 201460 213880 223580 213908
rect 201460 213868 201466 213880
rect 223574 213868 223580 213880
rect 223632 213868 223638 213920
rect 182358 213392 182364 213444
rect 182416 213432 182422 213444
rect 210694 213432 210700 213444
rect 182416 213404 210700 213432
rect 182416 213392 182422 213404
rect 210694 213392 210700 213404
rect 210752 213392 210758 213444
rect 181990 213324 181996 213376
rect 182048 213364 182054 213376
rect 216490 213364 216496 213376
rect 182048 213336 216496 213364
rect 182048 213324 182054 213336
rect 216490 213324 216496 213336
rect 216548 213324 216554 213376
rect 157978 213256 157984 213308
rect 158036 213296 158042 213308
rect 201402 213296 201408 213308
rect 158036 213268 201408 213296
rect 158036 213256 158042 213268
rect 201402 213256 201408 213268
rect 201460 213256 201466 213308
rect 242526 213256 242532 213308
rect 242584 213296 242590 213308
rect 252554 213296 252560 213308
rect 242584 213268 252560 213296
rect 242584 213256 242590 213268
rect 252554 213256 252560 213268
rect 252612 213256 252618 213308
rect 184750 213188 184756 213240
rect 184808 213228 184814 213240
rect 244366 213228 244372 213240
rect 184808 213200 244372 213228
rect 184808 213188 184814 213200
rect 244366 213188 244372 213200
rect 244424 213188 244430 213240
rect 250622 213188 250628 213240
rect 250680 213228 250686 213240
rect 311158 213228 311164 213240
rect 250680 213200 311164 213228
rect 250680 213188 250686 213200
rect 311158 213188 311164 213200
rect 311216 213188 311222 213240
rect 175734 212440 175740 212492
rect 175792 212480 175798 212492
rect 180058 212480 180064 212492
rect 175792 212452 180064 212480
rect 175792 212440 175798 212452
rect 180058 212440 180064 212452
rect 180116 212440 180122 212492
rect 199378 212440 199384 212492
rect 199436 212480 199442 212492
rect 220354 212480 220360 212492
rect 199436 212452 220360 212480
rect 199436 212440 199442 212452
rect 220354 212440 220360 212452
rect 220412 212440 220418 212492
rect 173894 212372 173900 212424
rect 173952 212412 173958 212424
rect 178678 212412 178684 212424
rect 173952 212384 178684 212412
rect 173952 212372 173958 212384
rect 178678 212372 178684 212384
rect 178736 212372 178742 212424
rect 181254 212372 181260 212424
rect 181312 212412 181318 212424
rect 184198 212412 184204 212424
rect 181312 212384 184204 212412
rect 181312 212372 181318 212384
rect 184198 212372 184204 212384
rect 184256 212372 184262 212424
rect 184382 212372 184388 212424
rect 184440 212412 184446 212424
rect 205542 212412 205548 212424
rect 184440 212384 186314 212412
rect 184440 212372 184446 212384
rect 176654 212304 176660 212356
rect 176712 212344 176718 212356
rect 176930 212344 176936 212356
rect 176712 212316 176936 212344
rect 176712 212304 176718 212316
rect 176930 212304 176936 212316
rect 176988 212304 176994 212356
rect 183554 212304 183560 212356
rect 183612 212344 183618 212356
rect 184290 212344 184296 212356
rect 183612 212316 184296 212344
rect 183612 212304 183618 212316
rect 184290 212304 184296 212316
rect 184348 212304 184354 212356
rect 184934 212304 184940 212356
rect 184992 212344 184998 212356
rect 185394 212344 185400 212356
rect 184992 212316 185400 212344
rect 184992 212304 184998 212316
rect 185394 212304 185400 212316
rect 185452 212304 185458 212356
rect 186286 212344 186314 212384
rect 195946 212384 205548 212412
rect 195946 212344 195974 212384
rect 205542 212372 205548 212384
rect 205600 212372 205606 212424
rect 186286 212316 195974 212344
rect 197078 212304 197084 212356
rect 197136 212344 197142 212356
rect 197136 212316 205634 212344
rect 197136 212304 197142 212316
rect 164234 212236 164240 212288
rect 164292 212276 164298 212288
rect 164786 212276 164792 212288
rect 164292 212248 164792 212276
rect 164292 212236 164298 212248
rect 164786 212236 164792 212248
rect 164844 212236 164850 212288
rect 165706 212236 165712 212288
rect 165764 212276 165770 212288
rect 166902 212276 166908 212288
rect 165764 212248 166908 212276
rect 165764 212236 165770 212248
rect 166902 212236 166908 212248
rect 166960 212236 166966 212288
rect 176838 212236 176844 212288
rect 176896 212276 176902 212288
rect 177666 212276 177672 212288
rect 176896 212248 177672 212276
rect 176896 212236 176902 212248
rect 177666 212236 177672 212248
rect 177724 212236 177730 212288
rect 178034 212236 178040 212288
rect 178092 212276 178098 212288
rect 178770 212276 178776 212288
rect 178092 212248 178776 212276
rect 178092 212236 178098 212248
rect 178770 212236 178776 212248
rect 178828 212236 178834 212288
rect 183646 212236 183652 212288
rect 183704 212276 183710 212288
rect 183922 212276 183928 212288
rect 183704 212248 183928 212276
rect 183704 212236 183710 212248
rect 183922 212236 183928 212248
rect 183980 212236 183986 212288
rect 185118 212236 185124 212288
rect 185176 212276 185182 212288
rect 185762 212276 185768 212288
rect 185176 212248 185768 212276
rect 185176 212236 185182 212248
rect 185762 212236 185768 212248
rect 185820 212236 185826 212288
rect 185854 212236 185860 212288
rect 185912 212276 185918 212288
rect 188338 212276 188344 212288
rect 185912 212248 188344 212276
rect 185912 212236 185918 212248
rect 188338 212236 188344 212248
rect 188396 212236 188402 212288
rect 195974 212236 195980 212288
rect 196032 212276 196038 212288
rect 196434 212276 196440 212288
rect 196032 212248 196440 212276
rect 196032 212236 196038 212248
rect 196434 212236 196440 212248
rect 196492 212236 196498 212288
rect 197354 212236 197360 212288
rect 197412 212276 197418 212288
rect 198550 212276 198556 212288
rect 197412 212248 198556 212276
rect 197412 212236 197418 212248
rect 198550 212236 198556 212248
rect 198608 212236 198614 212288
rect 198918 212236 198924 212288
rect 198976 212276 198982 212288
rect 200022 212276 200028 212288
rect 198976 212248 200028 212276
rect 198976 212236 198982 212248
rect 200022 212236 200028 212248
rect 200080 212236 200086 212288
rect 205606 212276 205634 212316
rect 221642 212276 221648 212288
rect 205606 212248 221648 212276
rect 221642 212236 221648 212248
rect 221700 212236 221706 212288
rect 173526 212168 173532 212220
rect 173584 212208 173590 212220
rect 173802 212208 173808 212220
rect 173584 212180 173808 212208
rect 173584 212168 173590 212180
rect 173802 212168 173808 212180
rect 173860 212208 173866 212220
rect 188798 212208 188804 212220
rect 173860 212180 188804 212208
rect 173860 212168 173866 212180
rect 188798 212168 188804 212180
rect 188856 212168 188862 212220
rect 194134 212168 194140 212220
rect 194192 212208 194198 212220
rect 221550 212208 221556 212220
rect 194192 212180 221556 212208
rect 194192 212168 194198 212180
rect 221550 212168 221556 212180
rect 221608 212168 221614 212220
rect 175366 212100 175372 212152
rect 175424 212140 175430 212152
rect 216582 212140 216588 212152
rect 175424 212112 216588 212140
rect 175424 212100 175430 212112
rect 216582 212100 216588 212112
rect 216640 212100 216646 212152
rect 159266 212032 159272 212084
rect 159324 212072 159330 212084
rect 201218 212072 201224 212084
rect 159324 212044 201224 212072
rect 159324 212032 159330 212044
rect 201218 212032 201224 212044
rect 201276 212032 201282 212084
rect 202690 212032 202696 212084
rect 202748 212072 202754 212084
rect 203334 212072 203340 212084
rect 202748 212044 203340 212072
rect 202748 212032 202754 212044
rect 203334 212032 203340 212044
rect 203392 212032 203398 212084
rect 204070 212032 204076 212084
rect 204128 212072 204134 212084
rect 204806 212072 204812 212084
rect 204128 212044 204812 212072
rect 204128 212032 204134 212044
rect 204806 212032 204812 212044
rect 204864 212032 204870 212084
rect 180518 211964 180524 212016
rect 180576 212004 180582 212016
rect 221734 212004 221740 212016
rect 180576 211976 221740 212004
rect 180576 211964 180582 211976
rect 221734 211964 221740 211976
rect 221792 211964 221798 212016
rect 165706 211896 165712 211948
rect 165764 211936 165770 211948
rect 165890 211936 165896 211948
rect 165764 211908 165896 211936
rect 165764 211896 165770 211908
rect 165890 211896 165896 211908
rect 165948 211896 165954 211948
rect 172054 211896 172060 211948
rect 172112 211936 172118 211948
rect 213730 211936 213736 211948
rect 172112 211908 213736 211936
rect 172112 211896 172118 211908
rect 213730 211896 213736 211908
rect 213788 211896 213794 211948
rect 155218 211828 155224 211880
rect 155276 211868 155282 211880
rect 204070 211868 204076 211880
rect 155276 211840 204076 211868
rect 155276 211828 155282 211840
rect 204070 211828 204076 211840
rect 204128 211828 204134 211880
rect 28258 211760 28264 211812
rect 28316 211800 28322 211812
rect 202690 211800 202696 211812
rect 28316 211772 202696 211800
rect 28316 211760 28322 211772
rect 202690 211760 202696 211772
rect 202748 211760 202754 211812
rect 203702 211760 203708 211812
rect 203760 211800 203766 211812
rect 272058 211800 272064 211812
rect 203760 211772 272064 211800
rect 203760 211760 203766 211772
rect 272058 211760 272064 211772
rect 272116 211760 272122 211812
rect 167638 211692 167644 211744
rect 167696 211732 167702 211744
rect 168282 211732 168288 211744
rect 167696 211704 168288 211732
rect 167696 211692 167702 211704
rect 168282 211692 168288 211704
rect 168340 211692 168346 211744
rect 178586 211692 178592 211744
rect 178644 211732 178650 211744
rect 185854 211732 185860 211744
rect 178644 211704 185860 211732
rect 178644 211692 178650 211704
rect 185854 211692 185860 211704
rect 185912 211692 185918 211744
rect 195974 211692 195980 211744
rect 196032 211732 196038 211744
rect 196158 211732 196164 211744
rect 196032 211704 196164 211732
rect 196032 211692 196038 211704
rect 196158 211692 196164 211704
rect 196216 211692 196222 211744
rect 168742 211352 168748 211404
rect 168800 211392 168806 211404
rect 169662 211392 169668 211404
rect 168800 211364 169668 211392
rect 168800 211352 168806 211364
rect 169662 211352 169668 211364
rect 169720 211392 169726 211404
rect 187326 211392 187332 211404
rect 169720 211364 187332 211392
rect 169720 211352 169726 211364
rect 187326 211352 187332 211364
rect 187384 211352 187390 211404
rect 187786 211352 187792 211404
rect 187844 211392 187850 211404
rect 202138 211392 202144 211404
rect 187844 211364 202144 211392
rect 187844 211352 187850 211364
rect 202138 211352 202144 211364
rect 202196 211352 202202 211404
rect 169754 211284 169760 211336
rect 169812 211324 169818 211336
rect 173526 211324 173532 211336
rect 169812 211296 173532 211324
rect 169812 211284 169818 211296
rect 173526 211284 173532 211296
rect 173584 211284 173590 211336
rect 178678 211284 178684 211336
rect 178736 211324 178742 211336
rect 203702 211324 203708 211336
rect 178736 211296 203708 211324
rect 178736 211284 178742 211296
rect 203702 211284 203708 211296
rect 203760 211284 203766 211336
rect 162578 211216 162584 211268
rect 162636 211256 162642 211268
rect 166534 211256 166540 211268
rect 162636 211228 166540 211256
rect 162636 211216 162642 211228
rect 166534 211216 166540 211228
rect 166592 211216 166598 211268
rect 168282 211216 168288 211268
rect 168340 211256 168346 211268
rect 196250 211256 196256 211268
rect 168340 211228 196256 211256
rect 168340 211216 168346 211228
rect 196250 211216 196256 211228
rect 196308 211216 196314 211268
rect 157886 211148 157892 211200
rect 157944 211188 157950 211200
rect 202322 211188 202328 211200
rect 157944 211160 202328 211188
rect 157944 211148 157950 211160
rect 202322 211148 202328 211160
rect 202380 211148 202386 211200
rect 197354 211080 197360 211132
rect 197412 211120 197418 211132
rect 197538 211120 197544 211132
rect 197412 211092 197544 211120
rect 197412 211080 197418 211092
rect 197538 211080 197544 211092
rect 197596 211080 197602 211132
rect 179598 210876 179604 210928
rect 179656 210916 179662 210928
rect 179782 210916 179788 210928
rect 179656 210888 179788 210916
rect 179656 210876 179662 210888
rect 179782 210876 179788 210888
rect 179840 210876 179846 210928
rect 200206 210808 200212 210860
rect 200264 210848 200270 210860
rect 201126 210848 201132 210860
rect 200264 210820 201132 210848
rect 200264 210808 200270 210820
rect 201126 210808 201132 210820
rect 201184 210808 201190 210860
rect 184934 210740 184940 210792
rect 184992 210780 184998 210792
rect 185210 210780 185216 210792
rect 184992 210752 185216 210780
rect 184992 210740 184998 210752
rect 185210 210740 185216 210752
rect 185268 210740 185274 210792
rect 3510 210536 3516 210588
rect 3568 210576 3574 210588
rect 178678 210576 178684 210588
rect 3568 210548 178684 210576
rect 3568 210536 3574 210548
rect 178678 210536 178684 210548
rect 178736 210536 178742 210588
rect 183094 210536 183100 210588
rect 183152 210576 183158 210588
rect 213178 210576 213184 210588
rect 183152 210548 213184 210576
rect 183152 210536 183158 210548
rect 213178 210536 213184 210548
rect 213236 210536 213242 210588
rect 3418 210468 3424 210520
rect 3476 210508 3482 210520
rect 184382 210508 184388 210520
rect 3476 210480 184388 210508
rect 3476 210468 3482 210480
rect 184382 210468 184388 210480
rect 184440 210468 184446 210520
rect 3602 210400 3608 210452
rect 3660 210440 3666 210452
rect 187786 210440 187792 210452
rect 3660 210412 187792 210440
rect 3660 210400 3666 210412
rect 187786 210400 187792 210412
rect 187844 210400 187850 210452
rect 205266 210400 205272 210452
rect 205324 210440 205330 210452
rect 218790 210440 218796 210452
rect 205324 210412 218796 210440
rect 205324 210400 205330 210412
rect 218790 210400 218796 210412
rect 218848 210400 218854 210452
rect 198366 209992 198372 210044
rect 198424 210032 198430 210044
rect 204346 210032 204352 210044
rect 198424 210004 204352 210032
rect 198424 209992 198430 210004
rect 204346 209992 204352 210004
rect 204404 210032 204410 210044
rect 205358 210032 205364 210044
rect 204404 210004 205364 210032
rect 204404 209992 204410 210004
rect 205358 209992 205364 210004
rect 205416 209992 205422 210044
rect 160554 209924 160560 209976
rect 160612 209964 160618 209976
rect 200206 209964 200212 209976
rect 160612 209936 200212 209964
rect 160612 209924 160618 209936
rect 200206 209924 200212 209936
rect 200264 209924 200270 209976
rect 156598 209856 156604 209908
rect 156656 209896 156662 209908
rect 156656 209868 199516 209896
rect 156656 209856 156662 209868
rect 153838 209788 153844 209840
rect 153896 209828 153902 209840
rect 198366 209828 198372 209840
rect 153896 209800 198372 209828
rect 153896 209788 153902 209800
rect 198366 209788 198372 209800
rect 198424 209788 198430 209840
rect 199488 209828 199516 209868
rect 199562 209856 199568 209908
rect 199620 209896 199626 209908
rect 199930 209896 199936 209908
rect 199620 209868 199936 209896
rect 199620 209856 199626 209868
rect 199930 209856 199936 209868
rect 199988 209856 199994 209908
rect 204254 209828 204260 209840
rect 199488 209800 204260 209828
rect 204254 209788 204260 209800
rect 204312 209788 204318 209840
rect 203150 209556 203156 209568
rect 202064 209528 203156 209556
rect 159450 209380 159456 209432
rect 159508 209420 159514 209432
rect 163590 209420 163596 209432
rect 159508 209392 163596 209420
rect 159508 209380 159514 209392
rect 163590 209380 163596 209392
rect 163648 209380 163654 209432
rect 201678 209420 201684 209432
rect 176626 209392 201684 209420
rect 160646 209176 160652 209228
rect 160704 209216 160710 209228
rect 176626 209216 176654 209392
rect 201678 209380 201684 209392
rect 201736 209380 201742 209432
rect 160704 209188 176654 209216
rect 160704 209176 160710 209188
rect 146938 209108 146944 209160
rect 146996 209148 147002 209160
rect 202064 209148 202092 209528
rect 203150 209516 203156 209528
rect 203208 209556 203214 209568
rect 203886 209556 203892 209568
rect 203208 209528 203892 209556
rect 203208 209516 203214 209528
rect 203886 209516 203892 209528
rect 203944 209516 203950 209568
rect 202874 209488 202880 209500
rect 146996 209120 202092 209148
rect 202156 209460 202880 209488
rect 146996 209108 147002 209120
rect 120810 209040 120816 209092
rect 120868 209080 120874 209092
rect 202156 209080 202184 209460
rect 202874 209448 202880 209460
rect 202932 209448 202938 209500
rect 204990 209420 204996 209432
rect 120868 209052 202184 209080
rect 202248 209392 204996 209420
rect 120868 209040 120874 209052
rect 202248 209012 202276 209392
rect 204990 209380 204996 209392
rect 205048 209380 205054 209432
rect 195946 208984 202276 209012
rect 11698 208360 11704 208412
rect 11756 208400 11762 208412
rect 195946 208400 195974 208984
rect 11756 208372 195974 208400
rect 11756 208360 11762 208372
rect 209314 207680 209320 207732
rect 209372 207720 209378 207732
rect 264514 207720 264520 207732
rect 209372 207692 264520 207720
rect 209372 207680 209378 207692
rect 264514 207680 264520 207692
rect 264572 207680 264578 207732
rect 209406 207612 209412 207664
rect 209464 207652 209470 207664
rect 265802 207652 265808 207664
rect 209464 207624 265808 207652
rect 209464 207612 209470 207624
rect 265802 207612 265808 207624
rect 265860 207612 265866 207664
rect 209590 206320 209596 206372
rect 209648 206360 209654 206372
rect 260282 206360 260288 206372
rect 209648 206332 260288 206360
rect 209648 206320 209654 206332
rect 260282 206320 260288 206332
rect 260340 206320 260346 206372
rect 209498 206252 209504 206304
rect 209556 206292 209562 206304
rect 264422 206292 264428 206304
rect 209556 206264 264428 206292
rect 209556 206252 209562 206264
rect 264422 206252 264428 206264
rect 264480 206252 264486 206304
rect 209682 204960 209688 205012
rect 209740 205000 209746 205012
rect 261662 205000 261668 205012
rect 209740 204972 261668 205000
rect 209740 204960 209746 204972
rect 261662 204960 261668 204972
rect 261720 204960 261726 205012
rect 249794 204892 249800 204944
rect 249852 204932 249858 204944
rect 250438 204932 250444 204944
rect 249852 204904 250444 204932
rect 249852 204892 249858 204904
rect 250438 204892 250444 204904
rect 250496 204932 250502 204944
rect 250496 204904 316034 204932
rect 250496 204892 250502 204904
rect 316006 204864 316034 204904
rect 327258 204864 327264 204876
rect 316006 204836 327264 204864
rect 327258 204824 327264 204836
rect 327316 204864 327322 204876
rect 327810 204864 327816 204876
rect 327316 204836 327816 204864
rect 327316 204824 327322 204836
rect 327810 204824 327816 204836
rect 327868 204824 327874 204876
rect 247954 203600 247960 203652
rect 248012 203640 248018 203652
rect 332594 203640 332600 203652
rect 248012 203612 332600 203640
rect 248012 203600 248018 203612
rect 332594 203600 332600 203612
rect 332652 203600 332658 203652
rect 229002 203532 229008 203584
rect 229060 203572 229066 203584
rect 342254 203572 342260 203584
rect 229060 203544 342260 203572
rect 229060 203532 229066 203544
rect 342254 203532 342260 203544
rect 342312 203532 342318 203584
rect 3326 202784 3332 202836
rect 3384 202824 3390 202836
rect 159266 202824 159272 202836
rect 3384 202796 159272 202824
rect 3384 202784 3390 202796
rect 159266 202784 159272 202796
rect 159324 202784 159330 202836
rect 208946 202104 208952 202156
rect 209004 202144 209010 202156
rect 266722 202144 266728 202156
rect 209004 202116 266728 202144
rect 209004 202104 209010 202116
rect 266722 202104 266728 202116
rect 266780 202104 266786 202156
rect 210510 200744 210516 200796
rect 210568 200784 210574 200796
rect 224586 200784 224592 200796
rect 210568 200756 224592 200784
rect 210568 200744 210574 200756
rect 224586 200744 224592 200756
rect 224644 200744 224650 200796
rect 210694 199384 210700 199436
rect 210752 199424 210758 199436
rect 225138 199424 225144 199436
rect 210752 199396 225144 199424
rect 210752 199384 210758 199396
rect 225138 199384 225144 199396
rect 225196 199384 225202 199436
rect 577498 193128 577504 193180
rect 577556 193168 577562 193180
rect 579614 193168 579620 193180
rect 577556 193140 579620 193168
rect 577556 193128 577562 193140
rect 579614 193128 579620 193140
rect 579672 193128 579678 193180
rect 3142 188980 3148 189032
rect 3200 189020 3206 189032
rect 160554 189020 160560 189032
rect 3200 188992 160560 189020
rect 3200 188980 3206 188992
rect 160554 188980 160560 188992
rect 160612 188980 160618 189032
rect 257522 187688 257528 187740
rect 257580 187728 257586 187740
rect 257798 187728 257804 187740
rect 257580 187700 257804 187728
rect 257580 187688 257586 187700
rect 257798 187688 257804 187700
rect 257856 187728 257862 187740
rect 449894 187728 449900 187740
rect 257856 187700 449900 187728
rect 257856 187688 257862 187700
rect 449894 187688 449900 187700
rect 449952 187688 449958 187740
rect 257614 186328 257620 186380
rect 257672 186368 257678 186380
rect 257982 186368 257988 186380
rect 257672 186340 257988 186368
rect 257672 186328 257678 186340
rect 257982 186328 257988 186340
rect 258040 186368 258046 186380
rect 447134 186368 447140 186380
rect 258040 186340 447140 186368
rect 258040 186328 258046 186340
rect 447134 186328 447140 186340
rect 447192 186328 447198 186380
rect 242618 184152 242624 184204
rect 242676 184192 242682 184204
rect 260834 184192 260840 184204
rect 242676 184164 260840 184192
rect 242676 184152 242682 184164
rect 260834 184152 260840 184164
rect 260892 184152 260898 184204
rect 256234 183540 256240 183592
rect 256292 183580 256298 183592
rect 256510 183580 256516 183592
rect 256292 183552 256516 183580
rect 256292 183540 256298 183552
rect 256510 183540 256516 183552
rect 256568 183580 256574 183592
rect 425054 183580 425060 183592
rect 256568 183552 425060 183580
rect 256568 183540 256574 183552
rect 425054 183540 425060 183552
rect 425112 183540 425118 183592
rect 210326 180072 210332 180124
rect 210384 180112 210390 180124
rect 222286 180112 222292 180124
rect 210384 180084 222292 180112
rect 210384 180072 210390 180084
rect 222286 180072 222292 180084
rect 222344 180072 222350 180124
rect 209222 175924 209228 175976
rect 209280 175964 209286 175976
rect 267182 175964 267188 175976
rect 209280 175936 267188 175964
rect 209280 175924 209286 175936
rect 267182 175924 267188 175936
rect 267240 175924 267246 175976
rect 248230 175244 248236 175296
rect 248288 175284 248294 175296
rect 325694 175284 325700 175296
rect 248288 175256 325700 175284
rect 248288 175244 248294 175256
rect 325694 175244 325700 175256
rect 325752 175244 325758 175296
rect 260282 175176 260288 175228
rect 260340 175216 260346 175228
rect 260742 175216 260748 175228
rect 260340 175188 260748 175216
rect 260340 175176 260346 175188
rect 260742 175176 260748 175188
rect 260800 175176 260806 175228
rect 260282 173884 260288 173936
rect 260340 173924 260346 173936
rect 478874 173924 478880 173936
rect 260340 173896 478880 173924
rect 260340 173884 260346 173896
rect 478874 173884 478880 173896
rect 478932 173884 478938 173936
rect 246758 171096 246764 171148
rect 246816 171136 246822 171148
rect 304994 171136 305000 171148
rect 246816 171108 305000 171136
rect 246816 171096 246822 171108
rect 304994 171096 305000 171108
rect 305052 171096 305058 171148
rect 245010 168376 245016 168428
rect 245068 168416 245074 168428
rect 245286 168416 245292 168428
rect 245068 168388 245292 168416
rect 245068 168376 245074 168388
rect 245286 168376 245292 168388
rect 245344 168416 245350 168428
rect 298094 168416 298100 168428
rect 245344 168388 298100 168416
rect 245344 168376 245350 168388
rect 298094 168376 298100 168388
rect 298152 168376 298158 168428
rect 283650 167016 283656 167068
rect 283708 167056 283714 167068
rect 284110 167056 284116 167068
rect 283708 167028 284116 167056
rect 283708 167016 283714 167028
rect 284110 167016 284116 167028
rect 284168 167056 284174 167068
rect 340874 167056 340880 167068
rect 284168 167028 340880 167056
rect 284168 167016 284174 167028
rect 340874 167016 340880 167028
rect 340932 167016 340938 167068
rect 3326 164160 3332 164212
rect 3384 164200 3390 164212
rect 160646 164200 160652 164212
rect 3384 164172 160652 164200
rect 3384 164160 3390 164172
rect 160646 164160 160652 164172
rect 160704 164160 160710 164212
rect 157794 162256 157800 162308
rect 157852 162296 157858 162308
rect 158070 162296 158076 162308
rect 157852 162268 158076 162296
rect 157852 162256 157858 162268
rect 158070 162256 158076 162268
rect 158128 162256 158134 162308
rect 161658 161508 161664 161560
rect 161716 161548 161722 161560
rect 162394 161548 162400 161560
rect 161716 161520 162400 161548
rect 161716 161508 161722 161520
rect 162394 161508 162400 161520
rect 162452 161508 162458 161560
rect 208394 161412 208400 161424
rect 182146 161384 208400 161412
rect 158714 161100 158720 161152
rect 158772 161140 158778 161152
rect 159634 161140 159640 161152
rect 158772 161112 159640 161140
rect 158772 161100 158778 161112
rect 159634 161100 159640 161112
rect 159692 161100 159698 161152
rect 182146 161140 182174 161384
rect 208394 161372 208400 161384
rect 208452 161372 208458 161424
rect 229554 161276 229560 161288
rect 169404 161112 182174 161140
rect 191806 161248 229560 161276
rect 155862 160624 155868 160676
rect 155920 160664 155926 160676
rect 162118 160664 162124 160676
rect 155920 160636 162124 160664
rect 155920 160624 155926 160636
rect 162118 160624 162124 160636
rect 162176 160624 162182 160676
rect 155494 160420 155500 160472
rect 155552 160460 155558 160472
rect 155552 160432 165200 160460
rect 155552 160420 155558 160432
rect 157058 160216 157064 160268
rect 157116 160256 157122 160268
rect 165172 160256 165200 160432
rect 157116 160228 163176 160256
rect 165172 160228 167776 160256
rect 157116 160216 157122 160228
rect 161842 160148 161848 160200
rect 161900 160188 161906 160200
rect 163148 160188 163176 160228
rect 161900 160160 163084 160188
rect 163148 160160 164234 160188
rect 161900 160148 161906 160160
rect 163056 160120 163084 160160
rect 163056 160092 163544 160120
rect 159910 160012 159916 160064
rect 159968 160052 159974 160064
rect 159968 160024 163360 160052
rect 159968 160012 159974 160024
rect 162118 159944 162124 159996
rect 162176 159984 162182 159996
rect 162176 159956 162992 159984
rect 162176 159944 162182 159956
rect 162964 159928 162992 159956
rect 163332 159928 163360 160024
rect 161750 159876 161756 159928
rect 161808 159916 161814 159928
rect 162670 159916 162676 159928
rect 161808 159888 162440 159916
rect 161808 159876 161814 159888
rect 150434 159808 150440 159860
rect 150492 159848 150498 159860
rect 159542 159848 159548 159860
rect 150492 159820 159548 159848
rect 150492 159808 150498 159820
rect 159542 159808 159548 159820
rect 159600 159848 159606 159860
rect 159910 159848 159916 159860
rect 159600 159820 159916 159848
rect 159600 159808 159606 159820
rect 159910 159808 159916 159820
rect 159968 159808 159974 159860
rect 162412 159848 162440 159888
rect 162596 159888 162676 159916
rect 162596 159848 162624 159888
rect 162670 159876 162676 159888
rect 162728 159876 162734 159928
rect 162946 159876 162952 159928
rect 163004 159876 163010 159928
rect 163314 159876 163320 159928
rect 163372 159876 163378 159928
rect 162412 159820 162624 159848
rect 163130 159808 163136 159860
rect 163188 159848 163194 159860
rect 163516 159848 163544 160092
rect 164206 159860 164234 160160
rect 164712 159956 167684 159984
rect 163188 159820 163544 159848
rect 163188 159808 163194 159820
rect 164142 159808 164148 159860
rect 164200 159820 164234 159860
rect 164200 159808 164206 159820
rect 164418 159808 164424 159860
rect 164476 159848 164482 159860
rect 164712 159848 164740 159956
rect 165522 159916 165528 159928
rect 164476 159820 164740 159848
rect 164476 159808 164482 159820
rect 164712 159792 164740 159820
rect 165448 159888 165528 159916
rect 132494 159740 132500 159792
rect 132552 159780 132558 159792
rect 132552 159752 164648 159780
rect 132552 159740 132558 159752
rect 135254 159672 135260 159724
rect 135312 159712 135318 159724
rect 164620 159712 164648 159752
rect 164694 159740 164700 159792
rect 164752 159740 164758 159792
rect 165338 159740 165344 159792
rect 165396 159780 165402 159792
rect 165448 159780 165476 159888
rect 165522 159876 165528 159888
rect 165580 159876 165586 159928
rect 166166 159808 166172 159860
rect 166224 159808 166230 159860
rect 167656 159848 167684 159956
rect 167748 159928 167776 160228
rect 167730 159876 167736 159928
rect 167788 159876 167794 159928
rect 169404 159848 169432 161112
rect 191806 160936 191834 161248
rect 229554 161236 229560 161248
rect 229612 161236 229618 161288
rect 207934 161168 207940 161220
rect 207992 161208 207998 161220
rect 208302 161208 208308 161220
rect 207992 161180 208308 161208
rect 207992 161168 207998 161180
rect 208302 161168 208308 161180
rect 208360 161168 208366 161220
rect 207474 161100 207480 161152
rect 207532 161140 207538 161152
rect 256142 161140 256148 161152
rect 207532 161112 256148 161140
rect 207532 161100 207538 161112
rect 256142 161100 256148 161112
rect 256200 161100 256206 161152
rect 207934 161032 207940 161084
rect 207992 161072 207998 161084
rect 254854 161072 254860 161084
rect 207992 161044 254860 161072
rect 207992 161032 207998 161044
rect 254854 161032 254860 161044
rect 254912 161032 254918 161084
rect 209222 160964 209228 161016
rect 209280 161004 209286 161016
rect 246298 161004 246304 161016
rect 209280 160976 246304 161004
rect 209280 160964 209286 160976
rect 246298 160964 246304 160976
rect 246356 160964 246362 161016
rect 169772 160908 191834 160936
rect 169772 159928 169800 160908
rect 208394 160896 208400 160948
rect 208452 160936 208458 160948
rect 224494 160936 224500 160948
rect 208452 160908 224500 160936
rect 208452 160896 208458 160908
rect 224494 160896 224500 160908
rect 224552 160896 224558 160948
rect 227438 160800 227444 160812
rect 205606 160772 227444 160800
rect 179524 160704 186820 160732
rect 179524 160664 179552 160704
rect 179432 160636 179552 160664
rect 179616 160636 183554 160664
rect 179432 160120 179460 160636
rect 169864 160092 179460 160120
rect 169754 159876 169760 159928
rect 169812 159876 169818 159928
rect 167656 159820 169432 159848
rect 165396 159752 165476 159780
rect 165396 159740 165402 159752
rect 165614 159740 165620 159792
rect 165672 159780 165678 159792
rect 166184 159780 166212 159808
rect 165672 159752 166212 159780
rect 165672 159740 165678 159752
rect 167546 159740 167552 159792
rect 167604 159780 167610 159792
rect 169864 159780 169892 160092
rect 173866 160024 176424 160052
rect 173866 159984 173894 160024
rect 172992 159956 173894 159984
rect 167604 159752 169892 159780
rect 170600 159888 172008 159916
rect 167604 159740 167610 159752
rect 135312 159684 164234 159712
rect 164620 159684 165292 159712
rect 135312 159672 135318 159684
rect 139394 159604 139400 159656
rect 139452 159644 139458 159656
rect 158438 159644 158444 159656
rect 139452 159616 158444 159644
rect 139452 159604 139458 159616
rect 158438 159604 158444 159616
rect 158496 159644 158502 159656
rect 158496 159616 159956 159644
rect 158496 159604 158502 159616
rect 125594 159536 125600 159588
rect 125652 159576 125658 159588
rect 159928 159576 159956 159616
rect 160002 159604 160008 159656
rect 160060 159644 160066 159656
rect 163038 159644 163044 159656
rect 160060 159616 163044 159644
rect 160060 159604 160066 159616
rect 163038 159604 163044 159616
rect 163096 159644 163102 159656
rect 163682 159644 163688 159656
rect 163096 159616 163688 159644
rect 163096 159604 163102 159616
rect 163682 159604 163688 159616
rect 163740 159604 163746 159656
rect 164206 159644 164234 159684
rect 165264 159644 165292 159684
rect 167454 159672 167460 159724
rect 167512 159712 167518 159724
rect 167730 159712 167736 159724
rect 167512 159684 167736 159712
rect 167512 159672 167518 159684
rect 167730 159672 167736 159684
rect 167788 159672 167794 159724
rect 170600 159644 170628 159888
rect 171980 159848 172008 159888
rect 172698 159848 172704 159860
rect 171980 159820 172704 159848
rect 172698 159808 172704 159820
rect 172756 159848 172762 159860
rect 172756 159820 172928 159848
rect 172756 159808 172762 159820
rect 172900 159792 172928 159820
rect 170950 159740 170956 159792
rect 171008 159780 171014 159792
rect 171008 159752 171916 159780
rect 171008 159740 171014 159752
rect 170674 159672 170680 159724
rect 170732 159672 170738 159724
rect 171226 159672 171232 159724
rect 171284 159712 171290 159724
rect 171778 159712 171784 159724
rect 171284 159684 171784 159712
rect 171284 159672 171290 159684
rect 171778 159672 171784 159684
rect 171836 159672 171842 159724
rect 171888 159712 171916 159752
rect 172882 159740 172888 159792
rect 172940 159740 172946 159792
rect 172992 159712 173020 159956
rect 176396 159928 176424 160024
rect 171888 159684 173020 159712
rect 173176 159888 176332 159916
rect 164206 159616 165200 159644
rect 165264 159616 170628 159644
rect 164418 159576 164424 159588
rect 125652 159548 157334 159576
rect 159928 159548 164424 159576
rect 125652 159536 125658 159548
rect 96614 159468 96620 159520
rect 96672 159508 96678 159520
rect 156874 159508 156880 159520
rect 96672 159480 156880 159508
rect 96672 159468 96678 159480
rect 156874 159468 156880 159480
rect 156932 159468 156938 159520
rect 78674 159400 78680 159452
rect 78732 159440 78738 159452
rect 152642 159440 152648 159452
rect 78732 159412 152648 159440
rect 78732 159400 78738 159412
rect 152642 159400 152648 159412
rect 152700 159440 152706 159452
rect 152918 159440 152924 159452
rect 152700 159412 152924 159440
rect 152700 159400 152706 159412
rect 152918 159400 152924 159412
rect 152976 159400 152982 159452
rect 157306 159440 157334 159548
rect 164418 159536 164424 159548
rect 164476 159536 164482 159588
rect 165172 159576 165200 159616
rect 170692 159588 170720 159672
rect 173176 159644 173204 159888
rect 174078 159848 174084 159860
rect 173268 159820 174084 159848
rect 173268 159656 173296 159820
rect 174078 159808 174084 159820
rect 174136 159808 174142 159860
rect 174814 159808 174820 159860
rect 174872 159808 174878 159860
rect 176304 159848 176332 159888
rect 176378 159876 176384 159928
rect 176436 159876 176442 159928
rect 177666 159916 177672 159928
rect 177592 159888 177672 159916
rect 177592 159848 177620 159888
rect 177666 159876 177672 159888
rect 177724 159876 177730 159928
rect 176304 159820 177620 159848
rect 177776 159820 178034 159848
rect 173894 159740 173900 159792
rect 173952 159740 173958 159792
rect 171612 159616 173204 159644
rect 168282 159576 168288 159588
rect 165172 159548 168288 159576
rect 168282 159536 168288 159548
rect 168340 159536 168346 159588
rect 170674 159536 170680 159588
rect 170732 159536 170738 159588
rect 161290 159468 161296 159520
rect 161348 159508 161354 159520
rect 171612 159508 171640 159616
rect 173250 159604 173256 159656
rect 173308 159604 173314 159656
rect 173912 159644 173940 159740
rect 173986 159644 173992 159656
rect 173912 159616 173992 159644
rect 173986 159604 173992 159616
rect 174044 159604 174050 159656
rect 174262 159604 174268 159656
rect 174320 159644 174326 159656
rect 174832 159644 174860 159808
rect 177776 159780 177804 159820
rect 174320 159616 174860 159644
rect 174924 159752 177804 159780
rect 178006 159780 178034 159820
rect 178954 159780 178960 159792
rect 178006 159752 178960 159780
rect 174320 159604 174326 159616
rect 171686 159536 171692 159588
rect 171744 159576 171750 159588
rect 174924 159576 174952 159752
rect 178954 159740 178960 159752
rect 179012 159740 179018 159792
rect 179616 159712 179644 160636
rect 183526 160460 183554 160636
rect 186792 160596 186820 160704
rect 205606 160596 205634 160772
rect 227438 160760 227444 160772
rect 227496 160760 227502 160812
rect 230106 160732 230112 160744
rect 186792 160568 205634 160596
rect 229066 160704 230112 160732
rect 229066 160528 229094 160704
rect 230106 160692 230112 160704
rect 230164 160692 230170 160744
rect 205606 160500 229094 160528
rect 183526 160432 195376 160460
rect 195348 160392 195376 160432
rect 205606 160392 205634 160500
rect 195348 160364 205634 160392
rect 209222 160256 209228 160268
rect 191944 160228 209228 160256
rect 186498 159876 186504 159928
rect 186556 159916 186562 159928
rect 191944 159916 191972 160228
rect 209222 160216 209228 160228
rect 209280 160216 209286 160268
rect 209590 160188 209596 160200
rect 192036 160160 198412 160188
rect 192036 159928 192064 160160
rect 193784 160092 197354 160120
rect 193784 159928 193812 160092
rect 186556 159888 191972 159916
rect 186556 159876 186562 159888
rect 192018 159876 192024 159928
rect 192076 159876 192082 159928
rect 193766 159876 193772 159928
rect 193824 159876 193830 159928
rect 197326 159780 197354 160092
rect 198384 159848 198412 160160
rect 200684 160160 208164 160188
rect 200684 159928 200712 160160
rect 207934 160120 207940 160132
rect 203536 160092 207940 160120
rect 199654 159916 199660 159928
rect 199396 159888 199660 159916
rect 198384 159820 198596 159848
rect 198568 159792 198596 159820
rect 199396 159792 199424 159888
rect 199654 159876 199660 159888
rect 199712 159876 199718 159928
rect 200666 159876 200672 159928
rect 200724 159876 200730 159928
rect 203536 159792 203564 160092
rect 207934 160080 207940 160092
rect 207992 160080 207998 160132
rect 208136 160052 208164 160160
rect 208366 160160 209596 160188
rect 208366 160052 208394 160160
rect 209590 160148 209596 160160
rect 209648 160148 209654 160200
rect 208136 160024 208394 160052
rect 208946 159984 208952 159996
rect 206480 159956 208952 159984
rect 206480 159928 206508 159956
rect 208946 159944 208952 159956
rect 209004 159944 209010 159996
rect 206462 159876 206468 159928
rect 206520 159876 206526 159928
rect 206738 159876 206744 159928
rect 206796 159916 206802 159928
rect 208762 159916 208768 159928
rect 206796 159888 208768 159916
rect 206796 159876 206802 159888
rect 208762 159876 208768 159888
rect 208820 159876 208826 159928
rect 205910 159808 205916 159860
rect 205968 159848 205974 159860
rect 207658 159848 207664 159860
rect 205968 159820 207664 159848
rect 205968 159808 205974 159820
rect 207658 159808 207664 159820
rect 207716 159808 207722 159860
rect 197906 159780 197912 159792
rect 197326 159752 197912 159780
rect 197906 159740 197912 159752
rect 197964 159740 197970 159792
rect 198550 159740 198556 159792
rect 198608 159740 198614 159792
rect 199378 159740 199384 159792
rect 199436 159740 199442 159792
rect 203518 159740 203524 159792
rect 203576 159740 203582 159792
rect 203794 159740 203800 159792
rect 203852 159780 203858 159792
rect 209038 159780 209044 159792
rect 203852 159752 209044 159780
rect 203852 159740 203858 159752
rect 209038 159740 209044 159752
rect 209096 159740 209102 159792
rect 207750 159712 207756 159724
rect 171744 159548 174952 159576
rect 175016 159684 179644 159712
rect 183526 159684 207756 159712
rect 171744 159536 171750 159548
rect 175016 159508 175044 159684
rect 183526 159644 183554 159684
rect 207750 159672 207756 159684
rect 207808 159672 207814 159724
rect 177868 159616 183554 159644
rect 161348 159480 171640 159508
rect 171704 159480 175044 159508
rect 161348 159468 161354 159480
rect 158530 159440 158536 159452
rect 157306 159412 158536 159440
rect 158530 159400 158536 159412
rect 158588 159440 158594 159452
rect 165522 159440 165528 159452
rect 158588 159412 165528 159440
rect 158588 159400 158594 159412
rect 165522 159400 165528 159412
rect 165580 159400 165586 159452
rect 166902 159400 166908 159452
rect 166960 159440 166966 159452
rect 167178 159440 167184 159452
rect 166960 159412 167184 159440
rect 166960 159400 166966 159412
rect 167178 159400 167184 159412
rect 167236 159400 167242 159452
rect 169570 159400 169576 159452
rect 169628 159440 169634 159452
rect 171704 159440 171732 159480
rect 175090 159468 175096 159520
rect 175148 159508 175154 159520
rect 177868 159508 177896 159616
rect 185394 159604 185400 159656
rect 185452 159644 185458 159656
rect 208578 159644 208584 159656
rect 185452 159616 208584 159644
rect 185452 159604 185458 159616
rect 208578 159604 208584 159616
rect 208636 159604 208642 159656
rect 182542 159536 182548 159588
rect 182600 159576 182606 159588
rect 242158 159576 242164 159588
rect 182600 159548 242164 159576
rect 182600 159536 182606 159548
rect 242158 159536 242164 159548
rect 242216 159536 242222 159588
rect 175148 159480 177896 159508
rect 175148 159468 175154 159480
rect 178954 159468 178960 159520
rect 179012 159508 179018 159520
rect 179012 159480 186314 159508
rect 179012 159468 179018 159480
rect 173250 159440 173256 159452
rect 169628 159412 171732 159440
rect 172256 159412 173256 159440
rect 169628 159400 169634 159412
rect 3694 159332 3700 159384
rect 3752 159372 3758 159384
rect 157886 159372 157892 159384
rect 3752 159344 157892 159372
rect 3752 159332 3758 159344
rect 157886 159332 157892 159344
rect 157944 159332 157950 159384
rect 159910 159332 159916 159384
rect 159968 159372 159974 159384
rect 172256 159372 172284 159412
rect 173250 159400 173256 159412
rect 173308 159400 173314 159452
rect 159968 159344 165476 159372
rect 159968 159332 159974 159344
rect 164234 159304 164240 159316
rect 157306 159276 164240 159304
rect 154390 159196 154396 159248
rect 154448 159236 154454 159248
rect 157306 159236 157334 159276
rect 164234 159264 164240 159276
rect 164292 159304 164298 159316
rect 165338 159304 165344 159316
rect 164292 159276 165344 159304
rect 164292 159264 164298 159276
rect 165338 159264 165344 159276
rect 165396 159264 165402 159316
rect 165448 159304 165476 159344
rect 165632 159344 172284 159372
rect 165632 159304 165660 159344
rect 172606 159332 172612 159384
rect 172664 159372 172670 159384
rect 173158 159372 173164 159384
rect 172664 159344 173164 159372
rect 172664 159332 172670 159344
rect 173158 159332 173164 159344
rect 173216 159372 173222 159384
rect 181714 159372 181720 159384
rect 173216 159344 181720 159372
rect 173216 159332 173222 159344
rect 181714 159332 181720 159344
rect 181772 159332 181778 159384
rect 186286 159372 186314 159480
rect 190178 159468 190184 159520
rect 190236 159508 190242 159520
rect 211798 159508 211804 159520
rect 190236 159480 211804 159508
rect 190236 159468 190242 159480
rect 211798 159468 211804 159480
rect 211856 159468 211862 159520
rect 195422 159400 195428 159452
rect 195480 159440 195486 159452
rect 219250 159440 219256 159452
rect 195480 159412 219256 159440
rect 195480 159400 195486 159412
rect 219250 159400 219256 159412
rect 219308 159400 219314 159452
rect 210234 159372 210240 159384
rect 186286 159344 210240 159372
rect 210234 159332 210240 159344
rect 210292 159332 210298 159384
rect 167362 159304 167368 159316
rect 165448 159276 165660 159304
rect 165724 159276 167368 159304
rect 154448 159208 157334 159236
rect 154448 159196 154454 159208
rect 161198 159196 161204 159248
rect 161256 159236 161262 159248
rect 161256 159208 163360 159236
rect 161256 159196 161262 159208
rect 161566 159128 161572 159180
rect 161624 159168 161630 159180
rect 162578 159168 162584 159180
rect 161624 159140 162584 159168
rect 161624 159128 161630 159140
rect 162578 159128 162584 159140
rect 162636 159128 162642 159180
rect 163332 159168 163360 159208
rect 164418 159196 164424 159248
rect 164476 159236 164482 159248
rect 165724 159236 165752 159276
rect 167362 159264 167368 159276
rect 167420 159264 167426 159316
rect 167730 159264 167736 159316
rect 167788 159304 167794 159316
rect 167788 159276 201264 159304
rect 167788 159264 167794 159276
rect 164476 159208 165752 159236
rect 164476 159196 164482 159208
rect 166534 159196 166540 159248
rect 166592 159236 166598 159248
rect 201236 159236 201264 159276
rect 201310 159264 201316 159316
rect 201368 159304 201374 159316
rect 208854 159304 208860 159316
rect 201368 159276 208860 159304
rect 201368 159264 201374 159276
rect 208854 159264 208860 159276
rect 208912 159264 208918 159316
rect 203794 159236 203800 159248
rect 166592 159208 200804 159236
rect 201236 159208 203800 159236
rect 166592 159196 166598 159208
rect 163332 159140 170996 159168
rect 153010 159060 153016 159112
rect 153068 159100 153074 159112
rect 161842 159100 161848 159112
rect 153068 159072 161848 159100
rect 153068 159060 153074 159072
rect 161842 159060 161848 159072
rect 161900 159060 161906 159112
rect 168926 159100 168932 159112
rect 162136 159072 168932 159100
rect 152734 158992 152740 159044
rect 152792 159032 152798 159044
rect 162136 159032 162164 159072
rect 168926 159060 168932 159072
rect 168984 159060 168990 159112
rect 170968 159100 170996 159140
rect 171042 159128 171048 159180
rect 171100 159168 171106 159180
rect 171100 159140 181484 159168
rect 171100 159128 171106 159140
rect 176194 159100 176200 159112
rect 170968 159072 176200 159100
rect 176194 159060 176200 159072
rect 176252 159060 176258 159112
rect 176838 159060 176844 159112
rect 176896 159100 176902 159112
rect 178954 159100 178960 159112
rect 176896 159072 178960 159100
rect 176896 159060 176902 159072
rect 178954 159060 178960 159072
rect 179012 159060 179018 159112
rect 168558 159032 168564 159044
rect 152792 159004 162164 159032
rect 162228 159004 168564 159032
rect 152792 158992 152798 159004
rect 152918 158924 152924 158976
rect 152976 158964 152982 158976
rect 162228 158964 162256 159004
rect 168558 158992 168564 159004
rect 168616 158992 168622 159044
rect 170766 158992 170772 159044
rect 170824 159032 170830 159044
rect 170824 159004 181392 159032
rect 170824 158992 170830 159004
rect 152976 158936 162256 158964
rect 152976 158924 152982 158936
rect 163130 158924 163136 158976
rect 163188 158964 163194 158976
rect 163406 158964 163412 158976
rect 163188 158936 163412 158964
rect 163188 158924 163194 158936
rect 163406 158924 163412 158936
rect 163464 158924 163470 158976
rect 164326 158924 164332 158976
rect 164384 158964 164390 158976
rect 165246 158964 165252 158976
rect 164384 158936 165252 158964
rect 164384 158924 164390 158936
rect 165246 158924 165252 158936
rect 165304 158924 165310 158976
rect 167178 158924 167184 158976
rect 167236 158964 167242 158976
rect 169938 158964 169944 158976
rect 167236 158936 169944 158964
rect 167236 158924 167242 158936
rect 169938 158924 169944 158936
rect 169996 158924 170002 158976
rect 171502 158924 171508 158976
rect 171560 158964 171566 158976
rect 172054 158964 172060 158976
rect 171560 158936 172060 158964
rect 171560 158924 171566 158936
rect 172054 158924 172060 158936
rect 172112 158964 172118 158976
rect 175090 158964 175096 158976
rect 172112 158936 175096 158964
rect 172112 158924 172118 158936
rect 175090 158924 175096 158936
rect 175148 158924 175154 158976
rect 161382 158856 161388 158908
rect 161440 158896 161446 158908
rect 178218 158896 178224 158908
rect 161440 158868 178224 158896
rect 161440 158856 161446 158868
rect 178218 158856 178224 158868
rect 178276 158896 178282 158908
rect 178276 158868 179368 158896
rect 178276 158856 178282 158868
rect 161934 158788 161940 158840
rect 161992 158828 161998 158840
rect 176010 158828 176016 158840
rect 161992 158800 176016 158828
rect 161992 158788 161998 158800
rect 176010 158788 176016 158800
rect 176068 158788 176074 158840
rect 164142 158720 164148 158772
rect 164200 158720 164206 158772
rect 164418 158720 164424 158772
rect 164476 158760 164482 158772
rect 164694 158760 164700 158772
rect 164476 158732 164700 158760
rect 164476 158720 164482 158732
rect 164694 158720 164700 158732
rect 164752 158720 164758 158772
rect 166810 158720 166816 158772
rect 166868 158720 166874 158772
rect 172146 158760 172152 158772
rect 166920 158732 172152 158760
rect 154298 158652 154304 158704
rect 154356 158692 154362 158704
rect 164160 158692 164188 158720
rect 154356 158664 157334 158692
rect 154356 158652 154362 158664
rect 157306 158624 157334 158664
rect 163884 158664 164188 158692
rect 163774 158624 163780 158636
rect 157306 158596 163780 158624
rect 163774 158584 163780 158596
rect 163832 158584 163838 158636
rect 163038 158516 163044 158568
rect 163096 158556 163102 158568
rect 163884 158556 163912 158664
rect 164326 158652 164332 158704
rect 164384 158692 164390 158704
rect 166828 158692 166856 158720
rect 164384 158664 166856 158692
rect 164384 158652 164390 158664
rect 164602 158584 164608 158636
rect 164660 158584 164666 158636
rect 165522 158584 165528 158636
rect 165580 158624 165586 158636
rect 166920 158624 166948 158732
rect 172146 158720 172152 158732
rect 172204 158720 172210 158772
rect 169864 158664 170168 158692
rect 165580 158596 166948 158624
rect 165580 158584 165586 158596
rect 169202 158584 169208 158636
rect 169260 158624 169266 158636
rect 169754 158624 169760 158636
rect 169260 158596 169760 158624
rect 169260 158584 169266 158596
rect 169754 158584 169760 158596
rect 169812 158584 169818 158636
rect 163096 158528 163912 158556
rect 163096 158516 163102 158528
rect 164326 158516 164332 158568
rect 164384 158556 164390 158568
rect 164620 158556 164648 158584
rect 169864 158556 169892 158664
rect 170140 158624 170168 158664
rect 172790 158652 172796 158704
rect 172848 158692 172854 158704
rect 173434 158692 173440 158704
rect 172848 158664 173440 158692
rect 172848 158652 172854 158664
rect 173434 158652 173440 158664
rect 173492 158652 173498 158704
rect 176562 158624 176568 158636
rect 170140 158596 176568 158624
rect 176562 158584 176568 158596
rect 176620 158584 176626 158636
rect 176838 158584 176844 158636
rect 176896 158584 176902 158636
rect 177114 158624 177120 158636
rect 177040 158596 177120 158624
rect 172974 158556 172980 158568
rect 164384 158528 164648 158556
rect 165448 158528 169892 158556
rect 170784 158528 172980 158556
rect 164384 158516 164390 158528
rect 162302 158448 162308 158500
rect 162360 158488 162366 158500
rect 165448 158488 165476 158528
rect 162360 158460 165476 158488
rect 162360 158448 162366 158460
rect 168282 158448 168288 158500
rect 168340 158488 168346 158500
rect 170784 158488 170812 158528
rect 172974 158516 172980 158528
rect 173032 158516 173038 158568
rect 176856 158556 176884 158584
rect 173866 158528 176884 158556
rect 173866 158488 173894 158528
rect 168340 158460 170812 158488
rect 170876 158460 173894 158488
rect 168340 158448 168346 158460
rect 151170 158380 151176 158432
rect 151228 158420 151234 158432
rect 151630 158420 151636 158432
rect 151228 158392 151636 158420
rect 151228 158380 151234 158392
rect 151630 158380 151636 158392
rect 151688 158420 151694 158432
rect 165614 158420 165620 158432
rect 151688 158392 165620 158420
rect 151688 158380 151694 158392
rect 165614 158380 165620 158392
rect 165672 158380 165678 158432
rect 167362 158380 167368 158432
rect 167420 158420 167426 158432
rect 170582 158420 170588 158432
rect 167420 158392 170588 158420
rect 167420 158380 167426 158392
rect 170582 158380 170588 158392
rect 170640 158380 170646 158432
rect 153930 158312 153936 158364
rect 153988 158352 153994 158364
rect 164326 158352 164332 158364
rect 153988 158324 164332 158352
rect 153988 158312 153994 158324
rect 164326 158312 164332 158324
rect 164384 158312 164390 158364
rect 165890 158312 165896 158364
rect 165948 158352 165954 158364
rect 166350 158352 166356 158364
rect 165948 158324 166356 158352
rect 165948 158312 165954 158324
rect 166350 158312 166356 158324
rect 166408 158312 166414 158364
rect 170876 158352 170904 158460
rect 176838 158448 176844 158500
rect 176896 158488 176902 158500
rect 177040 158488 177068 158596
rect 177114 158584 177120 158596
rect 177172 158584 177178 158636
rect 179340 158624 179368 158868
rect 181364 158828 181392 159004
rect 181456 158964 181484 159140
rect 190822 159128 190828 159180
rect 190880 159168 190886 159180
rect 191282 159168 191288 159180
rect 190880 159140 191288 159168
rect 190880 159128 190886 159140
rect 191282 159128 191288 159140
rect 191340 159128 191346 159180
rect 195514 159128 195520 159180
rect 195572 159168 195578 159180
rect 200666 159168 200672 159180
rect 195572 159140 200672 159168
rect 195572 159128 195578 159140
rect 200666 159128 200672 159140
rect 200724 159128 200730 159180
rect 200776 159168 200804 159208
rect 203794 159196 203800 159208
rect 203852 159196 203858 159248
rect 204530 159196 204536 159248
rect 204588 159236 204594 159248
rect 204588 159208 209774 159236
rect 204588 159196 204594 159208
rect 201310 159168 201316 159180
rect 200776 159140 201316 159168
rect 201310 159128 201316 159140
rect 201368 159128 201374 159180
rect 202322 159128 202328 159180
rect 202380 159168 202386 159180
rect 203426 159168 203432 159180
rect 202380 159140 203432 159168
rect 202380 159128 202386 159140
rect 203426 159128 203432 159140
rect 203484 159128 203490 159180
rect 205082 159128 205088 159180
rect 205140 159168 205146 159180
rect 205542 159168 205548 159180
rect 205140 159140 205548 159168
rect 205140 159128 205146 159140
rect 205542 159128 205548 159140
rect 205600 159128 205606 159180
rect 206738 159128 206744 159180
rect 206796 159168 206802 159180
rect 207474 159168 207480 159180
rect 206796 159140 207480 159168
rect 206796 159128 206802 159140
rect 207474 159128 207480 159140
rect 207532 159128 207538 159180
rect 207750 159128 207756 159180
rect 207808 159168 207814 159180
rect 209222 159168 209228 159180
rect 207808 159140 209228 159168
rect 207808 159128 207814 159140
rect 209222 159128 209228 159140
rect 209280 159128 209286 159180
rect 209746 159168 209774 159208
rect 264238 159168 264244 159180
rect 209746 159140 264244 159168
rect 264238 159128 264244 159140
rect 264296 159128 264302 159180
rect 181714 159060 181720 159112
rect 181772 159100 181778 159112
rect 232866 159100 232872 159112
rect 181772 159072 232872 159100
rect 181772 159060 181778 159072
rect 232866 159060 232872 159072
rect 232924 159060 232930 159112
rect 181898 158992 181904 159044
rect 181956 159032 181962 159044
rect 232498 159032 232504 159044
rect 181956 159004 232504 159032
rect 181956 158992 181962 159004
rect 232498 158992 232504 159004
rect 232556 158992 232562 159044
rect 229922 158964 229928 158976
rect 181456 158936 229928 158964
rect 229922 158924 229928 158936
rect 229980 158924 229986 158976
rect 184198 158856 184204 158908
rect 184256 158896 184262 158908
rect 243630 158896 243636 158908
rect 184256 158868 243636 158896
rect 184256 158856 184262 158868
rect 243630 158856 243636 158868
rect 243688 158856 243694 158908
rect 181364 158800 188384 158828
rect 182358 158720 182364 158772
rect 182416 158760 182422 158772
rect 183278 158760 183284 158772
rect 182416 158732 183284 158760
rect 182416 158720 182422 158732
rect 183278 158720 183284 158732
rect 183336 158720 183342 158772
rect 183646 158720 183652 158772
rect 183704 158760 183710 158772
rect 184198 158760 184204 158772
rect 183704 158732 184204 158760
rect 183704 158720 183710 158732
rect 184198 158720 184204 158732
rect 184256 158720 184262 158772
rect 188356 158760 188384 158800
rect 189350 158788 189356 158840
rect 189408 158828 189414 158840
rect 189626 158828 189632 158840
rect 189408 158800 189632 158828
rect 189408 158788 189414 158800
rect 189626 158788 189632 158800
rect 189684 158788 189690 158840
rect 196158 158788 196164 158840
rect 196216 158828 196222 158840
rect 197170 158828 197176 158840
rect 196216 158800 197176 158828
rect 196216 158788 196222 158800
rect 197170 158788 197176 158800
rect 197228 158788 197234 158840
rect 198550 158788 198556 158840
rect 198608 158828 198614 158840
rect 199654 158828 199660 158840
rect 198608 158800 199660 158828
rect 198608 158788 198614 158800
rect 199654 158788 199660 158800
rect 199712 158788 199718 158840
rect 200666 158788 200672 158840
rect 200724 158828 200730 158840
rect 256234 158828 256240 158840
rect 200724 158800 256240 158828
rect 200724 158788 200730 158800
rect 256234 158788 256240 158800
rect 256292 158788 256298 158840
rect 231486 158760 231492 158772
rect 188356 158732 231492 158760
rect 231486 158720 231492 158732
rect 231544 158720 231550 158772
rect 182266 158652 182272 158704
rect 182324 158692 182330 158704
rect 183462 158692 183468 158704
rect 182324 158664 183468 158692
rect 182324 158652 182330 158664
rect 183462 158652 183468 158664
rect 183520 158652 183526 158704
rect 184382 158652 184388 158704
rect 184440 158692 184446 158704
rect 186314 158692 186320 158704
rect 184440 158664 186320 158692
rect 184440 158652 184446 158664
rect 186314 158652 186320 158664
rect 186372 158652 186378 158704
rect 188246 158652 188252 158704
rect 188304 158692 188310 158704
rect 189350 158692 189356 158704
rect 188304 158664 189356 158692
rect 188304 158652 188310 158664
rect 189350 158652 189356 158664
rect 189408 158652 189414 158704
rect 189902 158652 189908 158704
rect 189960 158692 189966 158704
rect 194410 158692 194416 158704
rect 189960 158664 194416 158692
rect 189960 158652 189966 158664
rect 194410 158652 194416 158664
rect 194468 158652 194474 158704
rect 195146 158652 195152 158704
rect 195204 158692 195210 158704
rect 196618 158692 196624 158704
rect 195204 158664 196624 158692
rect 195204 158652 195210 158664
rect 196618 158652 196624 158664
rect 196676 158652 196682 158704
rect 200022 158652 200028 158704
rect 200080 158692 200086 158704
rect 202322 158692 202328 158704
rect 200080 158664 202328 158692
rect 200080 158652 200086 158664
rect 202322 158652 202328 158664
rect 202380 158652 202386 158704
rect 202874 158652 202880 158704
rect 202932 158692 202938 158704
rect 203334 158692 203340 158704
rect 202932 158664 203340 158692
rect 202932 158652 202938 158664
rect 203334 158652 203340 158664
rect 203392 158652 203398 158704
rect 206738 158692 206744 158704
rect 203628 158664 206744 158692
rect 184750 158624 184756 158636
rect 179340 158596 184756 158624
rect 184750 158584 184756 158596
rect 184808 158584 184814 158636
rect 186866 158584 186872 158636
rect 186924 158624 186930 158636
rect 188522 158624 188528 158636
rect 186924 158596 188528 158624
rect 186924 158584 186930 158596
rect 188522 158584 188528 158596
rect 188580 158584 188586 158636
rect 194318 158584 194324 158636
rect 194376 158624 194382 158636
rect 203518 158624 203524 158636
rect 194376 158596 203524 158624
rect 194376 158584 194382 158596
rect 203518 158584 203524 158596
rect 203576 158584 203582 158636
rect 187142 158516 187148 158568
rect 187200 158556 187206 158568
rect 189902 158556 189908 158568
rect 187200 158528 189908 158556
rect 187200 158516 187206 158528
rect 189902 158516 189908 158528
rect 189960 158516 189966 158568
rect 190178 158516 190184 158568
rect 190236 158556 190242 158568
rect 201310 158556 201316 158568
rect 190236 158528 201316 158556
rect 190236 158516 190242 158528
rect 201310 158516 201316 158528
rect 201368 158516 201374 158568
rect 176896 158460 177068 158488
rect 176896 158448 176902 158460
rect 177114 158448 177120 158500
rect 177172 158488 177178 158500
rect 177390 158488 177396 158500
rect 177172 158460 177396 158488
rect 177172 158448 177178 158460
rect 177390 158448 177396 158460
rect 177448 158448 177454 158500
rect 182726 158448 182732 158500
rect 182784 158488 182790 158500
rect 188246 158488 188252 158500
rect 182784 158460 188252 158488
rect 182784 158448 182790 158460
rect 188246 158448 188252 158460
rect 188304 158448 188310 158500
rect 188338 158448 188344 158500
rect 188396 158488 188402 158500
rect 191190 158488 191196 158500
rect 188396 158460 191196 158488
rect 188396 158448 188402 158460
rect 191190 158448 191196 158460
rect 191248 158448 191254 158500
rect 196526 158448 196532 158500
rect 196584 158488 196590 158500
rect 203628 158488 203656 158664
rect 206738 158652 206744 158664
rect 206796 158652 206802 158704
rect 207198 158652 207204 158704
rect 207256 158692 207262 158704
rect 251818 158692 251824 158704
rect 207256 158664 251824 158692
rect 207256 158652 207262 158664
rect 251818 158652 251824 158664
rect 251876 158652 251882 158704
rect 203794 158584 203800 158636
rect 203852 158624 203858 158636
rect 204162 158624 204168 158636
rect 203852 158596 204168 158624
rect 203852 158584 203858 158596
rect 204162 158584 204168 158596
rect 204220 158584 204226 158636
rect 204806 158584 204812 158636
rect 204864 158624 204870 158636
rect 209498 158624 209504 158636
rect 204864 158596 209504 158624
rect 204864 158584 204870 158596
rect 209498 158584 209504 158596
rect 209556 158584 209562 158636
rect 204254 158516 204260 158568
rect 204312 158556 204318 158568
rect 209314 158556 209320 158568
rect 204312 158528 209320 158556
rect 204312 158516 204318 158528
rect 209314 158516 209320 158528
rect 209372 158516 209378 158568
rect 196584 158460 203656 158488
rect 196584 158448 196590 158460
rect 203702 158448 203708 158500
rect 203760 158488 203766 158500
rect 247678 158488 247684 158500
rect 203760 158460 247684 158488
rect 203760 158448 203766 158460
rect 247678 158448 247684 158460
rect 247736 158448 247742 158500
rect 172606 158380 172612 158432
rect 172664 158420 172670 158432
rect 172664 158392 176608 158420
rect 172664 158380 172670 158392
rect 166460 158324 170904 158352
rect 148318 158244 148324 158296
rect 148376 158284 148382 158296
rect 160554 158284 160560 158296
rect 148376 158256 160560 158284
rect 148376 158244 148382 158256
rect 160554 158244 160560 158256
rect 160612 158244 160618 158296
rect 162210 158244 162216 158296
rect 162268 158284 162274 158296
rect 166460 158284 166488 158324
rect 171686 158312 171692 158364
rect 171744 158352 171750 158364
rect 172054 158352 172060 158364
rect 171744 158324 172060 158352
rect 171744 158312 171750 158324
rect 172054 158312 172060 158324
rect 172112 158312 172118 158364
rect 174630 158312 174636 158364
rect 174688 158352 174694 158364
rect 175550 158352 175556 158364
rect 174688 158324 175556 158352
rect 174688 158312 174694 158324
rect 175550 158312 175556 158324
rect 175608 158312 175614 158364
rect 176580 158352 176608 158392
rect 176856 158392 200896 158420
rect 176856 158352 176884 158392
rect 176580 158324 176884 158352
rect 176948 158324 200528 158352
rect 162268 158256 166488 158284
rect 162268 158244 162274 158256
rect 166718 158244 166724 158296
rect 166776 158284 166782 158296
rect 172330 158284 172336 158296
rect 166776 158256 172336 158284
rect 166776 158244 166782 158256
rect 172330 158244 172336 158256
rect 172388 158244 172394 158296
rect 166902 158216 166908 158228
rect 164068 158188 166908 158216
rect 124858 158108 124864 158160
rect 124916 158148 124922 158160
rect 163958 158148 163964 158160
rect 124916 158120 163964 158148
rect 124916 158108 124922 158120
rect 163958 158108 163964 158120
rect 164016 158108 164022 158160
rect 60734 158040 60740 158092
rect 60792 158080 60798 158092
rect 164068 158080 164096 158188
rect 166902 158176 166908 158188
rect 166960 158176 166966 158228
rect 168282 158176 168288 158228
rect 168340 158216 168346 158228
rect 172422 158216 172428 158228
rect 168340 158188 172428 158216
rect 168340 158176 168346 158188
rect 172422 158176 172428 158188
rect 172480 158176 172486 158228
rect 171226 158108 171232 158160
rect 171284 158148 171290 158160
rect 171502 158148 171508 158160
rect 171284 158120 171508 158148
rect 171284 158108 171290 158120
rect 171502 158108 171508 158120
rect 171560 158148 171566 158160
rect 171560 158120 173894 158148
rect 171560 158108 171566 158120
rect 60792 158052 164096 158080
rect 60792 158040 60798 158052
rect 169754 158040 169760 158092
rect 169812 158080 169818 158092
rect 170122 158080 170128 158092
rect 169812 158052 170128 158080
rect 169812 158040 169818 158052
rect 170122 158040 170128 158052
rect 170180 158080 170186 158092
rect 172606 158080 172612 158092
rect 170180 158052 172612 158080
rect 170180 158040 170186 158052
rect 172606 158040 172612 158052
rect 172664 158040 172670 158092
rect 173866 158080 173894 158120
rect 176948 158080 176976 158324
rect 186314 158244 186320 158296
rect 186372 158284 186378 158296
rect 192018 158284 192024 158296
rect 186372 158256 192024 158284
rect 186372 158244 186378 158256
rect 192018 158244 192024 158256
rect 192076 158244 192082 158296
rect 177390 158176 177396 158228
rect 177448 158216 177454 158228
rect 177666 158216 177672 158228
rect 177448 158188 177672 158216
rect 177448 158176 177454 158188
rect 177666 158176 177672 158188
rect 177724 158176 177730 158228
rect 184106 158176 184112 158228
rect 184164 158216 184170 158228
rect 197998 158216 198004 158228
rect 184164 158188 198004 158216
rect 184164 158176 184170 158188
rect 197998 158176 198004 158188
rect 198056 158176 198062 158228
rect 181346 158108 181352 158160
rect 181404 158148 181410 158160
rect 190270 158148 190276 158160
rect 181404 158120 190276 158148
rect 181404 158108 181410 158120
rect 190270 158108 190276 158120
rect 190328 158108 190334 158160
rect 191006 158108 191012 158160
rect 191064 158148 191070 158160
rect 191064 158120 191512 158148
rect 191064 158108 191070 158120
rect 173866 158052 176976 158080
rect 180518 158040 180524 158092
rect 180576 158080 180582 158092
rect 191098 158080 191104 158092
rect 180576 158052 191104 158080
rect 180576 158040 180582 158052
rect 191098 158040 191104 158052
rect 191156 158040 191162 158092
rect 46198 157972 46204 158024
rect 46256 158012 46262 158024
rect 161474 158012 161480 158024
rect 46256 157984 161480 158012
rect 46256 157972 46262 157984
rect 161474 157972 161480 157984
rect 161532 158012 161538 158024
rect 162762 158012 162768 158024
rect 161532 157984 162768 158012
rect 161532 157972 161538 157984
rect 162762 157972 162768 157984
rect 162820 157972 162826 158024
rect 163498 157972 163504 158024
rect 163556 158012 163562 158024
rect 174262 158012 174268 158024
rect 163556 157984 174268 158012
rect 163556 157972 163562 157984
rect 174262 157972 174268 157984
rect 174320 157972 174326 158024
rect 180242 157972 180248 158024
rect 180300 158012 180306 158024
rect 190178 158012 190184 158024
rect 180300 157984 190184 158012
rect 180300 157972 180306 157984
rect 190178 157972 190184 157984
rect 190236 157972 190242 158024
rect 156690 157904 156696 157956
rect 156748 157944 156754 157956
rect 165154 157944 165160 157956
rect 156748 157916 165160 157944
rect 156748 157904 156754 157916
rect 165154 157904 165160 157916
rect 165212 157904 165218 157956
rect 168926 157904 168932 157956
rect 168984 157944 168990 157956
rect 169294 157944 169300 157956
rect 168984 157916 169300 157944
rect 168984 157904 168990 157916
rect 169294 157904 169300 157916
rect 169352 157904 169358 157956
rect 169478 157904 169484 157956
rect 169536 157944 169542 157956
rect 176102 157944 176108 157956
rect 169536 157916 176108 157944
rect 169536 157904 169542 157916
rect 176102 157904 176108 157916
rect 176160 157904 176166 157956
rect 178954 157904 178960 157956
rect 179012 157944 179018 157956
rect 184106 157944 184112 157956
rect 179012 157916 184112 157944
rect 179012 157904 179018 157916
rect 184106 157904 184112 157916
rect 184164 157904 184170 157956
rect 184750 157904 184756 157956
rect 184808 157944 184814 157956
rect 186498 157944 186504 157956
rect 184808 157916 186504 157944
rect 184808 157904 184814 157916
rect 186498 157904 186504 157916
rect 186556 157904 186562 157956
rect 160830 157836 160836 157888
rect 160888 157876 160894 157888
rect 164234 157876 164240 157888
rect 160888 157848 164240 157876
rect 160888 157836 160894 157848
rect 164234 157836 164240 157848
rect 164292 157836 164298 157888
rect 165338 157836 165344 157888
rect 165396 157876 165402 157888
rect 177114 157876 177120 157888
rect 165396 157848 177120 157876
rect 165396 157836 165402 157848
rect 177114 157836 177120 157848
rect 177172 157836 177178 157888
rect 191484 157876 191512 158120
rect 193490 158108 193496 158160
rect 193548 158148 193554 158160
rect 193548 158120 200436 158148
rect 193548 158108 193554 158120
rect 192662 158040 192668 158092
rect 192720 158080 192726 158092
rect 196342 158080 196348 158092
rect 192720 158052 196348 158080
rect 192720 158040 192726 158052
rect 196342 158040 196348 158052
rect 196400 158040 196406 158092
rect 192110 157972 192116 158024
rect 192168 158012 192174 158024
rect 194134 158012 194140 158024
rect 192168 157984 194140 158012
rect 192168 157972 192174 157984
rect 194134 157972 194140 157984
rect 194192 157972 194198 158024
rect 191558 157904 191564 157956
rect 191616 157944 191622 157956
rect 191616 157916 195974 157944
rect 191616 157904 191622 157916
rect 195606 157876 195612 157888
rect 191484 157848 195612 157876
rect 195606 157836 195612 157848
rect 195664 157836 195670 157888
rect 162026 157768 162032 157820
rect 162084 157808 162090 157820
rect 179046 157808 179052 157820
rect 162084 157780 179052 157808
rect 162084 157768 162090 157780
rect 179046 157768 179052 157780
rect 179104 157768 179110 157820
rect 185210 157768 185216 157820
rect 185268 157808 185274 157820
rect 190178 157808 190184 157820
rect 185268 157780 190184 157808
rect 185268 157768 185274 157780
rect 190178 157768 190184 157780
rect 190236 157768 190242 157820
rect 190270 157768 190276 157820
rect 190328 157808 190334 157820
rect 195422 157808 195428 157820
rect 190328 157780 195428 157808
rect 190328 157768 190334 157780
rect 195422 157768 195428 157780
rect 195480 157768 195486 157820
rect 161014 157700 161020 157752
rect 161072 157740 161078 157752
rect 176838 157740 176844 157752
rect 161072 157712 176844 157740
rect 161072 157700 161078 157712
rect 176838 157700 176844 157712
rect 176896 157740 176902 157752
rect 177666 157740 177672 157752
rect 176896 157712 177672 157740
rect 176896 157700 176902 157712
rect 177666 157700 177672 157712
rect 177724 157700 177730 157752
rect 188246 157700 188252 157752
rect 188304 157740 188310 157752
rect 195330 157740 195336 157752
rect 188304 157712 195336 157740
rect 188304 157700 188310 157712
rect 195330 157700 195336 157712
rect 195388 157700 195394 157752
rect 195946 157740 195974 157916
rect 197354 157836 197360 157888
rect 197412 157876 197418 157888
rect 200206 157876 200212 157888
rect 197412 157848 200212 157876
rect 197412 157836 197418 157848
rect 200206 157836 200212 157848
rect 200264 157836 200270 157888
rect 200408 157876 200436 158120
rect 200500 157944 200528 158324
rect 200868 158216 200896 158392
rect 201770 158380 201776 158432
rect 201828 158420 201834 158432
rect 209682 158420 209688 158432
rect 201828 158392 209688 158420
rect 201828 158380 201834 158392
rect 209682 158380 209688 158392
rect 209740 158380 209746 158432
rect 200942 158312 200948 158364
rect 201000 158352 201006 158364
rect 210694 158352 210700 158364
rect 201000 158324 210700 158352
rect 201000 158312 201006 158324
rect 210694 158312 210700 158324
rect 210752 158312 210758 158364
rect 207474 158244 207480 158296
rect 207532 158284 207538 158296
rect 252002 158284 252008 158296
rect 207532 158256 252008 158284
rect 207532 158244 207538 158256
rect 252002 158244 252008 158256
rect 252060 158244 252066 158296
rect 200868 158188 205634 158216
rect 205606 158080 205634 158188
rect 207566 158176 207572 158228
rect 207624 158216 207630 158228
rect 252094 158216 252100 158228
rect 207624 158188 252100 158216
rect 207624 158176 207630 158188
rect 252094 158176 252100 158188
rect 252152 158176 252158 158228
rect 207014 158108 207020 158160
rect 207072 158148 207078 158160
rect 253198 158148 253204 158160
rect 207072 158120 253204 158148
rect 207072 158108 207078 158120
rect 253198 158108 253204 158120
rect 253256 158108 253262 158160
rect 207842 158080 207848 158092
rect 205606 158052 207848 158080
rect 207842 158040 207848 158052
rect 207900 158040 207906 158092
rect 207934 158040 207940 158092
rect 207992 158080 207998 158092
rect 208302 158080 208308 158092
rect 207992 158052 208308 158080
rect 207992 158040 207998 158052
rect 208302 158040 208308 158052
rect 208360 158040 208366 158092
rect 208394 158040 208400 158092
rect 208452 158080 208458 158092
rect 272242 158080 272248 158092
rect 208452 158052 272248 158080
rect 208452 158040 208458 158052
rect 272242 158040 272248 158052
rect 272300 158040 272306 158092
rect 200666 157972 200672 158024
rect 200724 158012 200730 158024
rect 201218 158012 201224 158024
rect 200724 157984 201224 158012
rect 200724 157972 200730 157984
rect 201218 157972 201224 157984
rect 201276 157972 201282 158024
rect 209682 157972 209688 158024
rect 209740 158012 209746 158024
rect 283650 158012 283656 158024
rect 209740 157984 283656 158012
rect 209740 157972 209746 157984
rect 283650 157972 283656 157984
rect 283708 157972 283714 158024
rect 307110 157972 307116 158024
rect 307168 158012 307174 158024
rect 324406 158012 324412 158024
rect 307168 157984 324412 158012
rect 307168 157972 307174 157984
rect 324406 157972 324412 157984
rect 324464 157972 324470 158024
rect 200500 157916 205634 157944
rect 205174 157876 205180 157888
rect 200408 157848 205180 157876
rect 205174 157836 205180 157848
rect 205232 157836 205238 157888
rect 205606 157876 205634 157916
rect 207106 157904 207112 157956
rect 207164 157944 207170 157956
rect 249334 157944 249340 157956
rect 207164 157916 249340 157944
rect 207164 157904 207170 157916
rect 249334 157904 249340 157916
rect 249392 157904 249398 157956
rect 208026 157876 208032 157888
rect 205606 157848 208032 157876
rect 208026 157836 208032 157848
rect 208084 157836 208090 157888
rect 199286 157768 199292 157820
rect 199344 157808 199350 157820
rect 200114 157808 200120 157820
rect 199344 157780 200120 157808
rect 199344 157768 199350 157780
rect 200114 157768 200120 157780
rect 200172 157768 200178 157820
rect 208118 157808 208124 157820
rect 204272 157780 208124 157808
rect 204162 157740 204168 157752
rect 195946 157712 204168 157740
rect 204162 157700 204168 157712
rect 204220 157700 204226 157752
rect 160738 157632 160744 157684
rect 160796 157672 160802 157684
rect 165338 157672 165344 157684
rect 160796 157644 165344 157672
rect 160796 157632 160802 157644
rect 165338 157632 165344 157644
rect 165396 157632 165402 157684
rect 177482 157672 177488 157684
rect 165448 157644 177488 157672
rect 160922 157564 160928 157616
rect 160980 157604 160986 157616
rect 165448 157604 165476 157644
rect 177482 157632 177488 157644
rect 177540 157632 177546 157684
rect 195698 157632 195704 157684
rect 195756 157672 195762 157684
rect 199470 157672 199476 157684
rect 195756 157644 199476 157672
rect 195756 157632 195762 157644
rect 199470 157632 199476 157644
rect 199528 157632 199534 157684
rect 200206 157632 200212 157684
rect 200264 157672 200270 157684
rect 204272 157672 204300 157780
rect 208118 157768 208124 157780
rect 208176 157768 208182 157820
rect 258902 157740 258908 157752
rect 200264 157644 204300 157672
rect 205468 157712 258908 157740
rect 200264 157632 200270 157644
rect 170214 157604 170220 157616
rect 160980 157576 165476 157604
rect 165540 157576 170220 157604
rect 160980 157564 160986 157576
rect 163682 157496 163688 157548
rect 163740 157536 163746 157548
rect 165540 157536 165568 157576
rect 170214 157564 170220 157576
rect 170272 157564 170278 157616
rect 176562 157564 176568 157616
rect 176620 157604 176626 157616
rect 182726 157604 182732 157616
rect 176620 157576 182732 157604
rect 176620 157564 176626 157576
rect 182726 157564 182732 157576
rect 182784 157564 182790 157616
rect 191098 157564 191104 157616
rect 191156 157604 191162 157616
rect 198182 157604 198188 157616
rect 191156 157576 198188 157604
rect 191156 157564 191162 157576
rect 198182 157564 198188 157576
rect 198240 157564 198246 157616
rect 198274 157564 198280 157616
rect 198332 157604 198338 157616
rect 205468 157604 205496 157712
rect 258902 157700 258908 157712
rect 258960 157700 258966 157752
rect 255406 157672 255412 157684
rect 198332 157576 205496 157604
rect 205606 157644 255412 157672
rect 198332 157564 198338 157576
rect 163740 157508 165568 157536
rect 163740 157496 163746 157508
rect 166350 157496 166356 157548
rect 166408 157536 166414 157548
rect 200942 157536 200948 157548
rect 166408 157508 200948 157536
rect 166408 157496 166414 157508
rect 200942 157496 200948 157508
rect 201000 157496 201006 157548
rect 163498 157428 163504 157480
rect 163556 157468 163562 157480
rect 166718 157468 166724 157480
rect 163556 157440 166724 157468
rect 163556 157428 163562 157440
rect 166718 157428 166724 157440
rect 166776 157428 166782 157480
rect 171778 157428 171784 157480
rect 171836 157468 171842 157480
rect 171836 157440 176654 157468
rect 171836 157428 171842 157440
rect 157978 157360 157984 157412
rect 158036 157400 158042 157412
rect 162854 157400 162860 157412
rect 158036 157372 162860 157400
rect 158036 157360 158042 157372
rect 162854 157360 162860 157372
rect 162912 157400 162918 157412
rect 164142 157400 164148 157412
rect 162912 157372 164148 157400
rect 162912 157360 162918 157372
rect 164142 157360 164148 157372
rect 164200 157360 164206 157412
rect 164234 157360 164240 157412
rect 164292 157400 164298 157412
rect 169478 157400 169484 157412
rect 164292 157372 169484 157400
rect 164292 157360 164298 157372
rect 169478 157360 169484 157372
rect 169536 157360 169542 157412
rect 176626 157400 176654 157440
rect 185762 157428 185768 157480
rect 185820 157468 185826 157480
rect 187234 157468 187240 157480
rect 185820 157440 187240 157468
rect 185820 157428 185826 157440
rect 187234 157428 187240 157440
rect 187292 157428 187298 157480
rect 189626 157428 189632 157480
rect 189684 157468 189690 157480
rect 192662 157468 192668 157480
rect 189684 157440 192668 157468
rect 189684 157428 189690 157440
rect 192662 157428 192668 157440
rect 192720 157428 192726 157480
rect 195974 157428 195980 157480
rect 196032 157468 196038 157480
rect 205606 157468 205634 157644
rect 255406 157632 255412 157644
rect 255464 157632 255470 157684
rect 196032 157440 205634 157468
rect 196032 157428 196038 157440
rect 207290 157428 207296 157480
rect 207348 157468 207354 157480
rect 250438 157468 250444 157480
rect 207348 157440 250444 157468
rect 207348 157428 207354 157440
rect 250438 157428 250444 157440
rect 250496 157428 250502 157480
rect 207934 157400 207940 157412
rect 176626 157372 207940 157400
rect 207934 157360 207940 157372
rect 207992 157360 207998 157412
rect 204162 157292 204168 157344
rect 204220 157332 204226 157344
rect 207198 157332 207204 157344
rect 204220 157304 207204 157332
rect 204220 157292 204226 157304
rect 207198 157292 207204 157304
rect 207256 157292 207262 157344
rect 154482 157224 154488 157276
rect 154540 157264 154546 157276
rect 164970 157264 164976 157276
rect 154540 157236 164976 157264
rect 154540 157224 154546 157236
rect 164970 157224 164976 157236
rect 165028 157224 165034 157276
rect 208578 157224 208584 157276
rect 208636 157264 208642 157276
rect 270770 157264 270776 157276
rect 208636 157236 270776 157264
rect 208636 157224 208642 157236
rect 270770 157224 270776 157236
rect 270828 157264 270834 157276
rect 271782 157264 271788 157276
rect 270828 157236 271788 157264
rect 270828 157224 270834 157236
rect 271782 157224 271788 157236
rect 271840 157224 271846 157276
rect 162118 157156 162124 157208
rect 162176 157196 162182 157208
rect 162854 157196 162860 157208
rect 162176 157168 162860 157196
rect 162176 157156 162182 157168
rect 162854 157156 162860 157168
rect 162912 157156 162918 157208
rect 172974 157156 172980 157208
rect 173032 157196 173038 157208
rect 233510 157196 233516 157208
rect 173032 157168 233516 157196
rect 173032 157156 173038 157168
rect 233510 157156 233516 157168
rect 233568 157156 233574 157208
rect 162210 157088 162216 157140
rect 162268 157128 162274 157140
rect 171594 157128 171600 157140
rect 162268 157100 171600 157128
rect 162268 157088 162274 157100
rect 171594 157088 171600 157100
rect 171652 157088 171658 157140
rect 191098 157088 191104 157140
rect 191156 157128 191162 157140
rect 246574 157128 246580 157140
rect 191156 157100 246580 157128
rect 191156 157088 191162 157100
rect 246574 157088 246580 157100
rect 246632 157088 246638 157140
rect 174354 157020 174360 157072
rect 174412 157060 174418 157072
rect 234154 157060 234160 157072
rect 174412 157032 234160 157060
rect 174412 157020 174418 157032
rect 234154 157020 234160 157032
rect 234212 157020 234218 157072
rect 123478 156952 123484 157004
rect 123536 156992 123542 157004
rect 167638 156992 167644 157004
rect 123536 156964 167644 156992
rect 123536 156952 123542 156964
rect 167638 156952 167644 156964
rect 167696 156952 167702 157004
rect 175734 156952 175740 157004
rect 175792 156992 175798 157004
rect 235442 156992 235448 157004
rect 175792 156964 235448 156992
rect 175792 156952 175798 156964
rect 235442 156952 235448 156964
rect 235500 156952 235506 157004
rect 106274 156884 106280 156936
rect 106332 156924 106338 156936
rect 170674 156924 170680 156936
rect 106332 156896 170680 156924
rect 106332 156884 106338 156896
rect 170674 156884 170680 156896
rect 170732 156884 170738 156936
rect 181070 156884 181076 156936
rect 181128 156924 181134 156936
rect 240134 156924 240140 156936
rect 181128 156896 240140 156924
rect 181128 156884 181134 156896
rect 240134 156884 240140 156896
rect 240192 156924 240198 156936
rect 240962 156924 240968 156936
rect 240192 156896 240968 156924
rect 240192 156884 240198 156896
rect 240962 156884 240968 156896
rect 241020 156884 241026 156936
rect 99374 156816 99380 156868
rect 99432 156856 99438 156868
rect 162118 156856 162124 156868
rect 99432 156828 162124 156856
rect 99432 156816 99438 156828
rect 162118 156816 162124 156828
rect 162176 156816 162182 156868
rect 189350 156816 189356 156868
rect 189408 156856 189414 156868
rect 247954 156856 247960 156868
rect 189408 156828 247960 156856
rect 189408 156816 189414 156828
rect 247954 156816 247960 156828
rect 248012 156816 248018 156868
rect 85574 156748 85580 156800
rect 85632 156788 85638 156800
rect 169018 156788 169024 156800
rect 85632 156760 169024 156788
rect 85632 156748 85638 156760
rect 169018 156748 169024 156760
rect 169076 156748 169082 156800
rect 179598 156748 179604 156800
rect 179656 156788 179662 156800
rect 200850 156788 200856 156800
rect 179656 156760 200856 156788
rect 179656 156748 179662 156760
rect 200850 156748 200856 156760
rect 200908 156748 200914 156800
rect 81434 156680 81440 156732
rect 81492 156720 81498 156732
rect 168742 156720 168748 156732
rect 81492 156692 168748 156720
rect 81492 156680 81498 156692
rect 168742 156680 168748 156692
rect 168800 156680 168806 156732
rect 178494 156680 178500 156732
rect 178552 156720 178558 156732
rect 207750 156720 207756 156732
rect 178552 156692 207756 156720
rect 178552 156680 178558 156692
rect 207750 156680 207756 156692
rect 207808 156680 207814 156732
rect 271782 156680 271788 156732
rect 271840 156720 271846 156732
rect 289078 156720 289084 156732
rect 271840 156692 289084 156720
rect 271840 156680 271846 156692
rect 289078 156680 289084 156692
rect 289136 156680 289142 156732
rect 74534 156612 74540 156664
rect 74592 156652 74598 156664
rect 168190 156652 168196 156664
rect 74592 156624 168196 156652
rect 74592 156612 74598 156624
rect 168190 156612 168196 156624
rect 168248 156612 168254 156664
rect 171134 156612 171140 156664
rect 171192 156652 171198 156664
rect 171502 156652 171508 156664
rect 171192 156624 171508 156652
rect 171192 156612 171198 156624
rect 171502 156612 171508 156624
rect 171560 156612 171566 156664
rect 178770 156612 178776 156664
rect 178828 156652 178834 156664
rect 209498 156652 209504 156664
rect 178828 156624 209504 156652
rect 178828 156612 178834 156624
rect 209498 156612 209504 156624
rect 209556 156652 209562 156664
rect 213638 156652 213644 156664
rect 209556 156624 213644 156652
rect 209556 156612 209562 156624
rect 213638 156612 213644 156624
rect 213696 156612 213702 156664
rect 288526 156652 288532 156664
rect 277366 156624 288532 156652
rect 162118 156544 162124 156596
rect 162176 156584 162182 156596
rect 169754 156584 169760 156596
rect 162176 156556 169760 156584
rect 162176 156544 162182 156556
rect 169754 156544 169760 156556
rect 169812 156544 169818 156596
rect 186038 156544 186044 156596
rect 186096 156584 186102 156596
rect 191098 156584 191104 156596
rect 186096 156556 191104 156584
rect 186096 156544 186102 156556
rect 191098 156544 191104 156556
rect 191156 156544 191162 156596
rect 207014 156584 207020 156596
rect 195946 156556 207020 156584
rect 192938 156476 192944 156528
rect 192996 156516 193002 156528
rect 195946 156516 195974 156556
rect 207014 156544 207020 156556
rect 207072 156544 207078 156596
rect 220538 156516 220544 156528
rect 192996 156488 195974 156516
rect 200684 156488 220544 156516
rect 192996 156476 193002 156488
rect 151722 156408 151728 156460
rect 151780 156448 151786 156460
rect 163498 156448 163504 156460
rect 151780 156420 163504 156448
rect 151780 156408 151786 156420
rect 163498 156408 163504 156420
rect 163556 156408 163562 156460
rect 161382 156340 161388 156392
rect 161440 156380 161446 156392
rect 174906 156380 174912 156392
rect 161440 156352 174912 156380
rect 161440 156340 161446 156352
rect 174906 156340 174912 156352
rect 174964 156340 174970 156392
rect 172882 156272 172888 156324
rect 172940 156312 172946 156324
rect 200684 156312 200712 156488
rect 220538 156476 220544 156488
rect 220596 156476 220602 156528
rect 277366 156448 277394 156624
rect 288526 156612 288532 156624
rect 288584 156652 288590 156664
rect 430574 156652 430580 156664
rect 288584 156624 430580 156652
rect 288584 156612 288590 156624
rect 430574 156612 430580 156624
rect 430632 156612 430638 156664
rect 205606 156420 277394 156448
rect 205606 156380 205634 156420
rect 172940 156284 200712 156312
rect 200776 156352 205634 156380
rect 172940 156272 172946 156284
rect 164234 156204 164240 156256
rect 164292 156244 164298 156256
rect 164970 156244 164976 156256
rect 164292 156216 164976 156244
rect 164292 156204 164298 156216
rect 164970 156204 164976 156216
rect 165028 156204 165034 156256
rect 195790 156204 195796 156256
rect 195848 156244 195854 156256
rect 200776 156244 200804 156352
rect 200850 156272 200856 156324
rect 200908 156312 200914 156324
rect 211798 156312 211804 156324
rect 200908 156284 211804 156312
rect 200908 156272 200914 156284
rect 211798 156272 211804 156284
rect 211856 156272 211862 156324
rect 195848 156216 200804 156244
rect 195848 156204 195854 156216
rect 200114 156136 200120 156188
rect 200172 156176 200178 156188
rect 200942 156176 200948 156188
rect 200172 156148 200948 156176
rect 200172 156136 200178 156148
rect 200942 156136 200948 156148
rect 201000 156136 201006 156188
rect 167178 156068 167184 156120
rect 167236 156108 167242 156120
rect 168098 156108 168104 156120
rect 167236 156080 168104 156108
rect 167236 156068 167242 156080
rect 168098 156068 168104 156080
rect 168156 156068 168162 156120
rect 160738 155932 160744 155984
rect 160796 155972 160802 155984
rect 166350 155972 166356 155984
rect 160796 155944 166356 155972
rect 160796 155932 160802 155944
rect 166350 155932 166356 155944
rect 166408 155932 166414 155984
rect 168650 155932 168656 155984
rect 168708 155972 168714 155984
rect 169110 155972 169116 155984
rect 168708 155944 169116 155972
rect 168708 155932 168714 155944
rect 169110 155932 169116 155944
rect 169168 155932 169174 155984
rect 169938 155932 169944 155984
rect 169996 155972 170002 155984
rect 170306 155972 170312 155984
rect 169996 155944 170312 155972
rect 169996 155932 170002 155944
rect 170306 155932 170312 155944
rect 170364 155932 170370 155984
rect 171226 155932 171232 155984
rect 171284 155972 171290 155984
rect 171870 155972 171876 155984
rect 171284 155944 171876 155972
rect 171284 155932 171290 155944
rect 171870 155932 171876 155944
rect 171928 155932 171934 155984
rect 177114 155932 177120 155984
rect 177172 155972 177178 155984
rect 181438 155972 181444 155984
rect 177172 155944 181444 155972
rect 177172 155932 177178 155944
rect 181438 155932 181444 155944
rect 181496 155932 181502 155984
rect 211798 155932 211804 155984
rect 211856 155972 211862 155984
rect 212258 155972 212264 155984
rect 211856 155944 212264 155972
rect 211856 155932 211862 155944
rect 212258 155932 212264 155944
rect 212316 155932 212322 155984
rect 289354 155932 289360 155984
rect 289412 155972 289418 155984
rect 518894 155972 518900 155984
rect 289412 155944 518900 155972
rect 289412 155932 289418 155944
rect 518894 155932 518900 155944
rect 518952 155932 518958 155984
rect 149698 155864 149704 155916
rect 149756 155904 149762 155916
rect 150342 155904 150348 155916
rect 149756 155876 150348 155904
rect 149756 155864 149762 155876
rect 150342 155864 150348 155876
rect 150400 155904 150406 155916
rect 165062 155904 165068 155916
rect 150400 155876 165068 155904
rect 150400 155864 150406 155876
rect 165062 155864 165068 155876
rect 165120 155864 165126 155916
rect 169294 155864 169300 155916
rect 169352 155904 169358 155916
rect 169662 155904 169668 155916
rect 169352 155876 169668 155904
rect 169352 155864 169358 155876
rect 169662 155864 169668 155876
rect 169720 155864 169726 155916
rect 175458 155864 175464 155916
rect 175516 155904 175522 155916
rect 176378 155904 176384 155916
rect 175516 155876 176384 155904
rect 175516 155864 175522 155876
rect 176378 155864 176384 155876
rect 176436 155904 176442 155916
rect 176436 155876 176654 155904
rect 176436 155864 176442 155876
rect 155770 155728 155776 155780
rect 155828 155768 155834 155780
rect 166626 155768 166632 155780
rect 155828 155740 166632 155768
rect 155828 155728 155834 155740
rect 166626 155728 166632 155740
rect 166684 155728 166690 155780
rect 161842 155660 161848 155712
rect 161900 155700 161906 155712
rect 163222 155700 163228 155712
rect 161900 155672 163228 155700
rect 161900 155660 161906 155672
rect 163222 155660 163228 155672
rect 163280 155660 163286 155712
rect 168466 155660 168472 155712
rect 168524 155700 168530 155712
rect 169202 155700 169208 155712
rect 168524 155672 169208 155700
rect 168524 155660 168530 155672
rect 169202 155660 169208 155672
rect 169260 155660 169266 155712
rect 171134 155660 171140 155712
rect 171192 155700 171198 155712
rect 175734 155700 175740 155712
rect 171192 155672 175740 155700
rect 171192 155660 171198 155672
rect 175734 155660 175740 155672
rect 175792 155660 175798 155712
rect 176626 155700 176654 155876
rect 187510 155864 187516 155916
rect 187568 155904 187574 155916
rect 210602 155904 210608 155916
rect 187568 155876 210608 155904
rect 187568 155864 187574 155876
rect 210602 155864 210608 155876
rect 210660 155864 210666 155916
rect 203058 155796 203064 155848
rect 203116 155836 203122 155848
rect 282270 155836 282276 155848
rect 203116 155808 282276 155836
rect 203116 155796 203122 155808
rect 282270 155796 282276 155808
rect 282328 155836 282334 155848
rect 282546 155836 282552 155848
rect 282328 155808 282552 155836
rect 282328 155796 282334 155808
rect 282546 155796 282552 155808
rect 282604 155796 282610 155848
rect 178034 155728 178040 155780
rect 178092 155768 178098 155780
rect 201494 155768 201500 155780
rect 178092 155740 201500 155768
rect 178092 155728 178098 155740
rect 201494 155728 201500 155740
rect 201552 155728 201558 155780
rect 207198 155728 207204 155780
rect 207256 155768 207262 155780
rect 207750 155768 207756 155780
rect 207256 155740 207756 155768
rect 207256 155728 207262 155740
rect 207750 155728 207756 155740
rect 207808 155768 207814 155780
rect 215938 155768 215944 155780
rect 207808 155740 215944 155768
rect 207808 155728 207814 155740
rect 215938 155728 215944 155740
rect 215996 155728 216002 155780
rect 235258 155700 235264 155712
rect 176626 155672 235264 155700
rect 235258 155660 235264 155672
rect 235316 155660 235322 155712
rect 164786 155592 164792 155644
rect 164844 155632 164850 155644
rect 175182 155632 175188 155644
rect 164844 155604 175188 155632
rect 164844 155592 164850 155604
rect 175182 155592 175188 155604
rect 175240 155632 175246 155644
rect 219066 155632 219072 155644
rect 175240 155604 219072 155632
rect 175240 155592 175246 155604
rect 219066 155592 219072 155604
rect 219124 155592 219130 155644
rect 173342 155524 173348 155576
rect 173400 155564 173406 155576
rect 173526 155564 173532 155576
rect 173400 155536 173532 155564
rect 173400 155524 173406 155536
rect 173526 155524 173532 155536
rect 173584 155564 173590 155576
rect 215754 155564 215760 155576
rect 173584 155536 215760 155564
rect 173584 155524 173590 155536
rect 215754 155524 215760 155536
rect 215812 155524 215818 155576
rect 176286 155456 176292 155508
rect 176344 155496 176350 155508
rect 178034 155496 178040 155508
rect 176344 155468 178040 155496
rect 176344 155456 176350 155468
rect 178034 155456 178040 155468
rect 178092 155456 178098 155508
rect 180150 155456 180156 155508
rect 180208 155496 180214 155508
rect 220630 155496 220636 155508
rect 180208 155468 220636 155496
rect 180208 155456 180214 155468
rect 220630 155456 220636 155468
rect 220688 155496 220694 155508
rect 225598 155496 225604 155508
rect 220688 155468 225604 155496
rect 220688 155456 220694 155468
rect 225598 155456 225604 155468
rect 225656 155456 225662 155508
rect 252554 155456 252560 155508
rect 252612 155496 252618 155508
rect 253198 155496 253204 155508
rect 252612 155468 253204 155496
rect 252612 155456 252618 155468
rect 253198 155456 253204 155468
rect 253256 155456 253262 155508
rect 153194 155388 153200 155440
rect 153252 155428 153258 155440
rect 174354 155428 174360 155440
rect 153252 155400 174360 155428
rect 153252 155388 153258 155400
rect 174354 155388 174360 155400
rect 174412 155388 174418 155440
rect 202598 155388 202604 155440
rect 202656 155428 202662 155440
rect 237006 155428 237012 155440
rect 202656 155400 237012 155428
rect 202656 155388 202662 155400
rect 237006 155388 237012 155400
rect 237064 155388 237070 155440
rect 144914 155320 144920 155372
rect 144972 155360 144978 155372
rect 173710 155360 173716 155372
rect 144972 155332 173716 155360
rect 144972 155320 144978 155332
rect 173710 155320 173716 155332
rect 173768 155320 173774 155372
rect 179322 155320 179328 155372
rect 179380 155360 179386 155372
rect 210326 155360 210332 155372
rect 179380 155332 210332 155360
rect 179380 155320 179386 155332
rect 210326 155320 210332 155332
rect 210384 155320 210390 155372
rect 25498 155252 25504 155304
rect 25556 155292 25562 155304
rect 164326 155292 164332 155304
rect 25556 155264 164332 155292
rect 25556 155252 25562 155264
rect 164326 155252 164332 155264
rect 164384 155252 164390 155304
rect 197998 155252 198004 155304
rect 198056 155292 198062 155304
rect 221826 155292 221832 155304
rect 198056 155264 221832 155292
rect 198056 155252 198062 155264
rect 221826 155252 221832 155264
rect 221884 155252 221890 155304
rect 6914 155184 6920 155236
rect 6972 155224 6978 155236
rect 155862 155224 155868 155236
rect 6972 155196 155868 155224
rect 6972 155184 6978 155196
rect 155862 155184 155868 155196
rect 155920 155184 155926 155236
rect 155954 155184 155960 155236
rect 156012 155224 156018 155236
rect 174538 155224 174544 155236
rect 156012 155196 174544 155224
rect 156012 155184 156018 155196
rect 174538 155184 174544 155196
rect 174596 155184 174602 155236
rect 178034 155184 178040 155236
rect 178092 155224 178098 155236
rect 216306 155224 216312 155236
rect 178092 155196 216312 155224
rect 178092 155184 178098 155196
rect 216306 155184 216312 155196
rect 216364 155184 216370 155236
rect 282270 155184 282276 155236
rect 282328 155224 282334 155236
rect 522298 155224 522304 155236
rect 282328 155196 522304 155224
rect 282328 155184 282334 155196
rect 522298 155184 522304 155196
rect 522356 155184 522362 155236
rect 190730 155116 190736 155168
rect 190788 155156 190794 155168
rect 202138 155156 202144 155168
rect 190788 155128 202144 155156
rect 190788 155116 190794 155128
rect 202138 155116 202144 155128
rect 202196 155116 202202 155168
rect 203610 155116 203616 155168
rect 203668 155156 203674 155168
rect 204070 155156 204076 155168
rect 203668 155128 204076 155156
rect 203668 155116 203674 155128
rect 204070 155116 204076 155128
rect 204128 155116 204134 155168
rect 183738 155048 183744 155100
rect 183796 155088 183802 155100
rect 271138 155088 271144 155100
rect 183796 155060 271144 155088
rect 183796 155048 183802 155060
rect 271138 155048 271144 155060
rect 271196 155048 271202 155100
rect 179874 154980 179880 155032
rect 179932 155020 179938 155032
rect 212442 155020 212448 155032
rect 179932 154992 212448 155020
rect 179932 154980 179938 154992
rect 212442 154980 212448 154992
rect 212500 154980 212506 155032
rect 182450 154912 182456 154964
rect 182508 154952 182514 154964
rect 252554 154952 252560 154964
rect 182508 154924 252560 154952
rect 182508 154912 182514 154924
rect 252554 154912 252560 154924
rect 252612 154912 252618 154964
rect 188798 154844 188804 154896
rect 188856 154884 188862 154896
rect 207106 154884 207112 154896
rect 188856 154856 207112 154884
rect 188856 154844 188862 154856
rect 207106 154844 207112 154856
rect 207164 154844 207170 154896
rect 167546 154776 167552 154828
rect 167604 154816 167610 154828
rect 168282 154816 168288 154828
rect 167604 154788 168288 154816
rect 167604 154776 167610 154788
rect 168282 154776 168288 154788
rect 168340 154776 168346 154828
rect 177666 154776 177672 154828
rect 177724 154816 177730 154828
rect 180058 154816 180064 154828
rect 177724 154788 180064 154816
rect 177724 154776 177730 154788
rect 180058 154776 180064 154788
rect 180116 154776 180122 154828
rect 212442 154572 212448 154624
rect 212500 154612 212506 154624
rect 213178 154612 213184 154624
rect 212500 154584 213184 154612
rect 212500 154572 212506 154584
rect 213178 154572 213184 154584
rect 213236 154572 213242 154624
rect 275646 154572 275652 154624
rect 275704 154612 275710 154624
rect 494054 154612 494060 154624
rect 275704 154584 494060 154612
rect 275704 154572 275710 154584
rect 494054 154572 494060 154584
rect 494112 154572 494118 154624
rect 192386 154504 192392 154556
rect 192444 154544 192450 154556
rect 207566 154544 207572 154556
rect 192444 154516 207572 154544
rect 192444 154504 192450 154516
rect 207566 154504 207572 154516
rect 207624 154504 207630 154556
rect 200850 154476 200856 154488
rect 195946 154448 200856 154476
rect 178310 154368 178316 154420
rect 178368 154408 178374 154420
rect 195946 154408 195974 154448
rect 200850 154436 200856 154448
rect 200908 154436 200914 154488
rect 205818 154436 205824 154488
rect 205876 154476 205882 154488
rect 282270 154476 282276 154488
rect 205876 154448 282276 154476
rect 205876 154436 205882 154448
rect 282270 154436 282276 154448
rect 282328 154436 282334 154488
rect 178368 154380 195974 154408
rect 178368 154368 178374 154380
rect 197446 154368 197452 154420
rect 197504 154408 197510 154420
rect 197906 154408 197912 154420
rect 197504 154380 197912 154408
rect 197504 154368 197510 154380
rect 197906 154368 197912 154380
rect 197964 154368 197970 154420
rect 202046 154368 202052 154420
rect 202104 154408 202110 154420
rect 277394 154408 277400 154420
rect 202104 154380 277400 154408
rect 202104 154368 202110 154380
rect 277394 154368 277400 154380
rect 277452 154368 277458 154420
rect 175826 154300 175832 154352
rect 175884 154340 175890 154352
rect 176562 154340 176568 154352
rect 175884 154312 176568 154340
rect 175884 154300 175890 154312
rect 176562 154300 176568 154312
rect 176620 154340 176626 154352
rect 235626 154340 235632 154352
rect 176620 154312 235632 154340
rect 176620 154300 176626 154312
rect 235626 154300 235632 154312
rect 235684 154300 235690 154352
rect 173434 154232 173440 154284
rect 173492 154272 173498 154284
rect 173710 154272 173716 154284
rect 173492 154244 173716 154272
rect 173492 154232 173498 154244
rect 173710 154232 173716 154244
rect 173768 154272 173774 154284
rect 228542 154272 228548 154284
rect 173768 154244 228548 154272
rect 173768 154232 173774 154244
rect 228542 154232 228548 154244
rect 228600 154232 228606 154284
rect 182910 154164 182916 154216
rect 182968 154204 182974 154216
rect 233142 154204 233148 154216
rect 182968 154176 233148 154204
rect 182968 154164 182974 154176
rect 233142 154164 233148 154176
rect 233200 154204 233206 154216
rect 233200 154176 238754 154204
rect 233200 154164 233206 154176
rect 182174 154096 182180 154148
rect 182232 154136 182238 154148
rect 183186 154136 183192 154148
rect 182232 154108 183192 154136
rect 182232 154096 182238 154108
rect 183186 154096 183192 154108
rect 183244 154096 183250 154148
rect 187970 154096 187976 154148
rect 188028 154136 188034 154148
rect 238202 154136 238208 154148
rect 188028 154108 238208 154136
rect 188028 154096 188034 154108
rect 238202 154096 238208 154108
rect 238260 154096 238266 154148
rect 174998 154028 175004 154080
rect 175056 154068 175062 154080
rect 217318 154068 217324 154080
rect 175056 154040 217324 154068
rect 175056 154028 175062 154040
rect 217318 154028 217324 154040
rect 217376 154028 217382 154080
rect 138014 153960 138020 154012
rect 138072 154000 138078 154012
rect 172514 154000 172520 154012
rect 138072 153972 172520 154000
rect 138072 153960 138078 153972
rect 172514 153960 172520 153972
rect 172572 153960 172578 154012
rect 185486 153960 185492 154012
rect 185544 154000 185550 154012
rect 223298 154000 223304 154012
rect 185544 153972 223304 154000
rect 185544 153960 185550 153972
rect 223298 153960 223304 153972
rect 223356 153960 223362 154012
rect 92474 153892 92480 153944
rect 92532 153932 92538 153944
rect 169570 153932 169576 153944
rect 92532 153904 169576 153932
rect 92532 153892 92538 153904
rect 169570 153892 169576 153904
rect 169628 153892 169634 153944
rect 180610 153892 180616 153944
rect 180668 153932 180674 153944
rect 214558 153932 214564 153944
rect 180668 153904 214564 153932
rect 180668 153892 180674 153904
rect 214558 153892 214564 153904
rect 214616 153892 214622 153944
rect 57974 153824 57980 153876
rect 58032 153864 58038 153876
rect 156782 153864 156788 153876
rect 58032 153836 156788 153864
rect 58032 153824 58038 153836
rect 156782 153824 156788 153836
rect 156840 153824 156846 153876
rect 178586 153824 178592 153876
rect 178644 153864 178650 153876
rect 208394 153864 208400 153876
rect 178644 153836 208400 153864
rect 178644 153824 178650 153836
rect 208394 153824 208400 153836
rect 208452 153864 208458 153876
rect 209590 153864 209596 153876
rect 208452 153836 209596 153864
rect 208452 153824 208458 153836
rect 209590 153824 209596 153836
rect 209648 153824 209654 153876
rect 238726 153864 238754 154176
rect 269114 154096 269120 154148
rect 269172 154136 269178 154148
rect 270126 154136 270132 154148
rect 269172 154108 270132 154136
rect 269172 154096 269178 154108
rect 270126 154096 270132 154108
rect 270184 154096 270190 154148
rect 250438 153864 250444 153876
rect 238726 153836 250444 153864
rect 250438 153824 250444 153836
rect 250496 153824 250502 153876
rect 282270 153824 282276 153876
rect 282328 153864 282334 153876
rect 557534 153864 557540 153876
rect 282328 153836 557540 153864
rect 282328 153824 282334 153836
rect 557534 153824 557540 153836
rect 557592 153824 557598 153876
rect 189074 153756 189080 153808
rect 189132 153796 189138 153808
rect 202874 153796 202880 153808
rect 189132 153768 202880 153796
rect 189132 153756 189138 153768
rect 202874 153756 202880 153768
rect 202932 153756 202938 153808
rect 180702 153688 180708 153740
rect 180760 153728 180766 153740
rect 220722 153728 220728 153740
rect 180760 153700 220728 153728
rect 180760 153688 180766 153700
rect 220722 153688 220728 153700
rect 220780 153728 220786 153740
rect 228358 153728 228364 153740
rect 220780 153700 228364 153728
rect 220780 153688 220786 153700
rect 228358 153688 228364 153700
rect 228416 153688 228422 153740
rect 183830 153620 183836 153672
rect 183888 153660 183894 153672
rect 276290 153660 276296 153672
rect 183888 153632 276296 153660
rect 183888 153620 183894 153632
rect 276290 153620 276296 153632
rect 276348 153620 276354 153672
rect 195606 153552 195612 153604
rect 195664 153592 195670 153604
rect 207290 153592 207296 153604
rect 195664 153564 207296 153592
rect 195664 153552 195670 153564
rect 207290 153552 207296 153564
rect 207348 153552 207354 153604
rect 184934 153416 184940 153468
rect 184992 153456 184998 153468
rect 185854 153456 185860 153468
rect 184992 153428 185860 153456
rect 184992 153416 184998 153428
rect 185854 153416 185860 153428
rect 185912 153416 185918 153468
rect 197630 153348 197636 153400
rect 197688 153388 197694 153400
rect 197998 153388 198004 153400
rect 197688 153360 198004 153388
rect 197688 153348 197694 153360
rect 197998 153348 198004 153360
rect 198056 153348 198062 153400
rect 296622 153280 296628 153332
rect 296680 153320 296686 153332
rect 507854 153320 507860 153332
rect 296680 153292 507860 153320
rect 296680 153280 296686 153292
rect 507854 153280 507860 153292
rect 507912 153280 507918 153332
rect 205726 153212 205732 153264
rect 205784 153252 205790 153264
rect 206002 153252 206008 153264
rect 205784 153224 206008 153252
rect 205784 153212 205790 153224
rect 206002 153212 206008 153224
rect 206060 153212 206066 153264
rect 206186 153212 206192 153264
rect 206244 153252 206250 153264
rect 206646 153252 206652 153264
rect 206244 153224 206652 153252
rect 206244 153212 206250 153224
rect 206646 153212 206652 153224
rect 206704 153212 206710 153264
rect 209700 153224 209912 153252
rect 172606 153144 172612 153196
rect 172664 153184 172670 153196
rect 176562 153184 176568 153196
rect 172664 153156 176568 153184
rect 172664 153144 172670 153156
rect 176562 153144 176568 153156
rect 176620 153144 176626 153196
rect 202230 153144 202236 153196
rect 202288 153184 202294 153196
rect 202598 153184 202604 153196
rect 202288 153156 202604 153184
rect 202288 153144 202294 153156
rect 202598 153144 202604 153156
rect 202656 153144 202662 153196
rect 205634 153144 205640 153196
rect 205692 153184 205698 153196
rect 206370 153184 206376 153196
rect 205692 153156 206376 153184
rect 205692 153144 205698 153156
rect 206370 153144 206376 153156
rect 206428 153144 206434 153196
rect 175458 153076 175464 153128
rect 175516 153116 175522 153128
rect 176470 153116 176476 153128
rect 175516 153088 176476 153116
rect 175516 153076 175522 153088
rect 176470 153076 176476 153088
rect 176528 153076 176534 153128
rect 189258 153076 189264 153128
rect 189316 153116 189322 153128
rect 189626 153116 189632 153128
rect 189316 153088 189632 153116
rect 189316 153076 189322 153088
rect 189626 153076 189632 153088
rect 189684 153076 189690 153128
rect 205266 153076 205272 153128
rect 205324 153116 205330 153128
rect 209700 153116 209728 153224
rect 209884 153184 209912 153224
rect 270126 153212 270132 153264
rect 270184 153252 270190 153264
rect 483014 153252 483020 153264
rect 270184 153224 483020 153252
rect 270184 153212 270190 153224
rect 483014 153212 483020 153224
rect 483072 153212 483078 153264
rect 209884 153156 215294 153184
rect 205324 153088 209728 153116
rect 215266 153116 215294 153156
rect 217318 153144 217324 153196
rect 217376 153184 217382 153196
rect 217778 153184 217784 153196
rect 217376 153156 217784 153184
rect 217376 153144 217382 153156
rect 217778 153144 217784 153156
rect 217836 153144 217842 153196
rect 280430 153144 280436 153196
rect 280488 153184 280494 153196
rect 579890 153184 579896 153196
rect 280488 153156 579896 153184
rect 280488 153144 280494 153156
rect 579890 153144 579896 153156
rect 579948 153144 579954 153196
rect 287974 153116 287980 153128
rect 215266 153088 287980 153116
rect 205324 153076 205330 153088
rect 287974 153076 287980 153088
rect 288032 153116 288038 153128
rect 288342 153116 288348 153128
rect 288032 153088 288348 153116
rect 288032 153076 288038 153088
rect 288342 153076 288348 153088
rect 288400 153076 288406 153128
rect 188890 153008 188896 153060
rect 188948 153048 188954 153060
rect 209682 153048 209688 153060
rect 188948 153020 209688 153048
rect 188948 153008 188954 153020
rect 209682 153008 209688 153020
rect 209740 153008 209746 153060
rect 209774 153008 209780 153060
rect 209832 153048 209838 153060
rect 218974 153048 218980 153060
rect 209832 153020 218980 153048
rect 209832 153008 209838 153020
rect 218974 153008 218980 153020
rect 219032 153008 219038 153060
rect 175274 152940 175280 152992
rect 175332 152980 175338 152992
rect 176010 152980 176016 152992
rect 175332 152952 176016 152980
rect 175332 152940 175338 152952
rect 176010 152940 176016 152952
rect 176068 152940 176074 152992
rect 187694 152940 187700 152992
rect 187752 152980 187758 152992
rect 247770 152980 247776 152992
rect 187752 152952 247776 152980
rect 187752 152940 187758 152952
rect 247770 152940 247776 152952
rect 247828 152940 247834 152992
rect 183278 152872 183284 152924
rect 183336 152912 183342 152924
rect 241330 152912 241336 152924
rect 183336 152884 241336 152912
rect 183336 152872 183342 152884
rect 241330 152872 241336 152884
rect 241388 152912 241394 152924
rect 246298 152912 246304 152924
rect 241388 152884 246304 152912
rect 241388 152872 241394 152884
rect 246298 152872 246304 152884
rect 246356 152872 246362 152924
rect 176746 152804 176752 152856
rect 176804 152844 176810 152856
rect 179322 152844 179328 152856
rect 176804 152816 179328 152844
rect 176804 152804 176810 152816
rect 179322 152804 179328 152816
rect 179380 152804 179386 152856
rect 181806 152804 181812 152856
rect 181864 152844 181870 152856
rect 235350 152844 235356 152856
rect 181864 152816 235356 152844
rect 181864 152804 181870 152816
rect 235350 152804 235356 152816
rect 235408 152804 235414 152856
rect 195974 152736 195980 152788
rect 196032 152776 196038 152788
rect 196986 152776 196992 152788
rect 196032 152748 196992 152776
rect 196032 152736 196038 152748
rect 196986 152736 196992 152748
rect 197044 152736 197050 152788
rect 197170 152736 197176 152788
rect 197228 152776 197234 152788
rect 239582 152776 239588 152788
rect 197228 152748 239588 152776
rect 197228 152736 197234 152748
rect 239582 152736 239588 152748
rect 239640 152736 239646 152788
rect 174630 152668 174636 152720
rect 174688 152708 174694 152720
rect 215110 152708 215116 152720
rect 174688 152680 195100 152708
rect 174688 152668 174694 152680
rect 133874 152600 133880 152652
rect 133932 152640 133938 152652
rect 173710 152640 173716 152652
rect 133932 152612 173716 152640
rect 133932 152600 133938 152612
rect 173710 152600 173716 152612
rect 173768 152600 173774 152652
rect 186314 152600 186320 152652
rect 186372 152640 186378 152652
rect 187326 152640 187332 152652
rect 186372 152612 187332 152640
rect 186372 152600 186378 152612
rect 187326 152600 187332 152612
rect 187384 152600 187390 152652
rect 190546 152600 190552 152652
rect 190604 152640 190610 152652
rect 195072 152640 195100 152680
rect 195256 152680 215116 152708
rect 195256 152640 195284 152680
rect 215110 152668 215116 152680
rect 215168 152668 215174 152720
rect 190604 152612 195008 152640
rect 195072 152612 195284 152640
rect 190604 152600 190610 152612
rect 104894 152532 104900 152584
rect 104952 152572 104958 152584
rect 170858 152572 170864 152584
rect 104952 152544 170864 152572
rect 104952 152532 104958 152544
rect 170858 152532 170864 152544
rect 170916 152532 170922 152584
rect 173866 152544 178080 152572
rect 46934 152464 46940 152516
rect 46992 152504 46998 152516
rect 155586 152504 155592 152516
rect 46992 152476 155592 152504
rect 46992 152464 46998 152476
rect 155586 152464 155592 152476
rect 155644 152464 155650 152516
rect 165798 152464 165804 152516
rect 165856 152504 165862 152516
rect 166442 152504 166448 152516
rect 165856 152476 166448 152504
rect 165856 152464 165862 152476
rect 166442 152464 166448 152476
rect 166500 152464 166506 152516
rect 163222 152396 163228 152448
rect 163280 152436 163286 152448
rect 163774 152436 163780 152448
rect 163280 152408 163780 152436
rect 163280 152396 163286 152408
rect 163774 152396 163780 152408
rect 163832 152396 163838 152448
rect 173866 152380 173894 152544
rect 176654 152464 176660 152516
rect 176712 152504 176718 152516
rect 177022 152504 177028 152516
rect 176712 152476 177028 152504
rect 176712 152464 176718 152476
rect 177022 152464 177028 152476
rect 177080 152464 177086 152516
rect 177298 152464 177304 152516
rect 177356 152504 177362 152516
rect 177942 152504 177948 152516
rect 177356 152476 177948 152504
rect 177356 152464 177362 152476
rect 177942 152464 177948 152476
rect 178000 152464 178006 152516
rect 178052 152504 178080 152544
rect 179506 152532 179512 152584
rect 179564 152572 179570 152584
rect 180426 152572 180432 152584
rect 179564 152544 180432 152572
rect 179564 152532 179570 152544
rect 180426 152532 180432 152544
rect 180484 152532 180490 152584
rect 180978 152532 180984 152584
rect 181036 152572 181042 152584
rect 181036 152544 186314 152572
rect 181036 152532 181042 152544
rect 178052 152476 180196 152504
rect 176930 152396 176936 152448
rect 176988 152436 176994 152448
rect 177758 152436 177764 152448
rect 176988 152408 177764 152436
rect 176988 152396 176994 152408
rect 177758 152396 177764 152408
rect 177816 152396 177822 152448
rect 173250 152328 173256 152380
rect 173308 152368 173314 152380
rect 173802 152368 173808 152380
rect 173308 152340 173808 152368
rect 173308 152328 173314 152340
rect 173802 152328 173808 152340
rect 173860 152340 173894 152380
rect 180168 152368 180196 152476
rect 180886 152464 180892 152516
rect 180944 152504 180950 152516
rect 181990 152504 181996 152516
rect 180944 152476 181996 152504
rect 180944 152464 180950 152476
rect 181990 152464 181996 152476
rect 182048 152464 182054 152516
rect 182174 152464 182180 152516
rect 182232 152504 182238 152516
rect 182726 152504 182732 152516
rect 182232 152476 182732 152504
rect 182232 152464 182238 152476
rect 182726 152464 182732 152476
rect 182784 152464 182790 152516
rect 183738 152464 183744 152516
rect 183796 152504 183802 152516
rect 184566 152504 184572 152516
rect 183796 152476 184572 152504
rect 183796 152464 183802 152476
rect 184566 152464 184572 152476
rect 184624 152464 184630 152516
rect 186286 152504 186314 152544
rect 186498 152532 186504 152584
rect 186556 152572 186562 152584
rect 186958 152572 186964 152584
rect 186556 152544 186964 152572
rect 186556 152532 186562 152544
rect 186958 152532 186964 152544
rect 187016 152532 187022 152584
rect 187694 152532 187700 152584
rect 187752 152572 187758 152584
rect 188706 152572 188712 152584
rect 187752 152544 188712 152572
rect 187752 152532 187758 152544
rect 188706 152532 188712 152544
rect 188764 152532 188770 152584
rect 189074 152532 189080 152584
rect 189132 152572 189138 152584
rect 190362 152572 190368 152584
rect 189132 152544 190368 152572
rect 189132 152532 189138 152544
rect 190362 152532 190368 152544
rect 190420 152532 190426 152584
rect 194594 152532 194600 152584
rect 194652 152572 194658 152584
rect 194870 152572 194876 152584
rect 194652 152544 194876 152572
rect 194652 152532 194658 152544
rect 194870 152532 194876 152544
rect 194928 152532 194934 152584
rect 194980 152572 195008 152612
rect 207842 152600 207848 152652
rect 207900 152640 207906 152652
rect 307110 152640 307116 152652
rect 207900 152612 307116 152640
rect 207900 152600 207906 152612
rect 307110 152600 307116 152612
rect 307168 152600 307174 152652
rect 228726 152572 228732 152584
rect 194980 152544 228732 152572
rect 228726 152532 228732 152544
rect 228784 152532 228790 152584
rect 511994 152572 512000 152584
rect 287026 152544 512000 152572
rect 217318 152504 217324 152516
rect 186286 152476 217324 152504
rect 217318 152464 217324 152476
rect 217376 152464 217382 152516
rect 181162 152396 181168 152448
rect 181220 152436 181226 152448
rect 181898 152436 181904 152448
rect 181220 152408 181904 152436
rect 181220 152396 181226 152408
rect 181898 152396 181904 152408
rect 181956 152396 181962 152448
rect 183646 152396 183652 152448
rect 183704 152436 183710 152448
rect 184842 152436 184848 152448
rect 183704 152408 184848 152436
rect 183704 152396 183710 152408
rect 184842 152396 184848 152408
rect 184900 152396 184906 152448
rect 184934 152396 184940 152448
rect 184992 152436 184998 152448
rect 186222 152436 186228 152448
rect 184992 152408 186228 152436
rect 184992 152396 184998 152408
rect 186222 152396 186228 152408
rect 186280 152396 186286 152448
rect 186590 152396 186596 152448
rect 186648 152436 186654 152448
rect 187050 152436 187056 152448
rect 186648 152408 187056 152436
rect 186648 152396 186654 152408
rect 187050 152396 187056 152408
rect 187108 152396 187114 152448
rect 187786 152396 187792 152448
rect 187844 152436 187850 152448
rect 188430 152436 188436 152448
rect 187844 152408 188436 152436
rect 187844 152396 187850 152408
rect 188430 152396 188436 152408
rect 188488 152396 188494 152448
rect 189166 152396 189172 152448
rect 189224 152436 189230 152448
rect 189810 152436 189816 152448
rect 189224 152408 189816 152436
rect 189224 152396 189230 152408
rect 189810 152396 189816 152408
rect 189868 152396 189874 152448
rect 190638 152396 190644 152448
rect 190696 152436 190702 152448
rect 190914 152436 190920 152448
rect 190696 152408 190920 152436
rect 190696 152396 190702 152408
rect 190914 152396 190920 152408
rect 190972 152396 190978 152448
rect 191926 152396 191932 152448
rect 191984 152436 191990 152448
rect 192846 152436 192852 152448
rect 191984 152408 192852 152436
rect 191984 152396 191990 152408
rect 192846 152396 192852 152408
rect 192904 152396 192910 152448
rect 196158 152396 196164 152448
rect 196216 152436 196222 152448
rect 196434 152436 196440 152448
rect 196216 152408 196440 152436
rect 196216 152396 196222 152408
rect 196434 152396 196440 152408
rect 196492 152396 196498 152448
rect 197446 152396 197452 152448
rect 197504 152436 197510 152448
rect 197814 152436 197820 152448
rect 197504 152408 197820 152436
rect 197504 152396 197510 152408
rect 197814 152396 197820 152408
rect 197872 152396 197878 152448
rect 198734 152396 198740 152448
rect 198792 152436 198798 152448
rect 199378 152436 199384 152448
rect 198792 152408 199384 152436
rect 198792 152396 198798 152408
rect 199378 152396 199384 152408
rect 199436 152396 199442 152448
rect 200114 152396 200120 152448
rect 200172 152436 200178 152448
rect 200574 152436 200580 152448
rect 200172 152408 200580 152436
rect 200172 152396 200178 152408
rect 200574 152396 200580 152408
rect 200632 152396 200638 152448
rect 201678 152396 201684 152448
rect 201736 152436 201742 152448
rect 202506 152436 202512 152448
rect 201736 152408 202512 152436
rect 201736 152396 201742 152408
rect 202506 152396 202512 152408
rect 202564 152396 202570 152448
rect 202598 152396 202604 152448
rect 202656 152436 202662 152448
rect 284386 152436 284392 152448
rect 202656 152408 284392 152436
rect 202656 152396 202662 152408
rect 284386 152396 284392 152408
rect 284444 152436 284450 152448
rect 287026 152436 287054 152544
rect 511994 152532 512000 152544
rect 512052 152532 512058 152584
rect 288342 152464 288348 152516
rect 288400 152504 288406 152516
rect 550634 152504 550640 152516
rect 288400 152476 550640 152504
rect 288400 152464 288406 152476
rect 550634 152464 550640 152476
rect 550692 152464 550698 152516
rect 284444 152408 287054 152436
rect 284444 152396 284450 152408
rect 234062 152368 234068 152380
rect 180168 152340 234068 152368
rect 173860 152328 173866 152340
rect 234062 152328 234068 152340
rect 234120 152328 234126 152380
rect 179506 152260 179512 152312
rect 179564 152300 179570 152312
rect 179966 152300 179972 152312
rect 179564 152272 179972 152300
rect 179564 152260 179570 152272
rect 179966 152260 179972 152272
rect 180024 152260 180030 152312
rect 180150 152260 180156 152312
rect 180208 152300 180214 152312
rect 180208 152272 205864 152300
rect 180208 152260 180214 152272
rect 165614 152192 165620 152244
rect 165672 152232 165678 152244
rect 166534 152232 166540 152244
rect 165672 152204 166540 152232
rect 165672 152192 165678 152204
rect 166534 152192 166540 152204
rect 166592 152192 166598 152244
rect 178678 152192 178684 152244
rect 178736 152232 178742 152244
rect 178736 152204 195974 152232
rect 178736 152192 178742 152204
rect 179414 152124 179420 152176
rect 179472 152164 179478 152176
rect 179690 152164 179696 152176
rect 179472 152136 179696 152164
rect 179472 152124 179478 152136
rect 179690 152124 179696 152136
rect 179748 152124 179754 152176
rect 186498 152124 186504 152176
rect 186556 152164 186562 152176
rect 187602 152164 187608 152176
rect 186556 152136 187608 152164
rect 186556 152124 186562 152136
rect 187602 152124 187608 152136
rect 187660 152124 187666 152176
rect 192202 152124 192208 152176
rect 192260 152164 192266 152176
rect 193122 152164 193128 152176
rect 192260 152136 193128 152164
rect 192260 152124 192266 152136
rect 193122 152124 193128 152136
rect 193180 152124 193186 152176
rect 193490 152124 193496 152176
rect 193548 152164 193554 152176
rect 194042 152164 194048 152176
rect 193548 152136 194048 152164
rect 193548 152124 193554 152136
rect 194042 152124 194048 152136
rect 194100 152124 194106 152176
rect 177758 152056 177764 152108
rect 177816 152096 177822 152108
rect 180150 152096 180156 152108
rect 177816 152068 180156 152096
rect 177816 152056 177822 152068
rect 180150 152056 180156 152068
rect 180208 152056 180214 152108
rect 193214 152056 193220 152108
rect 193272 152096 193278 152108
rect 193858 152096 193864 152108
rect 193272 152068 193864 152096
rect 193272 152056 193278 152068
rect 193858 152056 193864 152068
rect 193916 152056 193922 152108
rect 195946 152096 195974 152204
rect 197630 152192 197636 152244
rect 197688 152232 197694 152244
rect 198642 152232 198648 152244
rect 197688 152204 198648 152232
rect 197688 152192 197694 152204
rect 198642 152192 198648 152204
rect 198700 152192 198706 152244
rect 201770 152192 201776 152244
rect 201828 152232 201834 152244
rect 202782 152232 202788 152244
rect 201828 152204 202788 152232
rect 201828 152192 201834 152204
rect 202782 152192 202788 152204
rect 202840 152192 202846 152244
rect 205836 152232 205864 152272
rect 205910 152260 205916 152312
rect 205968 152300 205974 152312
rect 206186 152300 206192 152312
rect 205968 152272 206192 152300
rect 205968 152260 205974 152272
rect 206186 152260 206192 152272
rect 206244 152260 206250 152312
rect 209866 152260 209872 152312
rect 209924 152300 209930 152312
rect 210878 152300 210884 152312
rect 209924 152272 210884 152300
rect 209924 152260 209930 152272
rect 210878 152260 210884 152272
rect 210936 152260 210942 152312
rect 211982 152232 211988 152244
rect 205836 152204 211988 152232
rect 211982 152192 211988 152204
rect 212040 152192 212046 152244
rect 209866 152096 209872 152108
rect 195946 152068 209872 152096
rect 209866 152056 209872 152068
rect 209924 152056 209930 152108
rect 193306 151988 193312 152040
rect 193364 152028 193370 152040
rect 194226 152028 194232 152040
rect 193364 152000 194232 152028
rect 193364 151988 193370 152000
rect 194226 151988 194232 152000
rect 194284 151988 194290 152040
rect 205634 151988 205640 152040
rect 205692 152028 205698 152040
rect 206922 152028 206928 152040
rect 205692 152000 206928 152028
rect 205692 151988 205698 152000
rect 206922 151988 206928 152000
rect 206980 151988 206986 152040
rect 194686 151784 194692 151836
rect 194744 151824 194750 151836
rect 195054 151824 195060 151836
rect 194744 151796 195060 151824
rect 194744 151784 194750 151796
rect 195054 151784 195060 151796
rect 195112 151784 195118 151836
rect 159726 151716 159732 151768
rect 159784 151756 159790 151768
rect 161474 151756 161480 151768
rect 159784 151728 161480 151756
rect 159784 151716 159790 151728
rect 161474 151716 161480 151728
rect 161532 151716 161538 151768
rect 181254 151716 181260 151768
rect 181312 151756 181318 151768
rect 214374 151756 214380 151768
rect 181312 151728 214380 151756
rect 181312 151716 181318 151728
rect 214374 151716 214380 151728
rect 214432 151756 214438 151768
rect 215202 151756 215208 151768
rect 214432 151728 215208 151756
rect 214432 151716 214438 151728
rect 215202 151716 215208 151728
rect 215260 151716 215266 151768
rect 186682 151648 186688 151700
rect 186740 151688 186746 151700
rect 213546 151688 213552 151700
rect 186740 151660 213552 151688
rect 186740 151648 186746 151660
rect 213546 151648 213552 151660
rect 213604 151648 213610 151700
rect 182634 151580 182640 151632
rect 182692 151620 182698 151632
rect 242710 151620 242716 151632
rect 182692 151592 242716 151620
rect 182692 151580 182698 151592
rect 242710 151580 242716 151592
rect 242768 151580 242774 151632
rect 185670 151512 185676 151564
rect 185728 151552 185734 151564
rect 245378 151552 245384 151564
rect 185728 151524 245384 151552
rect 185728 151512 185734 151524
rect 245378 151512 245384 151524
rect 245436 151512 245442 151564
rect 181622 151444 181628 151496
rect 181680 151484 181686 151496
rect 240778 151484 240784 151496
rect 181680 151456 240784 151484
rect 181680 151444 181686 151456
rect 240778 151444 240784 151456
rect 240836 151444 240842 151496
rect 183554 151376 183560 151428
rect 183612 151416 183618 151428
rect 243538 151416 243544 151428
rect 183612 151388 243544 151416
rect 183612 151376 183618 151388
rect 243538 151376 243544 151388
rect 243596 151376 243602 151428
rect 189902 151308 189908 151360
rect 189960 151348 189966 151360
rect 247862 151348 247868 151360
rect 189960 151320 247868 151348
rect 189960 151308 189966 151320
rect 247862 151308 247868 151320
rect 247920 151308 247926 151360
rect 188522 151240 188528 151292
rect 188580 151280 188586 151292
rect 246482 151280 246488 151292
rect 188580 151252 246488 151280
rect 188580 151240 188586 151252
rect 246482 151240 246488 151252
rect 246540 151240 246546 151292
rect 180794 151172 180800 151224
rect 180852 151212 180858 151224
rect 235994 151212 236000 151224
rect 180852 151184 236000 151212
rect 180852 151172 180858 151184
rect 235994 151172 236000 151184
rect 236052 151172 236058 151224
rect 151078 151104 151084 151156
rect 151136 151144 151142 151156
rect 174078 151144 174084 151156
rect 151136 151116 174084 151144
rect 151136 151104 151142 151116
rect 174078 151104 174084 151116
rect 174136 151104 174142 151156
rect 195422 151104 195428 151156
rect 195480 151144 195486 151156
rect 241514 151144 241520 151156
rect 195480 151116 241520 151144
rect 195480 151104 195486 151116
rect 241514 151104 241520 151116
rect 241572 151104 241578 151156
rect 245378 151104 245384 151156
rect 245436 151144 245442 151156
rect 295978 151144 295984 151156
rect 245436 151116 295984 151144
rect 245436 151104 245442 151116
rect 295978 151104 295984 151116
rect 296036 151104 296042 151156
rect 142154 151036 142160 151088
rect 142212 151076 142218 151088
rect 172698 151076 172704 151088
rect 142212 151048 172704 151076
rect 142212 151036 142218 151048
rect 172698 151036 172704 151048
rect 172756 151036 172762 151088
rect 198182 151036 198188 151088
rect 198240 151076 198246 151088
rect 233234 151076 233240 151088
rect 198240 151048 233240 151076
rect 198240 151036 198246 151048
rect 233234 151036 233240 151048
rect 233292 151036 233298 151088
rect 279694 151036 279700 151088
rect 279752 151076 279758 151088
rect 381630 151076 381636 151088
rect 279752 151048 381636 151076
rect 279752 151036 279758 151048
rect 381630 151036 381636 151048
rect 381688 151036 381694 151088
rect 201218 150968 201224 151020
rect 201276 151008 201282 151020
rect 229094 151008 229100 151020
rect 201276 150980 229100 151008
rect 201276 150968 201282 150980
rect 229094 150968 229100 150980
rect 229152 151008 229158 151020
rect 229830 151008 229836 151020
rect 229152 150980 229836 151008
rect 229152 150968 229158 150980
rect 229830 150968 229836 150980
rect 229888 150968 229894 151020
rect 183186 150900 183192 150952
rect 183244 150940 183250 150952
rect 251266 150940 251272 150952
rect 183244 150912 251272 150940
rect 183244 150900 183250 150912
rect 251266 150900 251272 150912
rect 251324 150900 251330 150952
rect 192294 150832 192300 150884
rect 192352 150872 192358 150884
rect 279694 150872 279700 150884
rect 192352 150844 279700 150872
rect 192352 150832 192358 150844
rect 279694 150832 279700 150844
rect 279752 150832 279758 150884
rect 235994 150492 236000 150544
rect 236052 150532 236058 150544
rect 236914 150532 236920 150544
rect 236052 150504 236920 150532
rect 236052 150492 236058 150504
rect 236914 150492 236920 150504
rect 236972 150492 236978 150544
rect 214374 150424 214380 150476
rect 214432 150464 214438 150476
rect 215938 150464 215944 150476
rect 214432 150436 215944 150464
rect 214432 150424 214438 150436
rect 215938 150424 215944 150436
rect 215996 150424 216002 150476
rect 233234 150424 233240 150476
rect 233292 150464 233298 150476
rect 233970 150464 233976 150476
rect 233292 150436 233976 150464
rect 233292 150424 233298 150436
rect 233970 150424 233976 150436
rect 234028 150424 234034 150476
rect 241514 150424 241520 150476
rect 241572 150464 241578 150476
rect 242158 150464 242164 150476
rect 241572 150436 242164 150464
rect 241572 150424 241578 150436
rect 242158 150424 242164 150436
rect 242216 150424 242222 150476
rect 242710 150424 242716 150476
rect 242768 150464 242774 150476
rect 243630 150464 243636 150476
rect 242768 150436 243636 150464
rect 242768 150424 242774 150436
rect 243630 150424 243636 150436
rect 243688 150424 243694 150476
rect 251266 150424 251272 150476
rect 251324 150464 251330 150476
rect 251818 150464 251824 150476
rect 251324 150436 251824 150464
rect 251324 150424 251330 150436
rect 251818 150424 251824 150436
rect 251876 150424 251882 150476
rect 197354 150356 197360 150408
rect 197412 150396 197418 150408
rect 292206 150396 292212 150408
rect 197412 150368 292212 150396
rect 197412 150356 197418 150368
rect 292206 150356 292212 150368
rect 292264 150356 292270 150408
rect 201494 150288 201500 150340
rect 201552 150328 201558 150340
rect 214650 150328 214656 150340
rect 201552 150300 214656 150328
rect 201552 150288 201558 150300
rect 214650 150288 214656 150300
rect 214708 150288 214714 150340
rect 184014 150220 184020 150272
rect 184072 150260 184078 150272
rect 274450 150260 274456 150272
rect 184072 150232 274456 150260
rect 184072 150220 184078 150232
rect 274450 150220 274456 150232
rect 274508 150220 274514 150272
rect 188062 150152 188068 150204
rect 188120 150192 188126 150204
rect 275186 150192 275192 150204
rect 188120 150164 275192 150192
rect 188120 150152 188126 150164
rect 275186 150152 275192 150164
rect 275244 150152 275250 150204
rect 195330 150084 195336 150136
rect 195388 150124 195394 150136
rect 260834 150124 260840 150136
rect 195388 150096 260840 150124
rect 195388 150084 195394 150096
rect 260834 150084 260840 150096
rect 260892 150084 260898 150136
rect 274634 150084 274640 150136
rect 274692 150124 274698 150136
rect 274910 150124 274916 150136
rect 274692 150096 274916 150124
rect 274692 150084 274698 150096
rect 274910 150084 274916 150096
rect 274968 150084 274974 150136
rect 190178 150016 190184 150068
rect 190236 150056 190242 150068
rect 244918 150056 244924 150068
rect 190236 150028 244924 150056
rect 190236 150016 190242 150028
rect 244918 150016 244924 150028
rect 244976 150016 244982 150068
rect 181530 149948 181536 150000
rect 181588 149988 181594 150000
rect 219434 149988 219440 150000
rect 181588 149960 219440 149988
rect 181588 149948 181594 149960
rect 219434 149948 219440 149960
rect 219492 149988 219498 150000
rect 220722 149988 220728 150000
rect 219492 149960 220728 149988
rect 219492 149948 219498 149960
rect 220722 149948 220728 149960
rect 220780 149948 220786 150000
rect 200850 149880 200856 149932
rect 200908 149920 200914 149932
rect 238386 149920 238392 149932
rect 200908 149892 238392 149920
rect 200908 149880 200914 149892
rect 238386 149880 238392 149892
rect 238444 149880 238450 149932
rect 178862 149812 178868 149864
rect 178920 149852 178926 149864
rect 211062 149852 211068 149864
rect 178920 149824 211068 149852
rect 178920 149812 178926 149824
rect 211062 149812 211068 149824
rect 211120 149812 211126 149864
rect 191834 149744 191840 149796
rect 191892 149784 191898 149796
rect 223206 149784 223212 149796
rect 191892 149756 223212 149784
rect 191892 149744 191898 149756
rect 223206 149744 223212 149756
rect 223264 149744 223270 149796
rect 275186 149744 275192 149796
rect 275244 149784 275250 149796
rect 327074 149784 327080 149796
rect 275244 149756 327080 149784
rect 275244 149744 275250 149756
rect 327074 149744 327080 149756
rect 327132 149744 327138 149796
rect 71774 149676 71780 149728
rect 71832 149716 71838 149728
rect 156874 149716 156880 149728
rect 71832 149688 156880 149716
rect 71832 149676 71838 149688
rect 156874 149676 156880 149688
rect 156932 149676 156938 149728
rect 176562 149676 176568 149728
rect 176620 149716 176626 149728
rect 182082 149716 182088 149728
rect 176620 149688 182088 149716
rect 176620 149676 176626 149688
rect 182082 149676 182088 149688
rect 182140 149716 182146 149728
rect 217502 149716 217508 149728
rect 182140 149688 217508 149716
rect 182140 149676 182146 149688
rect 217502 149676 217508 149688
rect 217560 149676 217566 149728
rect 220722 149676 220728 149728
rect 220780 149716 220786 149728
rect 232498 149716 232504 149728
rect 220780 149688 232504 149716
rect 220780 149676 220786 149688
rect 232498 149676 232504 149688
rect 232556 149676 232562 149728
rect 292206 149676 292212 149728
rect 292264 149716 292270 149728
rect 451274 149716 451280 149728
rect 292264 149688 451280 149716
rect 292264 149676 292270 149688
rect 451274 149676 451280 149688
rect 451332 149676 451338 149728
rect 187234 149608 187240 149660
rect 187292 149648 187298 149660
rect 216214 149648 216220 149660
rect 187292 149620 216220 149648
rect 187292 149608 187298 149620
rect 216214 149608 216220 149620
rect 216272 149608 216278 149660
rect 185854 149540 185860 149592
rect 185912 149580 185918 149592
rect 218882 149580 218888 149592
rect 185912 149552 218888 149580
rect 185912 149540 185918 149552
rect 218882 149540 218888 149552
rect 218940 149540 218946 149592
rect 183002 149472 183008 149524
rect 183060 149512 183066 149524
rect 274634 149512 274640 149524
rect 183060 149484 274640 149512
rect 183060 149472 183066 149484
rect 274634 149472 274640 149484
rect 274692 149472 274698 149524
rect 151814 149064 151820 149116
rect 151872 149104 151878 149116
rect 174170 149104 174176 149116
rect 151872 149076 174176 149104
rect 151872 149064 151878 149076
rect 174170 149064 174176 149076
rect 174228 149064 174234 149116
rect 206002 149064 206008 149116
rect 206060 149104 206066 149116
rect 206554 149104 206560 149116
rect 206060 149076 206560 149104
rect 206060 149064 206066 149076
rect 206554 149064 206560 149076
rect 206612 149064 206618 149116
rect 274450 149064 274456 149116
rect 274508 149104 274514 149116
rect 275094 149104 275100 149116
rect 274508 149076 275100 149104
rect 274508 149064 274514 149076
rect 275094 149064 275100 149076
rect 275152 149064 275158 149116
rect 202874 148996 202880 149048
rect 202932 149036 202938 149048
rect 228818 149036 228824 149048
rect 202932 149008 228824 149036
rect 202932 148996 202938 149008
rect 228818 148996 228824 149008
rect 228876 148996 228882 149048
rect 201402 148928 201408 148980
rect 201460 148968 201466 148980
rect 270034 148968 270040 148980
rect 201460 148940 270040 148968
rect 201460 148928 201466 148940
rect 270034 148928 270040 148940
rect 270092 148968 270098 148980
rect 270310 148968 270316 148980
rect 270092 148940 270316 148968
rect 270092 148928 270098 148940
rect 270310 148928 270316 148940
rect 270368 148928 270374 148980
rect 202322 148860 202328 148912
rect 202380 148900 202386 148912
rect 269114 148900 269120 148912
rect 202380 148872 269120 148900
rect 202380 148860 202386 148872
rect 269114 148860 269120 148872
rect 269172 148860 269178 148912
rect 184382 148792 184388 148844
rect 184440 148832 184446 148844
rect 244090 148832 244096 148844
rect 184440 148804 244096 148832
rect 184440 148792 184446 148804
rect 244090 148792 244096 148804
rect 244148 148832 244154 148844
rect 244148 148804 248414 148832
rect 244148 148792 244154 148804
rect 187970 148724 187976 148776
rect 188028 148764 188034 148776
rect 248046 148764 248052 148776
rect 188028 148736 248052 148764
rect 188028 148724 188034 148736
rect 248046 148724 248052 148736
rect 248104 148724 248110 148776
rect 184658 148656 184664 148708
rect 184716 148696 184722 148708
rect 243722 148696 243728 148708
rect 184716 148668 243728 148696
rect 184716 148656 184722 148668
rect 243722 148656 243728 148668
rect 243780 148656 243786 148708
rect 248386 148696 248414 148804
rect 278038 148696 278044 148708
rect 248386 148668 278044 148696
rect 278038 148656 278044 148668
rect 278096 148656 278102 148708
rect 185578 148588 185584 148640
rect 185636 148628 185642 148640
rect 245010 148628 245016 148640
rect 185636 148600 245016 148628
rect 185636 148588 185642 148600
rect 245010 148588 245016 148600
rect 245068 148588 245074 148640
rect 151906 148520 151912 148572
rect 151964 148560 151970 148572
rect 173894 148560 173900 148572
rect 151964 148532 173900 148560
rect 151964 148520 151970 148532
rect 173894 148520 173900 148532
rect 173952 148520 173958 148572
rect 191190 148520 191196 148572
rect 191248 148560 191254 148572
rect 249242 148560 249248 148572
rect 191248 148532 249248 148560
rect 191248 148520 191254 148532
rect 249242 148520 249248 148532
rect 249300 148520 249306 148572
rect 133138 148452 133144 148504
rect 133196 148492 133202 148504
rect 171962 148492 171968 148504
rect 133196 148464 171968 148492
rect 133196 148452 133202 148464
rect 171962 148452 171968 148464
rect 172020 148452 172026 148504
rect 191282 148452 191288 148504
rect 191340 148492 191346 148504
rect 191558 148492 191564 148504
rect 191340 148464 191564 148492
rect 191340 148452 191346 148464
rect 191558 148452 191564 148464
rect 191616 148452 191622 148504
rect 194134 148452 194140 148504
rect 194192 148492 194198 148504
rect 251910 148492 251916 148504
rect 194192 148464 251916 148492
rect 194192 148452 194198 148464
rect 251910 148452 251916 148464
rect 251968 148452 251974 148504
rect 82814 148384 82820 148436
rect 82872 148424 82878 148436
rect 152826 148424 152832 148436
rect 82872 148396 152832 148424
rect 82872 148384 82878 148396
rect 152826 148384 152832 148396
rect 152884 148384 152890 148436
rect 192662 148384 192668 148436
rect 192720 148424 192726 148436
rect 249150 148424 249156 148436
rect 192720 148396 249156 148424
rect 192720 148384 192726 148396
rect 249150 148384 249156 148396
rect 249208 148384 249214 148436
rect 281534 148384 281540 148436
rect 281592 148424 281598 148436
rect 345014 148424 345020 148436
rect 281592 148396 345020 148424
rect 281592 148384 281598 148396
rect 345014 148384 345020 148396
rect 345072 148384 345078 148436
rect 15838 148316 15844 148368
rect 15896 148356 15902 148368
rect 163406 148356 163412 148368
rect 15896 148328 163412 148356
rect 15896 148316 15902 148328
rect 163406 148316 163412 148328
rect 163464 148316 163470 148368
rect 191374 148316 191380 148368
rect 191432 148356 191438 148368
rect 249426 148356 249432 148368
rect 191432 148328 249432 148356
rect 191432 148316 191438 148328
rect 249426 148316 249432 148328
rect 249484 148316 249490 148368
rect 270310 148316 270316 148368
rect 270368 148356 270374 148368
rect 500954 148356 500960 148368
rect 270368 148328 500960 148356
rect 270368 148316 270374 148328
rect 500954 148316 500960 148328
rect 501012 148316 501018 148368
rect 174170 148248 174176 148300
rect 174228 148288 174234 148300
rect 227346 148288 227352 148300
rect 174228 148260 227352 148288
rect 174228 148248 174234 148260
rect 227346 148248 227352 148260
rect 227404 148248 227410 148300
rect 194410 148180 194416 148232
rect 194468 148220 194474 148232
rect 227162 148220 227168 148232
rect 194468 148192 227168 148220
rect 194468 148180 194474 148192
rect 227162 148180 227168 148192
rect 227220 148180 227226 148232
rect 189626 148112 189632 148164
rect 189684 148152 189690 148164
rect 281534 148152 281540 148164
rect 189684 148124 281540 148152
rect 189684 148112 189690 148124
rect 281534 148112 281540 148124
rect 281592 148112 281598 148164
rect 200850 148044 200856 148096
rect 200908 148084 200914 148096
rect 201402 148084 201408 148096
rect 200908 148056 201408 148084
rect 200908 148044 200914 148056
rect 201402 148044 201408 148056
rect 201460 148044 201466 148096
rect 173894 147636 173900 147688
rect 173952 147676 173958 147688
rect 175366 147676 175372 147688
rect 173952 147648 175372 147676
rect 173952 147636 173958 147648
rect 175366 147636 175372 147648
rect 175424 147636 175430 147688
rect 176838 147568 176844 147620
rect 176896 147608 176902 147620
rect 182818 147608 182824 147620
rect 176896 147580 182824 147608
rect 176896 147568 176902 147580
rect 182818 147568 182824 147580
rect 182876 147568 182882 147620
rect 201954 147568 201960 147620
rect 202012 147608 202018 147620
rect 296622 147608 296628 147620
rect 202012 147580 296628 147608
rect 202012 147568 202018 147580
rect 296622 147568 296628 147580
rect 296680 147568 296686 147620
rect 187878 147500 187884 147552
rect 187936 147540 187942 147552
rect 276106 147540 276112 147552
rect 187936 147512 276112 147540
rect 187936 147500 187942 147512
rect 276106 147500 276112 147512
rect 276164 147540 276170 147552
rect 276382 147540 276388 147552
rect 276164 147512 276388 147540
rect 276164 147500 276170 147512
rect 276382 147500 276388 147512
rect 276440 147500 276446 147552
rect 206094 147432 206100 147484
rect 206152 147472 206158 147484
rect 284294 147472 284300 147484
rect 206152 147444 284300 147472
rect 206152 147432 206158 147444
rect 284294 147432 284300 147444
rect 284352 147432 284358 147484
rect 182358 147364 182364 147416
rect 182416 147404 182422 147416
rect 243446 147404 243452 147416
rect 182416 147376 243452 147404
rect 182416 147364 182422 147376
rect 243446 147364 243452 147376
rect 243504 147364 243510 147416
rect 249426 147364 249432 147416
rect 249484 147404 249490 147416
rect 249702 147404 249708 147416
rect 249484 147376 249708 147404
rect 249484 147364 249490 147376
rect 249702 147364 249708 147376
rect 249760 147404 249766 147416
rect 273254 147404 273260 147416
rect 249760 147376 273260 147404
rect 249760 147364 249766 147376
rect 273254 147364 273260 147376
rect 273312 147364 273318 147416
rect 193490 147296 193496 147348
rect 193548 147336 193554 147348
rect 254670 147336 254676 147348
rect 193548 147308 254676 147336
rect 193548 147296 193554 147308
rect 254670 147296 254676 147308
rect 254728 147296 254734 147348
rect 173618 147268 173624 147280
rect 161446 147240 173624 147268
rect 143534 147024 143540 147076
rect 143592 147064 143598 147076
rect 161446 147064 161474 147240
rect 173618 147228 173624 147240
rect 173676 147268 173682 147280
rect 233326 147268 233332 147280
rect 173676 147240 233332 147268
rect 173676 147228 173682 147240
rect 233326 147228 233332 147240
rect 233384 147228 233390 147280
rect 193950 147160 193956 147212
rect 194008 147200 194014 147212
rect 253750 147200 253756 147212
rect 194008 147172 253756 147200
rect 194008 147160 194014 147172
rect 253750 147160 253756 147172
rect 253808 147200 253814 147212
rect 253808 147172 258074 147200
rect 253808 147160 253814 147172
rect 193582 147092 193588 147144
rect 193640 147132 193646 147144
rect 253474 147132 253480 147144
rect 193640 147104 253480 147132
rect 193640 147092 193646 147104
rect 253474 147092 253480 147104
rect 253532 147092 253538 147144
rect 143592 147036 161474 147064
rect 143592 147024 143598 147036
rect 194870 147024 194876 147076
rect 194928 147064 194934 147076
rect 254578 147064 254584 147076
rect 194928 147036 254584 147064
rect 194928 147024 194934 147036
rect 254578 147024 254584 147036
rect 254636 147024 254642 147076
rect 68278 146956 68284 147008
rect 68336 146996 68342 147008
rect 151262 146996 151268 147008
rect 68336 146968 151268 146996
rect 68336 146956 68342 146968
rect 151262 146956 151268 146968
rect 151320 146956 151326 147008
rect 164878 146956 164884 147008
rect 164936 146996 164942 147008
rect 165246 146996 165252 147008
rect 164936 146968 165252 146996
rect 164936 146956 164942 146968
rect 165246 146956 165252 146968
rect 165304 146956 165310 147008
rect 165890 146956 165896 147008
rect 165948 146996 165954 147008
rect 166258 146996 166264 147008
rect 165948 146968 166264 146996
rect 165948 146956 165954 146968
rect 166258 146956 166264 146968
rect 166316 146996 166322 147008
rect 258046 146996 258074 147172
rect 276382 147024 276388 147076
rect 276440 147064 276446 147076
rect 316678 147064 316684 147076
rect 276440 147036 316684 147064
rect 276440 147024 276446 147036
rect 316678 147024 316684 147036
rect 316736 147024 316742 147076
rect 405734 146996 405740 147008
rect 166316 146968 171134 146996
rect 258046 146968 405740 146996
rect 166316 146956 166322 146968
rect 14458 146888 14464 146940
rect 14516 146928 14522 146940
rect 161658 146928 161664 146940
rect 14516 146900 161664 146928
rect 14516 146888 14522 146900
rect 161658 146888 161664 146900
rect 161716 146888 161722 146940
rect 171106 146928 171134 146968
rect 405734 146956 405740 146968
rect 405792 146956 405798 147008
rect 225414 146928 225420 146940
rect 171106 146900 225420 146928
rect 225414 146888 225420 146900
rect 225472 146888 225478 146940
rect 243446 146888 243452 146940
rect 243504 146928 243510 146940
rect 253290 146928 253296 146940
rect 243504 146900 253296 146928
rect 243504 146888 243510 146900
rect 253290 146888 253296 146900
rect 253348 146888 253354 146940
rect 284294 146888 284300 146940
rect 284352 146928 284358 146940
rect 285122 146928 285128 146940
rect 284352 146900 285128 146928
rect 284352 146888 284358 146900
rect 285122 146888 285128 146900
rect 285180 146928 285186 146940
rect 561674 146928 561680 146940
rect 285180 146900 561680 146928
rect 285180 146888 285186 146900
rect 561674 146888 561680 146900
rect 561732 146888 561738 146940
rect 181806 146820 181812 146872
rect 181864 146860 181870 146872
rect 239398 146860 239404 146872
rect 181864 146832 239404 146860
rect 181864 146820 181870 146832
rect 239398 146820 239404 146832
rect 239456 146820 239462 146872
rect 203702 146752 203708 146804
rect 203760 146792 203766 146804
rect 253566 146792 253572 146804
rect 203760 146764 253572 146792
rect 203760 146752 203766 146764
rect 253566 146752 253572 146764
rect 253624 146752 253630 146804
rect 202230 146684 202236 146736
rect 202288 146724 202294 146736
rect 250622 146724 250628 146736
rect 202288 146696 250628 146724
rect 202288 146684 202294 146696
rect 250622 146684 250628 146696
rect 250680 146684 250686 146736
rect 196250 146616 196256 146668
rect 196308 146656 196314 146668
rect 255958 146656 255964 146668
rect 196308 146628 255964 146656
rect 196308 146616 196314 146628
rect 255958 146616 255964 146628
rect 256016 146616 256022 146668
rect 154206 146208 154212 146260
rect 154264 146248 154270 146260
rect 154482 146248 154488 146260
rect 154264 146220 154488 146248
rect 154264 146208 154270 146220
rect 154482 146208 154488 146220
rect 154540 146248 154546 146260
rect 169294 146248 169300 146260
rect 154540 146220 169300 146248
rect 154540 146208 154546 146220
rect 169294 146208 169300 146220
rect 169352 146208 169358 146260
rect 175550 146208 175556 146260
rect 175608 146248 175614 146260
rect 176102 146248 176108 146260
rect 175608 146220 176108 146248
rect 175608 146208 175614 146220
rect 176102 146208 176108 146220
rect 176160 146208 176166 146260
rect 201678 146208 201684 146260
rect 201736 146248 201742 146260
rect 293954 146248 293960 146260
rect 201736 146220 293960 146248
rect 201736 146208 201742 146220
rect 293954 146208 293960 146220
rect 294012 146248 294018 146260
rect 294598 146248 294604 146260
rect 294012 146220 294604 146248
rect 294012 146208 294018 146220
rect 294598 146208 294604 146220
rect 294656 146208 294662 146260
rect 201770 146140 201776 146192
rect 201828 146180 201834 146192
rect 289354 146180 289360 146192
rect 201828 146152 289360 146180
rect 201828 146140 201834 146152
rect 289354 146140 289360 146152
rect 289412 146140 289418 146192
rect 190730 146072 190736 146124
rect 190788 146112 190794 146124
rect 270310 146112 270316 146124
rect 190788 146084 270316 146112
rect 190788 146072 190794 146084
rect 270310 146072 270316 146084
rect 270368 146072 270374 146124
rect 183738 146004 183744 146056
rect 183796 146044 183802 146056
rect 245470 146044 245476 146056
rect 183796 146016 245476 146044
rect 183796 146004 183802 146016
rect 245470 146004 245476 146016
rect 245528 146044 245534 146056
rect 245528 146016 258074 146044
rect 245528 146004 245534 146016
rect 189442 145936 189448 145988
rect 189500 145976 189506 145988
rect 250898 145976 250904 145988
rect 189500 145948 250904 145976
rect 189500 145936 189506 145948
rect 250898 145936 250904 145948
rect 250956 145936 250962 145988
rect 185302 145868 185308 145920
rect 185360 145908 185366 145920
rect 246666 145908 246672 145920
rect 185360 145880 246672 145908
rect 185360 145868 185366 145880
rect 246666 145868 246672 145880
rect 246724 145868 246730 145920
rect 176102 145800 176108 145852
rect 176160 145840 176166 145852
rect 236086 145840 236092 145852
rect 176160 145812 236092 145840
rect 176160 145800 176166 145812
rect 236086 145800 236092 145812
rect 236144 145800 236150 145852
rect 258046 145840 258074 146016
rect 282178 145840 282184 145852
rect 258046 145812 282184 145840
rect 282178 145800 282184 145812
rect 282236 145800 282242 145852
rect 197998 145732 198004 145784
rect 198056 145772 198062 145784
rect 257338 145772 257344 145784
rect 198056 145744 257344 145772
rect 198056 145732 198062 145744
rect 257338 145732 257344 145744
rect 257396 145732 257402 145784
rect 118694 145664 118700 145716
rect 118752 145704 118758 145716
rect 172054 145704 172060 145716
rect 118752 145676 172060 145704
rect 118752 145664 118758 145676
rect 172054 145664 172060 145676
rect 172112 145664 172118 145716
rect 198826 145664 198832 145716
rect 198884 145704 198890 145716
rect 258166 145704 258172 145716
rect 198884 145676 258172 145704
rect 198884 145664 198890 145676
rect 258166 145664 258172 145676
rect 258224 145664 258230 145716
rect 270310 145664 270316 145716
rect 270368 145704 270374 145716
rect 359458 145704 359464 145716
rect 270368 145676 359464 145704
rect 270368 145664 270374 145676
rect 359458 145664 359464 145676
rect 359516 145664 359522 145716
rect 95878 145596 95884 145648
rect 95936 145636 95942 145648
rect 154482 145636 154488 145648
rect 95936 145608 154488 145636
rect 95936 145596 95942 145608
rect 154482 145596 154488 145608
rect 154540 145596 154546 145648
rect 226978 145636 226984 145648
rect 171106 145608 226984 145636
rect 88978 145528 88984 145580
rect 89036 145568 89042 145580
rect 168650 145568 168656 145580
rect 89036 145540 168656 145568
rect 89036 145528 89042 145540
rect 168650 145528 168656 145540
rect 168708 145568 168714 145580
rect 171106 145568 171134 145608
rect 226978 145596 226984 145608
rect 227036 145596 227042 145648
rect 250898 145596 250904 145648
rect 250956 145636 250962 145648
rect 356054 145636 356060 145648
rect 250956 145608 356060 145636
rect 250956 145596 250962 145608
rect 356054 145596 356060 145608
rect 356112 145596 356118 145648
rect 168708 145540 171134 145568
rect 168708 145528 168714 145540
rect 200850 145528 200856 145580
rect 200908 145568 200914 145580
rect 258718 145568 258724 145580
rect 200908 145540 258724 145568
rect 200908 145528 200914 145540
rect 258718 145528 258724 145540
rect 258776 145528 258782 145580
rect 293954 145528 293960 145580
rect 294012 145568 294018 145580
rect 514018 145568 514024 145580
rect 294012 145540 514024 145568
rect 294012 145528 294018 145540
rect 514018 145528 514024 145540
rect 514076 145528 514082 145580
rect 179690 145460 179696 145512
rect 179748 145500 179754 145512
rect 218054 145500 218060 145512
rect 179748 145472 218060 145500
rect 179748 145460 179754 145472
rect 218054 145460 218060 145472
rect 218112 145460 218118 145512
rect 179322 145392 179328 145444
rect 179380 145432 179386 145444
rect 213270 145432 213276 145444
rect 179380 145404 213276 145432
rect 179380 145392 179386 145404
rect 213270 145392 213276 145404
rect 213328 145392 213334 145444
rect 175458 144848 175464 144900
rect 175516 144888 175522 144900
rect 176562 144888 176568 144900
rect 175516 144860 176568 144888
rect 175516 144848 175522 144860
rect 176562 144848 176568 144860
rect 176620 144848 176626 144900
rect 202874 144848 202880 144900
rect 202932 144888 202938 144900
rect 204070 144888 204076 144900
rect 202932 144860 204076 144888
rect 202932 144848 202938 144860
rect 204070 144848 204076 144860
rect 204128 144848 204134 144900
rect 218054 144848 218060 144900
rect 218112 144888 218118 144900
rect 227070 144888 227076 144900
rect 218112 144860 227076 144888
rect 218112 144848 218118 144860
rect 227070 144848 227076 144860
rect 227128 144848 227134 144900
rect 185210 144780 185216 144832
rect 185268 144820 185274 144832
rect 278222 144820 278228 144832
rect 185268 144792 278228 144820
rect 185268 144780 185274 144792
rect 278222 144780 278228 144792
rect 278280 144820 278286 144832
rect 284938 144820 284944 144832
rect 278280 144792 284944 144820
rect 278280 144780 278286 144792
rect 284938 144780 284944 144792
rect 284996 144780 285002 144832
rect 189350 144712 189356 144764
rect 189408 144752 189414 144764
rect 280246 144752 280252 144764
rect 189408 144724 280252 144752
rect 189408 144712 189414 144724
rect 280246 144712 280252 144724
rect 280304 144752 280310 144764
rect 281442 144752 281448 144764
rect 280304 144724 281448 144752
rect 280304 144712 280310 144724
rect 281442 144712 281448 144724
rect 281500 144712 281506 144764
rect 203886 144644 203892 144696
rect 203944 144684 203950 144696
rect 268930 144684 268936 144696
rect 203944 144656 268936 144684
rect 203944 144644 203950 144656
rect 268930 144644 268936 144656
rect 268988 144644 268994 144696
rect 201126 144576 201132 144628
rect 201184 144616 201190 144628
rect 259822 144616 259828 144628
rect 201184 144588 259828 144616
rect 201184 144576 201190 144588
rect 259822 144576 259828 144588
rect 259880 144576 259886 144628
rect 201218 144508 201224 144560
rect 201276 144548 201282 144560
rect 260098 144548 260104 144560
rect 201276 144520 260104 144548
rect 201276 144508 201282 144520
rect 260098 144508 260104 144520
rect 260156 144508 260162 144560
rect 176194 144440 176200 144492
rect 176252 144480 176258 144492
rect 221458 144480 221464 144492
rect 176252 144452 221464 144480
rect 176252 144440 176258 144452
rect 221458 144440 221464 144452
rect 221516 144440 221522 144492
rect 222010 144440 222016 144492
rect 222068 144480 222074 144492
rect 222194 144480 222200 144492
rect 222068 144452 222200 144480
rect 222068 144440 222074 144452
rect 222194 144440 222200 144452
rect 222252 144440 222258 144492
rect 179598 144372 179604 144424
rect 179656 144412 179662 144424
rect 222028 144412 222056 144440
rect 179656 144384 222056 144412
rect 179656 144372 179662 144384
rect 176562 144304 176568 144356
rect 176620 144344 176626 144356
rect 216030 144344 216036 144356
rect 176620 144316 216036 144344
rect 176620 144304 176626 144316
rect 216030 144304 216036 144316
rect 216088 144304 216094 144356
rect 281442 144304 281448 144356
rect 281500 144344 281506 144356
rect 319438 144344 319444 144356
rect 281500 144316 319444 144344
rect 281500 144304 281506 144316
rect 319438 144304 319444 144316
rect 319496 144304 319502 144356
rect 93854 144236 93860 144288
rect 93912 144276 93918 144288
rect 169110 144276 169116 144288
rect 93912 144248 169116 144276
rect 93912 144236 93918 144248
rect 169110 144236 169116 144248
rect 169168 144236 169174 144288
rect 200298 144236 200304 144288
rect 200356 144276 200362 144288
rect 201218 144276 201224 144288
rect 200356 144248 201224 144276
rect 200356 144236 200362 144248
rect 201218 144236 201224 144248
rect 201276 144236 201282 144288
rect 204070 144236 204076 144288
rect 204128 144276 204134 144288
rect 228634 144276 228640 144288
rect 204128 144248 228640 144276
rect 204128 144236 204134 144248
rect 228634 144236 228640 144248
rect 228692 144236 228698 144288
rect 290918 144236 290924 144288
rect 290976 144276 290982 144288
rect 436738 144276 436744 144288
rect 290976 144248 436744 144276
rect 290976 144236 290982 144248
rect 436738 144236 436744 144248
rect 436796 144236 436802 144288
rect 13078 144168 13084 144220
rect 13136 144208 13142 144220
rect 161566 144208 161572 144220
rect 13136 144180 161572 144208
rect 13136 144168 13142 144180
rect 161566 144168 161572 144180
rect 161624 144168 161630 144220
rect 202690 144168 202696 144220
rect 202748 144208 202754 144220
rect 262398 144208 262404 144220
rect 202748 144180 262404 144208
rect 202748 144168 202754 144180
rect 262398 144168 262404 144180
rect 262456 144168 262462 144220
rect 268930 144168 268936 144220
rect 268988 144208 268994 144220
rect 532694 144208 532700 144220
rect 268988 144180 532700 144208
rect 268988 144168 268994 144180
rect 532694 144168 532700 144180
rect 532752 144168 532758 144220
rect 196158 144100 196164 144152
rect 196216 144140 196222 144152
rect 290642 144140 290648 144152
rect 196216 144112 290648 144140
rect 196216 144100 196222 144112
rect 290642 144100 290648 144112
rect 290700 144140 290706 144152
rect 290918 144140 290924 144152
rect 290700 144112 290924 144140
rect 290700 144100 290706 144112
rect 290918 144100 290924 144112
rect 290976 144100 290982 144152
rect 174630 144032 174636 144084
rect 174688 144072 174694 144084
rect 176194 144072 176200 144084
rect 174688 144044 176200 144072
rect 174688 144032 174694 144044
rect 176194 144032 176200 144044
rect 176252 144032 176258 144084
rect 185118 143488 185124 143540
rect 185176 143528 185182 143540
rect 186222 143528 186228 143540
rect 185176 143500 186228 143528
rect 185176 143488 185182 143500
rect 186222 143488 186228 143500
rect 186280 143488 186286 143540
rect 186682 143488 186688 143540
rect 186740 143528 186746 143540
rect 269206 143528 269212 143540
rect 186740 143500 269212 143528
rect 186740 143488 186746 143500
rect 269206 143488 269212 143500
rect 269264 143488 269270 143540
rect 269298 143488 269304 143540
rect 269356 143528 269362 143540
rect 269758 143528 269764 143540
rect 269356 143500 269764 143528
rect 269356 143488 269362 143500
rect 269758 143488 269764 143500
rect 269816 143488 269822 143540
rect 185026 143420 185032 143472
rect 185084 143460 185090 143472
rect 269316 143460 269344 143488
rect 185084 143432 269344 143460
rect 185084 143420 185090 143432
rect 203610 143352 203616 143404
rect 203668 143392 203674 143404
rect 283098 143392 283104 143404
rect 203668 143364 283104 143392
rect 203668 143352 203674 143364
rect 283098 143352 283104 143364
rect 283156 143392 283162 143404
rect 283558 143392 283564 143404
rect 283156 143364 283564 143392
rect 283156 143352 283162 143364
rect 283558 143352 283564 143364
rect 283616 143352 283622 143404
rect 164510 143284 164516 143336
rect 164568 143324 164574 143336
rect 224310 143324 224316 143336
rect 164568 143296 224316 143324
rect 164568 143284 164574 143296
rect 224310 143284 224316 143296
rect 224368 143284 224374 143336
rect 187786 143216 187792 143268
rect 187844 143256 187850 143268
rect 243814 143256 243820 143268
rect 187844 143228 243820 143256
rect 187844 143216 187850 143228
rect 243814 143216 243820 143228
rect 243872 143216 243878 143268
rect 169754 143148 169760 143200
rect 169812 143188 169818 143200
rect 170122 143188 170128 143200
rect 169812 143160 170128 143188
rect 169812 143148 169818 143160
rect 170122 143148 170128 143160
rect 170180 143188 170186 143200
rect 222930 143188 222936 143200
rect 170180 143160 222936 143188
rect 170180 143148 170186 143160
rect 222930 143148 222936 143160
rect 222988 143148 222994 143200
rect 186222 143080 186228 143132
rect 186280 143120 186286 143132
rect 231118 143120 231124 143132
rect 186280 143092 231124 143120
rect 186280 143080 186286 143092
rect 231118 143080 231124 143092
rect 231176 143080 231182 143132
rect 143626 143012 143632 143064
rect 143684 143052 143690 143064
rect 173342 143052 173348 143064
rect 143684 143024 173348 143052
rect 143684 143012 143690 143024
rect 173342 143012 173348 143024
rect 173400 143012 173406 143064
rect 182266 143012 182272 143064
rect 182324 143052 182330 143064
rect 182324 143024 219434 143052
rect 182324 143012 182330 143024
rect 107654 142944 107660 142996
rect 107712 142984 107718 142996
rect 169754 142984 169760 142996
rect 107712 142956 169760 142984
rect 107712 142944 107718 142956
rect 169754 142944 169760 142956
rect 169812 142944 169818 142996
rect 49694 142876 49700 142928
rect 49752 142916 49758 142928
rect 165706 142916 165712 142928
rect 49752 142888 165712 142916
rect 49752 142876 49758 142888
rect 165706 142876 165712 142888
rect 165764 142876 165770 142928
rect 219406 142916 219434 143024
rect 222102 142916 222108 142928
rect 219406 142888 222108 142916
rect 222102 142876 222108 142888
rect 222160 142916 222166 142928
rect 264238 142916 264244 142928
rect 222160 142888 264244 142916
rect 222160 142876 222166 142888
rect 264238 142876 264244 142888
rect 264296 142876 264302 142928
rect 269206 142876 269212 142928
rect 269264 142916 269270 142928
rect 273438 142916 273444 142928
rect 269264 142888 273444 142916
rect 269264 142876 269270 142888
rect 273438 142876 273444 142888
rect 273496 142916 273502 142928
rect 309870 142916 309876 142928
rect 273496 142888 309876 142916
rect 273496 142876 273502 142888
rect 309870 142876 309876 142888
rect 309928 142876 309934 142928
rect 33134 142808 33140 142860
rect 33192 142848 33198 142860
rect 164234 142848 164240 142860
rect 33192 142820 164240 142848
rect 33192 142808 33198 142820
rect 164234 142808 164240 142820
rect 164292 142808 164298 142860
rect 197078 142808 197084 142860
rect 197136 142848 197142 142860
rect 255314 142848 255320 142860
rect 197136 142820 255320 142848
rect 197136 142808 197142 142820
rect 255314 142808 255320 142820
rect 255372 142808 255378 142860
rect 283098 142808 283104 142860
rect 283156 142848 283162 142860
rect 376018 142848 376024 142860
rect 283156 142820 376024 142848
rect 283156 142808 283162 142820
rect 376018 142808 376024 142820
rect 376076 142808 376082 142860
rect 187694 142060 187700 142112
rect 187752 142100 187758 142112
rect 283006 142100 283012 142112
rect 187752 142072 283012 142100
rect 187752 142060 187758 142072
rect 283006 142060 283012 142072
rect 283064 142060 283070 142112
rect 194778 141992 194784 142044
rect 194836 142032 194842 142044
rect 289170 142032 289176 142044
rect 194836 142004 289176 142032
rect 194836 141992 194842 142004
rect 289170 141992 289176 142004
rect 289228 141992 289234 142044
rect 204346 141924 204352 141976
rect 204404 141964 204410 141976
rect 278130 141964 278136 141976
rect 204404 141936 278136 141964
rect 204404 141924 204410 141936
rect 278130 141924 278136 141936
rect 278188 141924 278194 141976
rect 171226 141896 171232 141908
rect 161446 141868 171232 141896
rect 121454 141516 121460 141568
rect 121512 141556 121518 141568
rect 161446 141556 161474 141868
rect 171226 141856 171232 141868
rect 171284 141896 171290 141908
rect 234614 141896 234620 141908
rect 171284 141868 234620 141896
rect 171284 141856 171290 141868
rect 234614 141856 234620 141868
rect 234672 141856 234678 141908
rect 183646 141788 183652 141840
rect 183704 141828 183710 141840
rect 245194 141828 245200 141840
rect 183704 141800 245200 141828
rect 183704 141788 183710 141800
rect 245194 141788 245200 141800
rect 245252 141788 245258 141840
rect 189258 141720 189264 141772
rect 189316 141760 189322 141772
rect 190362 141760 190368 141772
rect 189316 141732 190368 141760
rect 189316 141720 189322 141732
rect 190362 141720 190368 141732
rect 190420 141760 190426 141772
rect 249058 141760 249064 141772
rect 190420 141732 249064 141760
rect 190420 141720 190426 141732
rect 249058 141720 249064 141732
rect 249116 141720 249122 141772
rect 205818 141652 205824 141704
rect 205876 141692 205882 141704
rect 265342 141692 265348 141704
rect 205876 141664 265348 141692
rect 205876 141652 205882 141664
rect 265342 141652 265348 141664
rect 265400 141652 265406 141704
rect 179138 141584 179144 141636
rect 179196 141624 179202 141636
rect 223114 141624 223120 141636
rect 179196 141596 223120 141624
rect 179196 141584 179202 141596
rect 223114 141584 223120 141596
rect 223172 141584 223178 141636
rect 121512 141528 161474 141556
rect 121512 141516 121518 141528
rect 178218 141516 178224 141568
rect 178276 141556 178282 141568
rect 179046 141556 179052 141568
rect 178276 141528 179052 141556
rect 178276 141516 178282 141528
rect 179046 141516 179052 141528
rect 179104 141556 179110 141568
rect 218698 141556 218704 141568
rect 179104 141528 218704 141556
rect 179104 141516 179110 141528
rect 218698 141516 218704 141528
rect 218756 141516 218762 141568
rect 243814 141516 243820 141568
rect 243872 141556 243878 141568
rect 323578 141556 323584 141568
rect 243872 141528 323584 141556
rect 243872 141516 243878 141528
rect 323578 141516 323584 141528
rect 323636 141516 323642 141568
rect 44174 141448 44180 141500
rect 44232 141488 44238 141500
rect 166258 141488 166264 141500
rect 44232 141460 166264 141488
rect 44232 141448 44238 141460
rect 166258 141448 166264 141460
rect 166316 141448 166322 141500
rect 177574 141448 177580 141500
rect 177632 141488 177638 141500
rect 179230 141488 179236 141500
rect 177632 141460 179236 141488
rect 177632 141448 177638 141460
rect 179230 141448 179236 141460
rect 179288 141488 179294 141500
rect 233878 141488 233884 141500
rect 179288 141460 233884 141488
rect 179288 141448 179294 141460
rect 233878 141448 233884 141460
rect 233936 141448 233942 141500
rect 245194 141448 245200 141500
rect 245252 141488 245258 141500
rect 266998 141488 267004 141500
rect 245252 141460 267004 141488
rect 245252 141448 245258 141460
rect 266998 141448 267004 141460
rect 267056 141448 267062 141500
rect 289170 141448 289176 141500
rect 289228 141488 289234 141500
rect 415394 141488 415400 141500
rect 289228 141460 415400 141488
rect 289228 141448 289234 141460
rect 415394 141448 415400 141460
rect 415452 141448 415458 141500
rect 31018 141380 31024 141432
rect 31076 141420 31082 141432
rect 164510 141420 164516 141432
rect 31076 141392 164516 141420
rect 31076 141380 31082 141392
rect 164510 141380 164516 141392
rect 164568 141380 164574 141432
rect 206922 141380 206928 141432
rect 206980 141420 206986 141432
rect 267918 141420 267924 141432
rect 206980 141392 267924 141420
rect 206980 141380 206986 141392
rect 267918 141380 267924 141392
rect 267976 141380 267982 141432
rect 278130 141380 278136 141432
rect 278188 141420 278194 141432
rect 547138 141420 547144 141432
rect 278188 141392 547144 141420
rect 278188 141380 278194 141392
rect 547138 141380 547144 141392
rect 547196 141380 547202 141432
rect 205910 140836 205916 140888
rect 205968 140876 205974 140888
rect 206922 140876 206928 140888
rect 205968 140848 206928 140876
rect 205968 140836 205974 140848
rect 206922 140836 206928 140848
rect 206980 140836 206986 140888
rect 205818 140768 205824 140820
rect 205876 140808 205882 140820
rect 206462 140808 206468 140820
rect 205876 140780 206468 140808
rect 205876 140768 205882 140780
rect 206462 140768 206468 140780
rect 206520 140768 206526 140820
rect 190638 140700 190644 140752
rect 190696 140740 190702 140752
rect 285030 140740 285036 140752
rect 190696 140712 285036 140740
rect 190696 140700 190702 140712
rect 285030 140700 285036 140712
rect 285088 140700 285094 140752
rect 197630 140632 197636 140684
rect 197688 140672 197694 140684
rect 272610 140672 272616 140684
rect 197688 140644 272616 140672
rect 197688 140632 197694 140644
rect 272610 140632 272616 140644
rect 272668 140632 272674 140684
rect 167270 140564 167276 140616
rect 167328 140604 167334 140616
rect 229462 140604 229468 140616
rect 167328 140576 229468 140604
rect 167328 140564 167334 140576
rect 229462 140564 229468 140576
rect 229520 140564 229526 140616
rect 184934 140496 184940 140548
rect 184992 140536 184998 140548
rect 246850 140536 246856 140548
rect 184992 140508 246856 140536
rect 184992 140496 184998 140508
rect 246850 140496 246856 140508
rect 246908 140536 246914 140548
rect 246908 140508 248414 140536
rect 246908 140496 246914 140508
rect 167362 140428 167368 140480
rect 167420 140468 167426 140480
rect 227254 140468 227260 140480
rect 167420 140440 227260 140468
rect 167420 140428 167426 140440
rect 227254 140428 227260 140440
rect 227312 140428 227318 140480
rect 169938 140360 169944 140412
rect 169996 140400 170002 140412
rect 170398 140400 170404 140412
rect 169996 140372 170404 140400
rect 169996 140360 170002 140372
rect 170398 140360 170404 140372
rect 170456 140400 170462 140412
rect 225690 140400 225696 140412
rect 170456 140372 225696 140400
rect 170456 140360 170462 140372
rect 225690 140360 225696 140372
rect 225748 140360 225754 140412
rect 169754 140292 169760 140344
rect 169812 140332 169818 140344
rect 170030 140332 170036 140344
rect 169812 140304 170036 140332
rect 169812 140292 169818 140304
rect 170030 140292 170036 140304
rect 170088 140332 170094 140344
rect 222838 140332 222844 140344
rect 170088 140304 222844 140332
rect 170088 140292 170094 140304
rect 222838 140292 222844 140304
rect 222896 140292 222902 140344
rect 115198 140156 115204 140208
rect 115256 140196 115262 140208
rect 171870 140196 171876 140208
rect 115256 140168 171876 140196
rect 115256 140156 115262 140168
rect 171870 140156 171876 140168
rect 171928 140156 171934 140208
rect 248386 140196 248414 140508
rect 302878 140196 302884 140208
rect 248386 140168 302884 140196
rect 302878 140156 302884 140168
rect 302936 140156 302942 140208
rect 40034 140088 40040 140140
rect 40092 140128 40098 140140
rect 165154 140128 165160 140140
rect 40092 140100 165160 140128
rect 40092 140088 40098 140100
rect 165154 140088 165160 140100
rect 165212 140088 165218 140140
rect 285030 140088 285036 140140
rect 285088 140128 285094 140140
rect 363598 140128 363604 140140
rect 285088 140100 363604 140128
rect 285088 140088 285094 140100
rect 363598 140088 363604 140100
rect 363656 140088 363662 140140
rect 17218 140020 17224 140072
rect 17276 140060 17282 140072
rect 163498 140060 163504 140072
rect 17276 140032 163504 140060
rect 17276 140020 17282 140032
rect 163498 140020 163504 140032
rect 163556 140020 163562 140072
rect 272610 140020 272616 140072
rect 272668 140060 272674 140072
rect 465074 140060 465080 140072
rect 272668 140032 465080 140060
rect 272668 140020 272674 140032
rect 465074 140020 465080 140032
rect 465132 140020 465138 140072
rect 167270 139408 167276 139460
rect 167328 139448 167334 139460
rect 167638 139448 167644 139460
rect 167328 139420 167644 139448
rect 167328 139408 167334 139420
rect 167638 139408 167644 139420
rect 167696 139408 167702 139460
rect 186590 139340 186596 139392
rect 186648 139380 186654 139392
rect 274818 139380 274824 139392
rect 186648 139352 274824 139380
rect 186648 139340 186654 139352
rect 274818 139340 274824 139352
rect 274876 139380 274882 139392
rect 275370 139380 275376 139392
rect 274876 139352 275376 139380
rect 274876 139340 274882 139352
rect 275370 139340 275376 139352
rect 275428 139340 275434 139392
rect 193398 139272 193404 139324
rect 193456 139312 193462 139324
rect 271966 139312 271972 139324
rect 193456 139284 271972 139312
rect 193456 139272 193462 139284
rect 271966 139272 271972 139284
rect 272024 139272 272030 139324
rect 205082 139204 205088 139256
rect 205140 139244 205146 139256
rect 269022 139244 269028 139256
rect 205140 139216 269028 139244
rect 205140 139204 205146 139216
rect 269022 139204 269028 139216
rect 269080 139204 269086 139256
rect 168098 139136 168104 139188
rect 168156 139176 168162 139188
rect 227990 139176 227996 139188
rect 168156 139148 227996 139176
rect 168156 139136 168162 139148
rect 227990 139136 227996 139148
rect 228048 139136 228054 139188
rect 179506 139068 179512 139120
rect 179564 139108 179570 139120
rect 226242 139108 226248 139120
rect 179564 139080 226248 139108
rect 179564 139068 179570 139080
rect 226242 139068 226248 139080
rect 226300 139068 226306 139120
rect 115934 138796 115940 138848
rect 115992 138836 115998 138848
rect 171318 138836 171324 138848
rect 115992 138808 171324 138836
rect 115992 138796 115998 138808
rect 171318 138796 171324 138808
rect 171376 138796 171382 138848
rect 275370 138796 275376 138848
rect 275428 138836 275434 138848
rect 314010 138836 314016 138848
rect 275428 138808 314016 138836
rect 275428 138796 275434 138808
rect 314010 138796 314016 138808
rect 314068 138796 314074 138848
rect 62114 138728 62120 138780
rect 62172 138768 62178 138780
rect 167362 138768 167368 138780
rect 62172 138740 167368 138768
rect 62172 138728 62178 138740
rect 167362 138728 167368 138740
rect 167420 138728 167426 138780
rect 271966 138728 271972 138780
rect 272024 138768 272030 138780
rect 399478 138768 399484 138780
rect 272024 138740 399484 138768
rect 272024 138728 272030 138740
rect 399478 138728 399484 138740
rect 399536 138728 399542 138780
rect 52454 138660 52460 138712
rect 52512 138700 52518 138712
rect 165798 138700 165804 138712
rect 52512 138672 165804 138700
rect 52512 138660 52518 138672
rect 165798 138660 165804 138672
rect 165856 138660 165862 138712
rect 269022 138660 269028 138712
rect 269080 138700 269086 138712
rect 554774 138700 554780 138712
rect 269080 138672 554780 138700
rect 269080 138660 269086 138672
rect 554774 138660 554780 138672
rect 554832 138660 554838 138712
rect 167730 137980 167736 138032
rect 167788 138020 167794 138032
rect 168098 138020 168104 138032
rect 167788 137992 168104 138020
rect 167788 137980 167794 137992
rect 168098 137980 168104 137992
rect 168156 137980 168162 138032
rect 194686 137912 194692 137964
rect 194744 137952 194750 137964
rect 285766 137952 285772 137964
rect 194744 137924 285772 137952
rect 194744 137912 194750 137924
rect 285766 137912 285772 137924
rect 285824 137912 285830 137964
rect 205726 137844 205732 137896
rect 205784 137884 205790 137896
rect 272242 137884 272248 137896
rect 205784 137856 272248 137884
rect 205784 137844 205790 137856
rect 272242 137844 272248 137856
rect 272300 137844 272306 137896
rect 146294 137300 146300 137352
rect 146352 137340 146358 137352
rect 173250 137340 173256 137352
rect 146352 137312 173256 137340
rect 146352 137300 146358 137312
rect 173250 137300 173256 137312
rect 173308 137300 173314 137352
rect 283006 137300 283012 137352
rect 283064 137340 283070 137352
rect 338114 137340 338120 137352
rect 283064 137312 338120 137340
rect 283064 137300 283070 137312
rect 338114 137300 338120 137312
rect 338172 137300 338178 137352
rect 26234 137232 26240 137284
rect 26292 137272 26298 137284
rect 164418 137272 164424 137284
rect 26292 137244 164424 137272
rect 26292 137232 26298 137244
rect 164418 137232 164424 137244
rect 164476 137232 164482 137284
rect 180426 137232 180432 137284
rect 180484 137272 180490 137284
rect 220078 137272 220084 137284
rect 180484 137244 220084 137272
rect 180484 137232 180490 137244
rect 220078 137232 220084 137244
rect 220136 137232 220142 137284
rect 285766 137232 285772 137284
rect 285824 137272 285830 137284
rect 419534 137272 419540 137284
rect 285824 137244 419540 137272
rect 285824 137232 285830 137244
rect 419534 137232 419540 137244
rect 419592 137232 419598 137284
rect 272242 136620 272248 136672
rect 272300 136660 272306 136672
rect 564434 136660 564440 136672
rect 272300 136632 564440 136660
rect 272300 136620 272306 136632
rect 564434 136620 564440 136632
rect 564492 136620 564498 136672
rect 196986 136552 196992 136604
rect 197044 136592 197050 136604
rect 261570 136592 261576 136604
rect 197044 136564 261576 136592
rect 197044 136552 197050 136564
rect 261570 136552 261576 136564
rect 261628 136592 261634 136604
rect 262122 136592 262128 136604
rect 261628 136564 262128 136592
rect 261628 136552 261634 136564
rect 262122 136552 262128 136564
rect 262180 136552 262186 136604
rect 205634 136484 205640 136536
rect 205692 136524 205698 136536
rect 270862 136524 270868 136536
rect 205692 136496 270868 136524
rect 205692 136484 205698 136496
rect 270862 136484 270868 136496
rect 270920 136524 270926 136536
rect 271782 136524 271788 136536
rect 270920 136496 271788 136524
rect 270920 136484 270926 136496
rect 271782 136484 271788 136496
rect 271840 136484 271846 136536
rect 189166 136416 189172 136468
rect 189224 136456 189230 136468
rect 249610 136456 249616 136468
rect 189224 136428 249616 136456
rect 189224 136416 189230 136428
rect 249610 136416 249616 136428
rect 249668 136416 249674 136468
rect 219434 136348 219440 136400
rect 219492 136388 219498 136400
rect 220078 136388 220084 136400
rect 219492 136360 220084 136388
rect 219492 136348 219498 136360
rect 220078 136348 220084 136360
rect 220136 136388 220142 136400
rect 238018 136388 238024 136400
rect 220136 136360 238024 136388
rect 220136 136348 220142 136360
rect 238018 136348 238024 136360
rect 238076 136348 238082 136400
rect 249610 136008 249616 136060
rect 249668 136048 249674 136060
rect 351914 136048 351920 136060
rect 249668 136020 351920 136048
rect 249668 136008 249674 136020
rect 351914 136008 351920 136020
rect 351972 136008 351978 136060
rect 262122 135940 262128 135992
rect 262180 135980 262186 135992
rect 440234 135980 440240 135992
rect 262180 135952 440240 135980
rect 262180 135940 262186 135952
rect 440234 135940 440240 135952
rect 440292 135940 440298 135992
rect 4798 135872 4804 135924
rect 4856 135912 4862 135924
rect 161750 135912 161756 135924
rect 4856 135884 161756 135912
rect 4856 135872 4862 135884
rect 161750 135872 161756 135884
rect 161808 135872 161814 135924
rect 180518 135872 180524 135924
rect 180576 135912 180582 135924
rect 223574 135912 223580 135924
rect 180576 135884 223580 135912
rect 180576 135872 180582 135884
rect 223574 135872 223580 135884
rect 223632 135872 223638 135924
rect 271782 135872 271788 135924
rect 271840 135912 271846 135924
rect 571978 135912 571984 135924
rect 271840 135884 571984 135912
rect 271840 135872 271846 135884
rect 571978 135872 571984 135884
rect 572036 135872 572042 135924
rect 191558 135192 191564 135244
rect 191616 135232 191622 135244
rect 250990 135232 250996 135244
rect 191616 135204 250996 135232
rect 191616 135192 191622 135204
rect 250990 135192 250996 135204
rect 251048 135192 251054 135244
rect 91094 134580 91100 134632
rect 91152 134620 91158 134632
rect 168374 134620 168380 134632
rect 91152 134592 168380 134620
rect 91152 134580 91158 134592
rect 168374 134580 168380 134592
rect 168432 134580 168438 134632
rect 181898 134580 181904 134632
rect 181956 134620 181962 134632
rect 241514 134620 241520 134632
rect 181956 134592 241520 134620
rect 181956 134580 181962 134592
rect 241514 134580 241520 134592
rect 241572 134580 241578 134632
rect 250990 134580 250996 134632
rect 251048 134620 251054 134632
rect 369854 134620 369860 134632
rect 251048 134592 369860 134620
rect 251048 134580 251054 134592
rect 369854 134580 369860 134592
rect 369912 134580 369918 134632
rect 8294 134512 8300 134564
rect 8352 134552 8358 134564
rect 162854 134552 162860 134564
rect 8352 134524 162860 134552
rect 8352 134512 8358 134524
rect 162854 134512 162860 134524
rect 162912 134512 162918 134564
rect 208118 134512 208124 134564
rect 208176 134552 208182 134564
rect 575474 134552 575480 134564
rect 208176 134524 575480 134552
rect 208176 134512 208182 134524
rect 575474 134512 575480 134524
rect 575532 134512 575538 134564
rect 191466 133832 191472 133884
rect 191524 133872 191530 133884
rect 285674 133872 285680 133884
rect 191524 133844 285680 133872
rect 191524 133832 191530 133844
rect 285674 133832 285680 133844
rect 285732 133832 285738 133884
rect 197446 133764 197452 133816
rect 197504 133804 197510 133816
rect 291930 133804 291936 133816
rect 197504 133776 291936 133804
rect 197504 133764 197510 133776
rect 291930 133764 291936 133776
rect 291988 133764 291994 133816
rect 186314 133696 186320 133748
rect 186372 133736 186378 133748
rect 246022 133736 246028 133748
rect 186372 133708 246028 133736
rect 186372 133696 186378 133708
rect 246022 133696 246028 133708
rect 246080 133696 246086 133748
rect 246022 133288 246028 133340
rect 246080 133328 246086 133340
rect 246942 133328 246948 133340
rect 246080 133300 246948 133328
rect 246080 133288 246086 133300
rect 246942 133288 246948 133300
rect 247000 133328 247006 133340
rect 320174 133328 320180 133340
rect 247000 133300 320180 133328
rect 247000 133288 247006 133300
rect 320174 133288 320180 133300
rect 320232 133288 320238 133340
rect 97994 133220 98000 133272
rect 98052 133260 98058 133272
rect 169754 133260 169760 133272
rect 98052 133232 169760 133260
rect 98052 133220 98058 133232
rect 169754 133220 169760 133232
rect 169812 133220 169818 133272
rect 285674 133220 285680 133272
rect 285732 133260 285738 133272
rect 376754 133260 376760 133272
rect 285732 133232 376760 133260
rect 285732 133220 285738 133232
rect 376754 133220 376760 133232
rect 376812 133220 376818 133272
rect 48314 133152 48320 133204
rect 48372 133192 48378 133204
rect 166166 133192 166172 133204
rect 48372 133164 166172 133192
rect 48372 133152 48378 133164
rect 166166 133152 166172 133164
rect 166224 133152 166230 133204
rect 166258 133152 166264 133204
rect 166316 133192 166322 133204
rect 174722 133192 174728 133204
rect 166316 133164 174728 133192
rect 166316 133152 166322 133164
rect 174722 133152 174728 133164
rect 174780 133152 174786 133204
rect 291930 133152 291936 133204
rect 291988 133192 291994 133204
rect 455414 133192 455420 133204
rect 291988 133164 455420 133192
rect 291988 133152 291994 133164
rect 455414 133152 455420 133164
rect 455472 133152 455478 133204
rect 192018 132404 192024 132456
rect 192076 132444 192082 132456
rect 287790 132444 287796 132456
rect 192076 132416 287796 132444
rect 192076 132404 192082 132416
rect 287790 132404 287796 132416
rect 287848 132404 287854 132456
rect 198918 132336 198924 132388
rect 198976 132376 198982 132388
rect 293218 132376 293224 132388
rect 198976 132348 293224 132376
rect 198976 132336 198982 132348
rect 293218 132336 293224 132348
rect 293276 132336 293282 132388
rect 186498 132268 186504 132320
rect 186556 132308 186562 132320
rect 247034 132308 247040 132320
rect 186556 132280 247040 132308
rect 186556 132268 186562 132280
rect 247034 132268 247040 132280
rect 247092 132268 247098 132320
rect 247034 131860 247040 131912
rect 247092 131900 247098 131912
rect 248322 131900 248328 131912
rect 247092 131872 248328 131900
rect 247092 131860 247098 131872
rect 248322 131860 248328 131872
rect 248380 131900 248386 131912
rect 301498 131900 301504 131912
rect 248380 131872 301504 131900
rect 248380 131860 248386 131872
rect 301498 131860 301504 131872
rect 301556 131860 301562 131912
rect 287790 131792 287796 131844
rect 287848 131832 287854 131844
rect 387794 131832 387800 131844
rect 287848 131804 387800 131832
rect 287848 131792 287854 131804
rect 387794 131792 387800 131804
rect 387852 131792 387858 131844
rect 110506 131724 110512 131776
rect 110564 131764 110570 131776
rect 170858 131764 170864 131776
rect 110564 131736 170864 131764
rect 110564 131724 110570 131736
rect 170858 131724 170864 131736
rect 170916 131724 170922 131776
rect 177758 131724 177764 131776
rect 177816 131764 177822 131776
rect 186314 131764 186320 131776
rect 177816 131736 186320 131764
rect 177816 131724 177822 131736
rect 186314 131724 186320 131736
rect 186372 131724 186378 131776
rect 293218 131724 293224 131776
rect 293276 131764 293282 131776
rect 468478 131764 468484 131776
rect 293276 131736 468484 131764
rect 293276 131724 293282 131736
rect 468478 131724 468484 131736
rect 468536 131724 468542 131776
rect 193306 131044 193312 131096
rect 193364 131084 193370 131096
rect 255222 131084 255228 131096
rect 193364 131056 255228 131084
rect 193364 131044 193370 131056
rect 255222 131044 255228 131056
rect 255280 131044 255286 131096
rect 169018 130364 169024 130416
rect 169076 130404 169082 130416
rect 176102 130404 176108 130416
rect 169076 130376 176108 130404
rect 169076 130364 169082 130376
rect 176102 130364 176108 130376
rect 176160 130364 176166 130416
rect 255222 130364 255228 130416
rect 255280 130404 255286 130416
rect 408494 130404 408500 130416
rect 255280 130376 408500 130404
rect 255280 130364 255286 130376
rect 408494 130364 408500 130376
rect 408552 130364 408558 130416
rect 195698 129684 195704 129736
rect 195756 129724 195762 129736
rect 268194 129724 268200 129736
rect 195756 129696 268200 129724
rect 195756 129684 195762 129696
rect 268194 129684 268200 129696
rect 268252 129724 268258 129736
rect 269022 129724 269028 129736
rect 268252 129696 269028 129724
rect 268252 129684 268258 129696
rect 269022 129684 269028 129696
rect 269080 129684 269086 129736
rect 199654 129616 199660 129668
rect 199712 129656 199718 129668
rect 270402 129656 270408 129668
rect 199712 129628 270408 129656
rect 199712 129616 199718 129628
rect 270402 129616 270408 129628
rect 270460 129616 270466 129668
rect 117314 129072 117320 129124
rect 117372 129112 117378 129124
rect 171778 129112 171784 129124
rect 117372 129084 171784 129112
rect 117372 129072 117378 129084
rect 171778 129072 171784 129084
rect 171836 129072 171842 129124
rect 269022 129072 269028 129124
rect 269080 129112 269086 129124
rect 422938 129112 422944 129124
rect 269080 129084 422944 129112
rect 269080 129072 269086 129084
rect 422938 129072 422944 129084
rect 422996 129072 423002 129124
rect 66254 129004 66260 129056
rect 66312 129044 66318 129056
rect 168282 129044 168288 129056
rect 66312 129016 168288 129044
rect 66312 129004 66318 129016
rect 168282 129004 168288 129016
rect 168340 129004 168346 129056
rect 181990 129004 181996 129056
rect 182048 129044 182054 129056
rect 237374 129044 237380 129056
rect 182048 129016 237380 129044
rect 182048 129004 182054 129016
rect 237374 129004 237380 129016
rect 237432 129004 237438 129056
rect 270402 129004 270408 129056
rect 270460 129044 270466 129056
rect 480254 129044 480260 129056
rect 270460 129016 480260 129044
rect 270460 129004 270466 129016
rect 480254 129004 480260 129016
rect 480312 129004 480318 129056
rect 200114 128256 200120 128308
rect 200172 128296 200178 128308
rect 274082 128296 274088 128308
rect 200172 128268 274088 128296
rect 200172 128256 200178 128268
rect 274082 128256 274088 128268
rect 274140 128296 274146 128308
rect 274542 128296 274548 128308
rect 274140 128268 274548 128296
rect 274140 128256 274146 128268
rect 274542 128256 274548 128268
rect 274600 128256 274606 128308
rect 195974 128188 195980 128240
rect 196032 128228 196038 128240
rect 256050 128228 256056 128240
rect 196032 128200 256056 128228
rect 196032 128188 196038 128200
rect 256050 128188 256056 128200
rect 256108 128188 256114 128240
rect 122098 127644 122104 127696
rect 122156 127684 122162 127696
rect 172422 127684 172428 127696
rect 122156 127656 172428 127684
rect 122156 127644 122162 127656
rect 172422 127644 172428 127656
rect 172480 127644 172486 127696
rect 256050 127644 256056 127696
rect 256108 127684 256114 127696
rect 256602 127684 256608 127696
rect 256108 127656 256608 127684
rect 256108 127644 256114 127656
rect 256602 127644 256608 127656
rect 256660 127684 256666 127696
rect 444374 127684 444380 127696
rect 256660 127656 444380 127684
rect 256660 127644 256666 127656
rect 444374 127644 444380 127656
rect 444432 127644 444438 127696
rect 69014 127576 69020 127628
rect 69072 127616 69078 127628
rect 167730 127616 167736 127628
rect 69072 127588 167736 127616
rect 69072 127576 69078 127588
rect 167730 127576 167736 127588
rect 167788 127576 167794 127628
rect 274082 127576 274088 127628
rect 274140 127616 274146 127628
rect 490006 127616 490012 127628
rect 274140 127588 490012 127616
rect 274140 127576 274146 127588
rect 490006 127576 490012 127588
rect 490064 127576 490070 127628
rect 186406 126896 186412 126948
rect 186464 126936 186470 126948
rect 280798 126936 280804 126948
rect 186464 126908 280804 126936
rect 186464 126896 186470 126908
rect 280798 126896 280804 126908
rect 280856 126936 280862 126948
rect 281442 126936 281448 126948
rect 280856 126908 281448 126936
rect 280856 126896 280862 126908
rect 281442 126896 281448 126908
rect 281500 126896 281506 126948
rect 198550 126828 198556 126880
rect 198608 126868 198614 126880
rect 288434 126868 288440 126880
rect 198608 126840 288440 126868
rect 198608 126828 198614 126840
rect 288434 126828 288440 126840
rect 288492 126868 288498 126880
rect 289722 126868 289728 126880
rect 288492 126840 289728 126868
rect 288492 126828 288498 126840
rect 289722 126828 289728 126840
rect 289780 126828 289786 126880
rect 191926 126760 191932 126812
rect 191984 126800 191990 126812
rect 253474 126800 253480 126812
rect 191984 126772 253480 126800
rect 191984 126760 191990 126772
rect 253474 126760 253480 126772
rect 253532 126800 253538 126812
rect 253842 126800 253848 126812
rect 253532 126772 253848 126800
rect 253532 126760 253538 126772
rect 253842 126760 253848 126772
rect 253900 126760 253906 126812
rect 281442 126352 281448 126404
rect 281500 126392 281506 126404
rect 307846 126392 307852 126404
rect 281500 126364 307852 126392
rect 281500 126352 281506 126364
rect 307846 126352 307852 126364
rect 307904 126352 307910 126404
rect 253474 126284 253480 126336
rect 253532 126324 253538 126336
rect 390554 126324 390560 126336
rect 253532 126296 390560 126324
rect 253532 126284 253538 126296
rect 390554 126284 390560 126296
rect 390612 126284 390618 126336
rect 289722 126216 289728 126268
rect 289780 126256 289786 126268
rect 458174 126256 458180 126268
rect 289780 126228 458180 126256
rect 289780 126216 289786 126228
rect 458174 126216 458180 126228
rect 458232 126216 458238 126268
rect 176562 125536 176568 125588
rect 176620 125576 176626 125588
rect 180150 125576 180156 125588
rect 176620 125548 180156 125576
rect 176620 125536 176626 125548
rect 180150 125536 180156 125548
rect 180208 125536 180214 125588
rect 198734 125536 198740 125588
rect 198792 125576 198798 125588
rect 274726 125576 274732 125588
rect 198792 125548 274732 125576
rect 198792 125536 198798 125548
rect 274726 125536 274732 125548
rect 274784 125576 274790 125588
rect 275370 125576 275376 125588
rect 274784 125548 275376 125576
rect 274784 125536 274790 125548
rect 275370 125536 275376 125548
rect 275428 125536 275434 125588
rect 189074 125468 189080 125520
rect 189132 125508 189138 125520
rect 251082 125508 251088 125520
rect 189132 125480 251088 125508
rect 189132 125468 189138 125480
rect 251082 125468 251088 125480
rect 251140 125468 251146 125520
rect 102134 124924 102140 124976
rect 102192 124964 102198 124976
rect 170398 124964 170404 124976
rect 102192 124936 170404 124964
rect 102192 124924 102198 124936
rect 170398 124924 170404 124936
rect 170456 124924 170462 124976
rect 251082 124924 251088 124976
rect 251140 124964 251146 124976
rect 337378 124964 337384 124976
rect 251140 124936 337384 124964
rect 251140 124924 251146 124936
rect 337378 124924 337384 124936
rect 337436 124924 337442 124976
rect 56594 124856 56600 124908
rect 56652 124896 56658 124908
rect 166074 124896 166080 124908
rect 56652 124868 166080 124896
rect 56652 124856 56658 124868
rect 166074 124856 166080 124868
rect 166132 124856 166138 124908
rect 275370 124856 275376 124908
rect 275428 124896 275434 124908
rect 476114 124896 476120 124908
rect 275428 124868 476120 124896
rect 275428 124856 275434 124868
rect 476114 124856 476120 124868
rect 476172 124856 476178 124908
rect 192938 124108 192944 124160
rect 192996 124148 193002 124160
rect 252462 124148 252468 124160
rect 192996 124120 252468 124148
rect 192996 124108 193002 124120
rect 252462 124108 252468 124120
rect 252520 124108 252526 124160
rect 201586 124040 201592 124092
rect 201644 124080 201650 124092
rect 261478 124080 261484 124092
rect 201644 124052 261484 124080
rect 201644 124040 201650 124052
rect 261478 124040 261484 124052
rect 261536 124080 261542 124092
rect 262122 124080 262128 124092
rect 261536 124052 262128 124080
rect 261536 124040 261542 124052
rect 262122 124040 262128 124052
rect 262180 124040 262186 124092
rect 252462 123496 252468 123548
rect 252520 123536 252526 123548
rect 394694 123536 394700 123548
rect 252520 123508 394700 123536
rect 252520 123496 252526 123508
rect 394694 123496 394700 123508
rect 394752 123496 394758 123548
rect 86954 123428 86960 123480
rect 87012 123468 87018 123480
rect 169478 123468 169484 123480
rect 87012 123440 169484 123468
rect 87012 123428 87018 123440
rect 169478 123428 169484 123440
rect 169536 123428 169542 123480
rect 262122 123428 262128 123480
rect 262180 123468 262186 123480
rect 503714 123468 503720 123480
rect 262180 123440 503720 123468
rect 262180 123428 262186 123440
rect 503714 123428 503720 123440
rect 503772 123428 503778 123480
rect 194502 122068 194508 122120
rect 194560 122108 194566 122120
rect 412634 122108 412640 122120
rect 194560 122080 412640 122108
rect 194560 122068 194566 122080
rect 412634 122068 412640 122080
rect 412692 122068 412698 122120
rect 60826 120708 60832 120760
rect 60884 120748 60890 120760
rect 167086 120748 167092 120760
rect 60884 120720 167092 120748
rect 60884 120708 60890 120720
rect 167086 120708 167092 120720
rect 167144 120708 167150 120760
rect 22738 119348 22744 119400
rect 22796 119388 22802 119400
rect 163222 119388 163228 119400
rect 22796 119360 163228 119388
rect 22796 119348 22802 119360
rect 163222 119348 163228 119360
rect 163280 119348 163286 119400
rect 184566 119348 184572 119400
rect 184624 119388 184630 119400
rect 273254 119388 273260 119400
rect 184624 119360 273260 119388
rect 184624 119348 184630 119360
rect 273254 119348 273260 119360
rect 273312 119348 273318 119400
rect 162854 117988 162860 118040
rect 162912 118028 162918 118040
rect 173986 118028 173992 118040
rect 162912 118000 173992 118028
rect 162912 117988 162918 118000
rect 173986 117988 173992 118000
rect 174044 117988 174050 118040
rect 24118 117920 24124 117972
rect 24176 117960 24182 117972
rect 163038 117960 163044 117972
rect 24176 117932 163044 117960
rect 24176 117920 24182 117932
rect 163038 117920 163044 117932
rect 163096 117920 163102 117972
rect 193214 117240 193220 117292
rect 193272 117280 193278 117292
rect 253382 117280 253388 117292
rect 193272 117252 253388 117280
rect 193272 117240 193278 117252
rect 253382 117240 253388 117252
rect 253440 117240 253446 117292
rect 39298 116560 39304 116612
rect 39356 116600 39362 116612
rect 164694 116600 164700 116612
rect 39356 116572 164700 116600
rect 39356 116560 39362 116572
rect 164694 116560 164700 116572
rect 164752 116560 164758 116612
rect 253382 116560 253388 116612
rect 253440 116600 253446 116612
rect 404354 116600 404360 116612
rect 253440 116572 404360 116600
rect 253440 116560 253446 116572
rect 404354 116560 404360 116572
rect 404412 116560 404418 116612
rect 43438 115200 43444 115252
rect 43496 115240 43502 115252
rect 166810 115240 166816 115252
rect 43496 115212 166816 115240
rect 43496 115200 43502 115212
rect 166810 115200 166816 115212
rect 166868 115200 166874 115252
rect 279418 113092 279424 113144
rect 279476 113132 279482 113144
rect 580166 113132 580172 113144
rect 279476 113104 580172 113132
rect 279476 113092 279482 113104
rect 580166 113092 580172 113104
rect 580224 113092 580230 113144
rect 9674 112412 9680 112464
rect 9732 112452 9738 112464
rect 163406 112452 163412 112464
rect 9732 112424 163412 112452
rect 9732 112412 9738 112424
rect 163406 112412 163412 112424
rect 163464 112412 163470 112464
rect 3142 111732 3148 111784
rect 3200 111772 3206 111784
rect 120810 111772 120816 111784
rect 3200 111744 120816 111772
rect 3200 111732 3206 111744
rect 120810 111732 120816 111744
rect 120868 111732 120874 111784
rect 131114 111052 131120 111104
rect 131172 111092 131178 111104
rect 173066 111092 173072 111104
rect 131172 111064 173072 111092
rect 131172 111052 131178 111064
rect 173066 111052 173072 111064
rect 173124 111052 173130 111104
rect 183462 111052 183468 111104
rect 183520 111092 183526 111104
rect 262214 111092 262220 111104
rect 183520 111064 262220 111092
rect 183520 111052 183526 111064
rect 262214 111052 262220 111064
rect 262272 111052 262278 111104
rect 52546 109692 52552 109744
rect 52604 109732 52610 109744
rect 165614 109732 165620 109744
rect 52604 109704 165620 109732
rect 52604 109692 52610 109704
rect 165614 109692 165620 109704
rect 165672 109692 165678 109744
rect 201126 109692 201132 109744
rect 201184 109732 201190 109744
rect 489178 109732 489184 109744
rect 201184 109704 489184 109732
rect 201184 109692 201190 109704
rect 489178 109692 489184 109704
rect 489236 109692 489242 109744
rect 70394 108264 70400 108316
rect 70452 108304 70458 108316
rect 167454 108304 167460 108316
rect 70452 108276 167460 108304
rect 70452 108264 70458 108276
rect 167454 108264 167460 108276
rect 167512 108264 167518 108316
rect 177298 108264 177304 108316
rect 177356 108304 177362 108316
rect 184290 108304 184296 108316
rect 177356 108276 184296 108304
rect 177356 108264 177362 108276
rect 184290 108264 184296 108276
rect 184348 108264 184354 108316
rect 201218 108264 201224 108316
rect 201276 108304 201282 108316
rect 492674 108304 492680 108316
rect 201276 108276 492680 108304
rect 201276 108264 201282 108276
rect 492674 108264 492680 108276
rect 492732 108264 492738 108316
rect 79318 106904 79324 106956
rect 79376 106944 79382 106956
rect 169202 106944 169208 106956
rect 79376 106916 169208 106944
rect 79376 106904 79382 106916
rect 169202 106904 169208 106916
rect 169260 106904 169266 106956
rect 179046 105612 179052 105664
rect 179104 105652 179110 105664
rect 201586 105652 201592 105664
rect 179104 105624 201592 105652
rect 179104 105612 179110 105624
rect 201586 105612 201592 105624
rect 201644 105612 201650 105664
rect 13814 105544 13820 105596
rect 13872 105584 13878 105596
rect 163130 105584 163136 105596
rect 13872 105556 163136 105584
rect 13872 105544 13878 105556
rect 163130 105544 163136 105556
rect 163188 105544 163194 105596
rect 190362 105544 190368 105596
rect 190420 105584 190426 105596
rect 347774 105584 347780 105596
rect 190420 105556 347780 105584
rect 190420 105544 190426 105556
rect 347774 105544 347780 105556
rect 347832 105544 347838 105596
rect 95234 104116 95240 104168
rect 95292 104156 95298 104168
rect 169846 104156 169852 104168
rect 95292 104128 169852 104156
rect 95292 104116 95298 104128
rect 169846 104116 169852 104128
rect 169904 104116 169910 104168
rect 31754 102756 31760 102808
rect 31812 102796 31818 102808
rect 164602 102796 164608 102808
rect 31812 102768 164608 102796
rect 31812 102756 31818 102768
rect 164602 102756 164608 102768
rect 164660 102756 164666 102808
rect 202690 101396 202696 101448
rect 202748 101436 202754 101448
rect 517514 101436 517520 101448
rect 202748 101408 517520 101436
rect 202748 101396 202754 101408
rect 517514 101396 517520 101408
rect 517572 101396 517578 101448
rect 341518 100648 341524 100700
rect 341576 100688 341582 100700
rect 580166 100688 580172 100700
rect 341576 100660 580172 100688
rect 341576 100648 341582 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 19334 99968 19340 100020
rect 19392 100008 19398 100020
rect 157886 100008 157892 100020
rect 19392 99980 157892 100008
rect 19392 99968 19398 99980
rect 157886 99968 157892 99980
rect 157944 99968 157950 100020
rect 111794 98608 111800 98660
rect 111852 98648 111858 98660
rect 171502 98648 171508 98660
rect 111852 98620 171508 98648
rect 111852 98608 111858 98620
rect 171502 98608 171508 98620
rect 171560 98608 171566 98660
rect 27614 97248 27620 97300
rect 27672 97288 27678 97300
rect 153930 97288 153936 97300
rect 27672 97260 153936 97288
rect 27672 97248 27678 97260
rect 153930 97248 153936 97260
rect 153988 97248 153994 97300
rect 35894 94460 35900 94512
rect 35952 94500 35958 94512
rect 156690 94500 156696 94512
rect 35952 94472 156696 94500
rect 35952 94460 35958 94472
rect 156690 94460 156696 94472
rect 156748 94460 156754 94512
rect 203978 94460 203984 94512
rect 204036 94500 204042 94512
rect 535454 94500 535460 94512
rect 204036 94472 535460 94500
rect 204036 94460 204042 94472
rect 535454 94460 535460 94472
rect 535512 94460 535518 94512
rect 11054 93100 11060 93152
rect 11112 93140 11118 93152
rect 148318 93140 148324 93152
rect 11112 93112 148324 93140
rect 11112 93100 11118 93112
rect 148318 93100 148324 93112
rect 148376 93100 148382 93152
rect 205542 91740 205548 91792
rect 205600 91780 205606 91792
rect 553394 91780 553400 91792
rect 205600 91752 553400 91780
rect 205600 91740 205606 91752
rect 553394 91740 553400 91752
rect 553452 91740 553458 91792
rect 206554 90312 206560 90364
rect 206612 90352 206618 90364
rect 556246 90352 556252 90364
rect 206612 90324 556252 90352
rect 206612 90312 206618 90324
rect 556246 90312 556252 90324
rect 556304 90312 556310 90364
rect 206462 88952 206468 89004
rect 206520 88992 206526 89004
rect 560294 88992 560300 89004
rect 206520 88964 560300 88992
rect 206520 88952 206526 88964
rect 560294 88952 560300 88964
rect 560352 88952 560358 89004
rect 206646 87592 206652 87644
rect 206704 87632 206710 87644
rect 564526 87632 564532 87644
rect 206704 87604 564532 87632
rect 206704 87592 206710 87604
rect 564526 87592 564532 87604
rect 564584 87592 564590 87644
rect 179138 86232 179144 86284
rect 179196 86272 179202 86284
rect 205634 86272 205640 86284
rect 179196 86244 205640 86272
rect 179196 86232 179202 86244
rect 205634 86232 205640 86244
rect 205692 86232 205698 86284
rect 206738 86232 206744 86284
rect 206796 86272 206802 86284
rect 567194 86272 567200 86284
rect 206796 86244 567200 86272
rect 206796 86232 206802 86244
rect 567194 86232 567200 86244
rect 567252 86232 567258 86284
rect 3510 85484 3516 85536
rect 3568 85524 3574 85536
rect 28258 85524 28264 85536
rect 3568 85496 28264 85524
rect 3568 85484 3574 85496
rect 28258 85484 28264 85496
rect 28316 85484 28322 85536
rect 206830 84804 206836 84856
rect 206888 84844 206894 84856
rect 569218 84844 569224 84856
rect 206888 84816 569224 84844
rect 206888 84804 206894 84816
rect 569218 84804 569224 84816
rect 569276 84804 569282 84856
rect 208210 83444 208216 83496
rect 208268 83484 208274 83496
rect 574094 83484 574100 83496
rect 208268 83456 574100 83484
rect 208268 83444 208274 83456
rect 574094 83444 574100 83456
rect 574152 83444 574158 83496
rect 208302 80656 208308 80708
rect 208360 80696 208366 80708
rect 578234 80696 578240 80708
rect 208360 80668 578240 80696
rect 208360 80656 208366 80668
rect 578234 80656 578240 80668
rect 578292 80656 578298 80708
rect 42794 77936 42800 77988
rect 42852 77976 42858 77988
rect 151170 77976 151176 77988
rect 42852 77948 151176 77976
rect 42852 77936 42858 77948
rect 151170 77936 151176 77948
rect 151228 77936 151234 77988
rect 198642 73788 198648 73840
rect 198700 73828 198706 73840
rect 454034 73828 454040 73840
rect 198700 73800 454040 73828
rect 198700 73788 198706 73800
rect 454034 73788 454040 73800
rect 454092 73788 454098 73840
rect 3510 71680 3516 71732
rect 3568 71720 3574 71732
rect 146938 71720 146944 71732
rect 3568 71692 146944 71720
rect 3568 71680 3574 71692
rect 146938 71680 146944 71692
rect 146996 71680 147002 71732
rect 176654 68280 176660 68332
rect 176712 68320 176718 68332
rect 187694 68320 187700 68332
rect 176712 68292 187700 68320
rect 176712 68280 176718 68292
rect 187694 68280 187700 68292
rect 187752 68280 187758 68332
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 155218 59344 155224 59356
rect 3108 59316 155224 59344
rect 3108 59304 3114 59316
rect 155218 59304 155224 59316
rect 155276 59304 155282 59356
rect 177942 58624 177948 58676
rect 178000 58664 178006 58676
rect 191098 58664 191104 58676
rect 178000 58636 191104 58664
rect 178000 58624 178006 58636
rect 191098 58624 191104 58636
rect 191156 58624 191162 58676
rect 3510 45500 3516 45552
rect 3568 45540 3574 45552
rect 156598 45540 156604 45552
rect 3568 45512 156604 45540
rect 3568 45500 3574 45512
rect 156598 45500 156604 45512
rect 156656 45500 156662 45552
rect 204162 37884 204168 37936
rect 204220 37924 204226 37936
rect 525794 37924 525800 37936
rect 204220 37896 525800 37924
rect 204220 37884 204226 37896
rect 525794 37884 525800 37896
rect 525852 37884 525858 37936
rect 206922 36524 206928 36576
rect 206980 36564 206986 36576
rect 568574 36564 568580 36576
rect 206980 36536 568580 36564
rect 206980 36524 206986 36536
rect 568574 36524 568580 36536
rect 568632 36524 568638 36576
rect 201310 35164 201316 35216
rect 201368 35204 201374 35216
rect 499574 35204 499580 35216
rect 201368 35176 499580 35204
rect 201368 35164 201374 35176
rect 499574 35164 499580 35176
rect 499632 35164 499638 35216
rect 204070 33736 204076 33788
rect 204128 33776 204134 33788
rect 524414 33776 524420 33788
rect 204128 33748 524420 33776
rect 204128 33736 204134 33748
rect 524414 33736 524420 33748
rect 524472 33736 524478 33788
rect 2866 33056 2872 33108
rect 2924 33096 2930 33108
rect 11698 33096 11704 33108
rect 2924 33068 11704 33096
rect 2924 33056 2930 33068
rect 11698 33056 11704 33068
rect 11756 33056 11762 33108
rect 176010 28908 176016 28960
rect 176068 28948 176074 28960
rect 176654 28948 176660 28960
rect 176068 28920 176660 28948
rect 176068 28908 176074 28920
rect 176654 28908 176660 28920
rect 176712 28908 176718 28960
rect 334618 20612 334624 20664
rect 334676 20652 334682 20664
rect 580074 20652 580080 20664
rect 334676 20624 580080 20652
rect 334676 20612 334682 20624
rect 580074 20612 580080 20624
rect 580132 20612 580138 20664
rect 205450 18572 205456 18624
rect 205508 18612 205514 18624
rect 539686 18612 539692 18624
rect 205508 18584 539692 18612
rect 205508 18572 205514 18584
rect 539686 18572 539692 18584
rect 539744 18572 539750 18624
rect 38654 17212 38660 17264
rect 38712 17252 38718 17264
rect 165430 17252 165436 17264
rect 38712 17224 165436 17252
rect 38712 17212 38718 17224
rect 165430 17212 165436 17224
rect 165488 17212 165494 17264
rect 197170 17212 197176 17264
rect 197228 17252 197234 17264
rect 433334 17252 433340 17264
rect 197228 17224 433340 17252
rect 197228 17212 197234 17224
rect 433334 17212 433340 17224
rect 433392 17212 433398 17264
rect 202782 15852 202788 15904
rect 202840 15892 202846 15904
rect 505370 15892 505376 15904
rect 202840 15864 505376 15892
rect 202840 15852 202846 15864
rect 505370 15852 505376 15864
rect 505428 15852 505434 15904
rect 88886 14424 88892 14476
rect 88944 14464 88950 14476
rect 168926 14464 168932 14476
rect 88944 14436 168932 14464
rect 88944 14424 88950 14436
rect 168926 14424 168932 14436
rect 168984 14424 168990 14476
rect 25314 13064 25320 13116
rect 25372 13104 25378 13116
rect 164878 13104 164884 13116
rect 25372 13076 164884 13104
rect 25372 13064 25378 13076
rect 164878 13064 164884 13076
rect 164936 13064 164942 13116
rect 143534 11772 143540 11824
rect 143592 11812 143598 11824
rect 144730 11812 144736 11824
rect 143592 11784 144736 11812
rect 143592 11772 143598 11784
rect 144730 11772 144736 11784
rect 144788 11772 144794 11824
rect 15746 11704 15752 11756
rect 15804 11744 15810 11756
rect 163774 11744 163780 11756
rect 15804 11716 163780 11744
rect 15804 11704 15810 11716
rect 163774 11704 163780 11716
rect 163832 11704 163838 11756
rect 20162 10276 20168 10328
rect 20220 10316 20226 10328
rect 124858 10316 124864 10328
rect 20220 10288 124864 10316
rect 20220 10276 20226 10288
rect 124858 10276 124864 10288
rect 124916 10276 124922 10328
rect 190454 10276 190460 10328
rect 190512 10316 190518 10328
rect 376018 10316 376024 10328
rect 190512 10288 376024 10316
rect 190512 10276 190518 10288
rect 376018 10276 376024 10288
rect 376076 10276 376082 10328
rect 195882 9052 195888 9104
rect 195940 9092 195946 9104
rect 422570 9092 422576 9104
rect 195940 9064 422576 9092
rect 195940 9052 195946 9064
rect 422570 9052 422576 9064
rect 422628 9052 422634 9104
rect 197078 8984 197084 9036
rect 197136 9024 197142 9036
rect 433242 9024 433248 9036
rect 197136 8996 433248 9024
rect 197136 8984 197142 8996
rect 433242 8984 433248 8996
rect 433300 8984 433306 9036
rect 103330 8916 103336 8968
rect 103388 8956 103394 8968
rect 170766 8956 170772 8968
rect 103388 8928 170772 8956
rect 103388 8916 103394 8928
rect 170766 8916 170772 8928
rect 170824 8916 170830 8968
rect 196066 8916 196072 8968
rect 196124 8956 196130 8968
rect 443822 8956 443828 8968
rect 196124 8928 443828 8956
rect 196124 8916 196130 8928
rect 443822 8916 443828 8928
rect 443880 8916 443886 8968
rect 73798 7556 73804 7608
rect 73856 7596 73862 7608
rect 167638 7596 167644 7608
rect 73856 7568 167644 7596
rect 73856 7556 73862 7568
rect 167638 7556 167644 7568
rect 167696 7556 167702 7608
rect 204254 7556 204260 7608
rect 204312 7596 204318 7608
rect 546678 7596 546684 7608
rect 204312 7568 546684 7596
rect 204312 7556 204318 7568
rect 546678 7556 546684 7568
rect 546736 7556 546742 7608
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 153838 6848 153844 6860
rect 3476 6820 153844 6848
rect 3476 6808 3482 6820
rect 153838 6808 153844 6820
rect 153896 6808 153902 6860
rect 193122 6264 193128 6316
rect 193180 6304 193186 6316
rect 383562 6304 383568 6316
rect 193180 6276 383568 6304
rect 193180 6264 193186 6276
rect 383562 6264 383568 6276
rect 383620 6264 383626 6316
rect 193030 6196 193036 6248
rect 193088 6236 193094 6248
rect 387150 6236 387156 6248
rect 193088 6208 387156 6236
rect 193088 6196 193094 6208
rect 387150 6196 387156 6208
rect 387208 6196 387214 6248
rect 199838 6128 199844 6180
rect 199896 6168 199902 6180
rect 475746 6168 475752 6180
rect 199896 6140 475752 6168
rect 199896 6128 199902 6140
rect 475746 6128 475752 6140
rect 475804 6128 475810 6180
rect 176286 5516 176292 5568
rect 176344 5556 176350 5568
rect 177850 5556 177856 5568
rect 176344 5528 177856 5556
rect 176344 5516 176350 5528
rect 177850 5516 177856 5528
rect 177908 5516 177914 5568
rect 5258 4768 5264 4820
rect 5316 4808 5322 4820
rect 46198 4808 46204 4820
rect 5316 4780 46204 4808
rect 5316 4768 5322 4780
rect 46198 4768 46204 4780
rect 46256 4768 46262 4820
rect 64322 4768 64328 4820
rect 64380 4808 64386 4820
rect 167914 4808 167920 4820
rect 64380 4780 167920 4808
rect 64380 4768 64386 4780
rect 167914 4768 167920 4780
rect 167972 4768 167978 4820
rect 209682 4088 209688 4140
rect 209740 4128 209746 4140
rect 210970 4128 210976 4140
rect 209740 4100 210976 4128
rect 209740 4088 209746 4100
rect 210970 4088 210976 4100
rect 211028 4088 211034 4140
rect 232498 4088 232504 4140
rect 232556 4128 232562 4140
rect 246390 4128 246396 4140
rect 232556 4100 246396 4128
rect 232556 4088 232562 4100
rect 246390 4088 246396 4100
rect 246448 4088 246454 4140
rect 250438 4088 250444 4140
rect 250496 4128 250502 4140
rect 264146 4128 264152 4140
rect 250496 4100 264152 4128
rect 250496 4088 250502 4100
rect 264146 4088 264152 4100
rect 264204 4088 264210 4140
rect 266998 4088 267004 4140
rect 267056 4128 267062 4140
rect 267056 4100 277394 4128
rect 267056 4088 267062 4100
rect 13538 4020 13544 4072
rect 13596 4060 13602 4072
rect 17218 4060 17224 4072
rect 13596 4032 17224 4060
rect 13596 4020 13602 4032
rect 17218 4020 17224 4032
rect 17276 4020 17282 4072
rect 235258 4020 235264 4072
rect 235316 4060 235322 4072
rect 235316 4032 238754 4060
rect 235316 4020 235322 4032
rect 211798 3952 211804 4004
rect 211856 3992 211862 4004
rect 221550 3992 221556 4004
rect 211856 3964 221556 3992
rect 211856 3952 211862 3964
rect 221550 3952 221556 3964
rect 221608 3952 221614 4004
rect 238726 3992 238754 4032
rect 242802 4020 242808 4072
rect 242860 4060 242866 4072
rect 267642 4060 267648 4072
rect 242860 4032 253244 4060
rect 242860 4020 242866 4032
rect 249978 3992 249984 4004
rect 238726 3964 249984 3992
rect 249978 3952 249984 3964
rect 250036 3952 250042 4004
rect 180150 3884 180156 3936
rect 180208 3924 180214 3936
rect 181438 3924 181444 3936
rect 180208 3896 181444 3924
rect 180208 3884 180214 3896
rect 181438 3884 181444 3896
rect 181496 3884 181502 3936
rect 184290 3884 184296 3936
rect 184348 3924 184354 3936
rect 194410 3924 194416 3936
rect 184348 3896 194416 3924
rect 184348 3884 184354 3896
rect 194410 3884 194416 3896
rect 194468 3884 194474 3936
rect 213178 3884 213184 3936
rect 213236 3924 213242 3936
rect 225138 3924 225144 3936
rect 213236 3896 225144 3924
rect 213236 3884 213242 3896
rect 225138 3884 225144 3896
rect 225196 3884 225202 3936
rect 228358 3884 228364 3936
rect 228416 3924 228422 3936
rect 235810 3924 235816 3936
rect 228416 3896 235816 3924
rect 228416 3884 228422 3896
rect 235810 3884 235816 3896
rect 235868 3884 235874 3936
rect 243630 3884 243636 3936
rect 243688 3924 243694 3936
rect 253106 3924 253112 3936
rect 243688 3896 253112 3924
rect 243688 3884 243694 3896
rect 253106 3884 253112 3896
rect 253164 3884 253170 3936
rect 253216 3924 253244 4032
rect 258046 4032 267648 4060
rect 253290 3952 253296 4004
rect 253348 3992 253354 4004
rect 258046 3992 258074 4032
rect 267642 4020 267648 4032
rect 267700 4020 267706 4072
rect 253348 3964 258074 3992
rect 253348 3952 253354 3964
rect 265342 3952 265348 4004
rect 265400 3992 265406 4004
rect 274634 3992 274640 4004
rect 265400 3964 274640 3992
rect 265400 3952 265406 3964
rect 274634 3952 274640 3964
rect 274692 3952 274698 4004
rect 277366 3992 277394 4100
rect 302878 4088 302884 4140
rect 302936 4128 302942 4140
rect 306742 4128 306748 4140
rect 302936 4100 306748 4128
rect 302936 4088 302942 4100
rect 306742 4088 306748 4100
rect 306800 4088 306806 4140
rect 307018 4088 307024 4140
rect 307076 4128 307082 4140
rect 322106 4128 322112 4140
rect 307076 4100 322112 4128
rect 307076 4088 307082 4100
rect 322106 4088 322112 4100
rect 322164 4088 322170 4140
rect 323578 4088 323584 4140
rect 323636 4128 323642 4140
rect 327534 4128 327540 4140
rect 323636 4100 327540 4128
rect 323636 4088 323642 4100
rect 327534 4088 327540 4100
rect 327592 4088 327598 4140
rect 331582 4128 331588 4140
rect 327736 4100 331588 4128
rect 284938 4020 284944 4072
rect 284996 4060 285002 4072
rect 303154 4060 303160 4072
rect 284996 4032 303160 4060
rect 284996 4020 285002 4032
rect 303154 4020 303160 4032
rect 303212 4020 303218 4072
rect 315298 4020 315304 4072
rect 315356 4060 315362 4072
rect 316218 4060 316224 4072
rect 315356 4032 316224 4060
rect 315356 4020 315362 4032
rect 316218 4020 316224 4032
rect 316276 4020 316282 4072
rect 319438 4020 319444 4072
rect 319496 4060 319502 4072
rect 319496 4032 320956 4060
rect 319496 4020 319502 4032
rect 288986 3992 288992 4004
rect 277366 3964 288992 3992
rect 288986 3952 288992 3964
rect 289044 3952 289050 4004
rect 311158 3952 311164 4004
rect 311216 3992 311222 4004
rect 320818 3992 320824 4004
rect 311216 3964 320824 3992
rect 311216 3952 311222 3964
rect 320818 3952 320824 3964
rect 320876 3952 320882 4004
rect 320928 3992 320956 4032
rect 321094 4020 321100 4072
rect 321152 4060 321158 4072
rect 327736 4060 327764 4100
rect 331582 4088 331588 4100
rect 331640 4088 331646 4140
rect 363598 4088 363604 4140
rect 363656 4128 363662 4140
rect 367002 4128 367008 4140
rect 363656 4100 367008 4128
rect 363656 4088 363662 4100
rect 367002 4088 367008 4100
rect 367060 4088 367066 4140
rect 429838 4088 429844 4140
rect 429896 4128 429902 4140
rect 432046 4128 432052 4140
rect 429896 4100 432052 4128
rect 429896 4088 429902 4100
rect 432046 4088 432052 4100
rect 432104 4088 432110 4140
rect 489178 4088 489184 4140
rect 489236 4128 489242 4140
rect 489914 4128 489920 4140
rect 489236 4100 489920 4128
rect 489236 4088 489242 4100
rect 489914 4088 489920 4100
rect 489972 4088 489978 4140
rect 547138 4088 547144 4140
rect 547196 4128 547202 4140
rect 547874 4128 547880 4140
rect 547196 4100 547880 4128
rect 547196 4088 547202 4100
rect 547874 4088 547880 4100
rect 547932 4088 547938 4140
rect 321152 4032 327764 4060
rect 321152 4020 321158 4032
rect 327810 4020 327816 4072
rect 327868 4060 327874 4072
rect 329282 4060 329288 4072
rect 327868 4032 329288 4060
rect 327868 4020 327874 4032
rect 329282 4020 329288 4032
rect 329340 4020 329346 4072
rect 337378 4020 337384 4072
rect 337436 4060 337442 4072
rect 359918 4060 359924 4072
rect 337436 4032 359924 4060
rect 337436 4020 337442 4032
rect 359918 4020 359924 4032
rect 359976 4020 359982 4072
rect 349154 3992 349160 4004
rect 320928 3964 349160 3992
rect 349154 3952 349160 3964
rect 349212 3952 349218 4004
rect 268838 3924 268844 3936
rect 253216 3896 268844 3924
rect 268838 3884 268844 3896
rect 268896 3884 268902 3936
rect 269758 3884 269764 3936
rect 269816 3924 269822 3936
rect 292574 3924 292580 3936
rect 269816 3896 292580 3924
rect 269816 3884 269822 3896
rect 292574 3884 292580 3896
rect 292632 3884 292638 3936
rect 309778 3884 309784 3936
rect 309836 3924 309842 3936
rect 346946 3924 346952 3936
rect 309836 3896 346952 3924
rect 309836 3884 309842 3896
rect 346946 3884 346952 3896
rect 347004 3884 347010 3936
rect 381630 3884 381636 3936
rect 381688 3924 381694 3936
rect 384758 3924 384764 3936
rect 381688 3896 384764 3924
rect 381688 3884 381694 3896
rect 384758 3884 384764 3896
rect 384816 3884 384822 3936
rect 180058 3816 180064 3868
rect 180116 3856 180122 3868
rect 189718 3856 189724 3868
rect 180116 3828 189724 3856
rect 180116 3816 180122 3828
rect 189718 3816 189724 3828
rect 189776 3816 189782 3868
rect 214558 3816 214564 3868
rect 214616 3856 214622 3868
rect 232222 3856 232228 3868
rect 214616 3828 232228 3856
rect 214616 3816 214622 3828
rect 232222 3816 232228 3828
rect 232280 3816 232286 3868
rect 243538 3816 243544 3868
rect 243596 3856 243602 3868
rect 272426 3856 272432 3868
rect 243596 3828 272432 3856
rect 243596 3816 243602 3828
rect 272426 3816 272432 3828
rect 272484 3816 272490 3868
rect 301498 3816 301504 3868
rect 301556 3856 301562 3868
rect 324314 3856 324320 3868
rect 301556 3828 324320 3856
rect 301556 3816 301562 3828
rect 324314 3816 324320 3828
rect 324372 3816 324378 3868
rect 327718 3816 327724 3868
rect 327776 3856 327782 3868
rect 329190 3856 329196 3868
rect 327776 3828 329196 3856
rect 327776 3816 327782 3828
rect 329190 3816 329196 3828
rect 329248 3816 329254 3868
rect 329282 3816 329288 3868
rect 329340 3856 329346 3868
rect 368198 3856 368204 3868
rect 329340 3828 368204 3856
rect 329340 3816 329346 3828
rect 368198 3816 368204 3828
rect 368256 3816 368262 3868
rect 384298 3816 384304 3868
rect 384356 3856 384362 3868
rect 398834 3856 398840 3868
rect 384356 3828 398840 3856
rect 384356 3816 384362 3828
rect 398834 3816 398840 3828
rect 398892 3816 398898 3868
rect 186958 3748 186964 3800
rect 187016 3788 187022 3800
rect 203886 3788 203892 3800
rect 187016 3760 203892 3788
rect 187016 3748 187022 3760
rect 203886 3748 203892 3760
rect 203944 3748 203950 3800
rect 217318 3748 217324 3800
rect 217376 3788 217382 3800
rect 239306 3788 239312 3800
rect 217376 3760 239312 3788
rect 217376 3748 217382 3760
rect 239306 3748 239312 3760
rect 239364 3748 239370 3800
rect 243722 3748 243728 3800
rect 243780 3788 243786 3800
rect 286594 3788 286600 3800
rect 243780 3760 286600 3788
rect 243780 3748 243786 3760
rect 286594 3748 286600 3760
rect 286652 3748 286658 3800
rect 313918 3748 313924 3800
rect 313976 3788 313982 3800
rect 403618 3788 403624 3800
rect 313976 3760 403624 3788
rect 313976 3748 313982 3760
rect 403618 3748 403624 3760
rect 403676 3748 403682 3800
rect 520734 3788 520740 3800
rect 509206 3760 520740 3788
rect 123478 3680 123484 3732
rect 123536 3720 123542 3732
rect 133138 3720 133144 3732
rect 123536 3692 133144 3720
rect 123536 3680 123542 3692
rect 133138 3680 133144 3692
rect 133196 3680 133202 3732
rect 135254 3680 135260 3732
rect 135312 3720 135318 3732
rect 136450 3720 136456 3732
rect 135312 3692 136456 3720
rect 135312 3680 135318 3692
rect 136450 3680 136456 3692
rect 136508 3680 136514 3732
rect 186038 3680 186044 3732
rect 186096 3720 186102 3732
rect 291378 3720 291384 3732
rect 186096 3692 291384 3720
rect 186096 3680 186102 3692
rect 291378 3680 291384 3692
rect 291436 3680 291442 3732
rect 305638 3680 305644 3732
rect 305696 3720 305702 3732
rect 311434 3720 311440 3732
rect 305696 3692 311440 3720
rect 305696 3680 305702 3692
rect 311434 3680 311440 3692
rect 311492 3680 311498 3732
rect 314010 3680 314016 3732
rect 314068 3720 314074 3732
rect 317322 3720 317328 3732
rect 314068 3692 317328 3720
rect 314068 3680 314074 3692
rect 317322 3680 317328 3692
rect 317380 3680 317386 3732
rect 320818 3680 320824 3732
rect 320876 3720 320882 3732
rect 364610 3720 364616 3732
rect 320876 3692 364616 3720
rect 320876 3680 320882 3692
rect 364610 3680 364616 3692
rect 364668 3680 364674 3732
rect 381538 3680 381544 3732
rect 381596 3720 381602 3732
rect 509206 3720 509234 3760
rect 520734 3748 520740 3760
rect 520792 3748 520798 3800
rect 381596 3692 509234 3720
rect 381596 3680 381602 3692
rect 12342 3612 12348 3664
rect 12400 3652 12406 3664
rect 15838 3652 15844 3664
rect 12400 3624 15844 3652
rect 12400 3612 12406 3624
rect 15838 3612 15844 3624
rect 15896 3612 15902 3664
rect 37182 3612 37188 3664
rect 37240 3652 37246 3664
rect 68278 3652 68284 3664
rect 37240 3624 68284 3652
rect 37240 3612 37246 3624
rect 68278 3612 68284 3624
rect 68336 3612 68342 3664
rect 68388 3624 74534 3652
rect 2866 3544 2872 3596
rect 2924 3584 2930 3596
rect 13078 3584 13084 3596
rect 2924 3556 13084 3584
rect 2924 3544 2930 3556
rect 13078 3544 13084 3556
rect 13136 3544 13142 3596
rect 60734 3544 60740 3596
rect 60792 3584 60798 3596
rect 61654 3584 61660 3596
rect 60792 3556 61660 3584
rect 60792 3544 60798 3556
rect 61654 3544 61660 3556
rect 61712 3544 61718 3596
rect 67910 3544 67916 3596
rect 67968 3584 67974 3596
rect 68388 3584 68416 3624
rect 67968 3556 68416 3584
rect 67968 3544 67974 3556
rect 69106 3544 69112 3596
rect 69164 3584 69170 3596
rect 71038 3584 71044 3596
rect 69164 3556 71044 3584
rect 69164 3544 69170 3556
rect 71038 3544 71044 3556
rect 71096 3544 71102 3596
rect 74506 3584 74534 3624
rect 77386 3612 77392 3664
rect 77444 3652 77450 3664
rect 80698 3652 80704 3664
rect 77444 3624 80704 3652
rect 77444 3612 77450 3624
rect 80698 3612 80704 3624
rect 80756 3612 80762 3664
rect 86862 3612 86868 3664
rect 86920 3652 86926 3664
rect 88978 3652 88984 3664
rect 86920 3624 88984 3652
rect 86920 3612 86926 3624
rect 88978 3612 88984 3624
rect 89036 3612 89042 3664
rect 109310 3612 109316 3664
rect 109368 3652 109374 3664
rect 112438 3652 112444 3664
rect 109368 3624 112444 3652
rect 109368 3612 109374 3624
rect 112438 3612 112444 3624
rect 112496 3612 112502 3664
rect 118786 3612 118792 3664
rect 118844 3652 118850 3664
rect 120718 3652 120724 3664
rect 118844 3624 120724 3652
rect 118844 3612 118850 3624
rect 120718 3612 120724 3624
rect 120776 3612 120782 3664
rect 121086 3612 121092 3664
rect 121144 3652 121150 3664
rect 122098 3652 122104 3664
rect 121144 3624 122104 3652
rect 121144 3612 121150 3624
rect 122098 3612 122104 3624
rect 122156 3612 122162 3664
rect 124674 3612 124680 3664
rect 124732 3652 124738 3664
rect 124732 3624 128400 3652
rect 124732 3612 124738 3624
rect 123386 3584 123392 3596
rect 74506 3556 123392 3584
rect 123386 3544 123392 3556
rect 123444 3544 123450 3596
rect 126974 3544 126980 3596
rect 127032 3584 127038 3596
rect 128170 3584 128176 3596
rect 127032 3556 128176 3584
rect 127032 3544 127038 3556
rect 128170 3544 128176 3556
rect 128228 3544 128234 3596
rect 128372 3584 128400 3624
rect 129366 3612 129372 3664
rect 129424 3652 129430 3664
rect 160186 3652 160192 3664
rect 129424 3624 160192 3652
rect 129424 3612 129430 3624
rect 160186 3612 160192 3624
rect 160244 3612 160250 3664
rect 170766 3612 170772 3664
rect 170824 3652 170830 3664
rect 174630 3652 174636 3664
rect 170824 3624 174636 3652
rect 170824 3612 170830 3624
rect 174630 3612 174636 3624
rect 174688 3612 174694 3664
rect 179230 3612 179236 3664
rect 179288 3652 179294 3664
rect 200298 3652 200304 3664
rect 179288 3624 200304 3652
rect 179288 3612 179294 3624
rect 200298 3612 200304 3624
rect 200356 3612 200362 3664
rect 215938 3612 215944 3664
rect 215996 3652 216002 3664
rect 242894 3652 242900 3664
rect 215996 3624 242900 3652
rect 215996 3612 216002 3624
rect 242894 3612 242900 3624
rect 242952 3612 242958 3664
rect 251818 3612 251824 3664
rect 251876 3652 251882 3664
rect 254670 3652 254676 3664
rect 251876 3624 254676 3652
rect 251876 3612 251882 3624
rect 254670 3612 254676 3624
rect 254728 3612 254734 3664
rect 254762 3612 254768 3664
rect 254820 3652 254826 3664
rect 373994 3652 374000 3664
rect 254820 3624 374000 3652
rect 254820 3612 254826 3624
rect 373994 3612 374000 3624
rect 374052 3612 374058 3664
rect 387058 3612 387064 3664
rect 387116 3652 387122 3664
rect 573910 3652 573916 3664
rect 387116 3624 573916 3652
rect 387116 3612 387122 3624
rect 573910 3612 573916 3624
rect 573968 3612 573974 3664
rect 162118 3584 162124 3596
rect 128372 3556 162124 3584
rect 162118 3544 162124 3556
rect 162176 3544 162182 3596
rect 169570 3544 169576 3596
rect 169628 3584 169634 3596
rect 174538 3584 174544 3596
rect 169628 3556 174544 3584
rect 169628 3544 169634 3556
rect 174538 3544 174544 3556
rect 174596 3544 174602 3596
rect 179322 3544 179328 3596
rect 179380 3584 179386 3596
rect 184934 3584 184940 3596
rect 179380 3556 184940 3584
rect 179380 3544 179386 3556
rect 184934 3544 184940 3556
rect 184992 3544 184998 3596
rect 186222 3544 186228 3596
rect 186280 3584 186286 3596
rect 294874 3584 294880 3596
rect 186280 3556 294880 3584
rect 186280 3544 186286 3556
rect 294874 3544 294880 3556
rect 294932 3544 294938 3596
rect 295978 3544 295984 3596
rect 296036 3584 296042 3596
rect 299474 3584 299480 3596
rect 296036 3556 299480 3584
rect 296036 3544 296042 3556
rect 299474 3544 299480 3556
rect 299532 3544 299538 3596
rect 299566 3544 299572 3596
rect 299624 3584 299630 3596
rect 300762 3584 300768 3596
rect 299624 3556 300768 3584
rect 299624 3544 299630 3556
rect 300762 3544 300768 3556
rect 300820 3544 300826 3596
rect 305730 3544 305736 3596
rect 305788 3584 305794 3596
rect 307662 3584 307668 3596
rect 305788 3556 307668 3584
rect 305788 3544 305794 3556
rect 307662 3544 307668 3556
rect 307720 3544 307726 3596
rect 307846 3544 307852 3596
rect 307904 3584 307910 3596
rect 309042 3584 309048 3596
rect 307904 3556 309048 3584
rect 307904 3544 307910 3556
rect 309042 3544 309048 3556
rect 309100 3544 309106 3596
rect 316678 3544 316684 3596
rect 316736 3584 316742 3596
rect 321094 3584 321100 3596
rect 316736 3556 321100 3584
rect 316736 3544 316742 3556
rect 321094 3544 321100 3556
rect 321152 3544 321158 3596
rect 321462 3544 321468 3596
rect 321520 3584 321526 3596
rect 510062 3584 510068 3596
rect 321520 3556 510068 3584
rect 321520 3544 321526 3556
rect 510062 3544 510068 3556
rect 510120 3544 510126 3596
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 14458 3516 14464 3528
rect 1728 3488 14464 3516
rect 1728 3476 1734 3488
rect 14458 3476 14464 3488
rect 14516 3476 14522 3528
rect 17034 3476 17040 3528
rect 17092 3516 17098 3528
rect 18598 3516 18604 3528
rect 17092 3488 18604 3516
rect 17092 3476 17098 3488
rect 18598 3476 18604 3488
rect 18656 3476 18662 3528
rect 23014 3476 23020 3528
rect 23072 3516 23078 3528
rect 24118 3516 24124 3528
rect 23072 3488 24124 3516
rect 23072 3476 23078 3488
rect 24118 3476 24124 3488
rect 24176 3476 24182 3528
rect 38378 3476 38384 3528
rect 38436 3516 38442 3528
rect 39298 3516 39304 3528
rect 38436 3488 39304 3516
rect 38436 3476 38442 3488
rect 39298 3476 39304 3488
rect 39356 3476 39362 3528
rect 41874 3476 41880 3528
rect 41932 3516 41938 3528
rect 43438 3516 43444 3528
rect 41932 3488 43444 3516
rect 41932 3476 41938 3488
rect 43438 3476 43444 3488
rect 43496 3476 43502 3528
rect 46658 3476 46664 3528
rect 46716 3516 46722 3528
rect 46716 3488 158116 3516
rect 46716 3476 46722 3488
rect 6454 3408 6460 3460
rect 6512 3448 6518 3460
rect 157978 3448 157984 3460
rect 6512 3420 157984 3448
rect 6512 3408 6518 3420
rect 157978 3408 157984 3420
rect 158036 3408 158042 3460
rect 158088 3448 158116 3488
rect 160094 3476 160100 3528
rect 160152 3516 160158 3528
rect 161290 3516 161296 3528
rect 160152 3488 161296 3516
rect 160152 3476 160158 3488
rect 161290 3476 161296 3488
rect 161348 3476 161354 3528
rect 168374 3476 168380 3528
rect 168432 3516 168438 3528
rect 176378 3516 176384 3528
rect 168432 3488 176384 3516
rect 168432 3476 168438 3488
rect 176378 3476 176384 3488
rect 176436 3476 176442 3528
rect 182082 3476 182088 3528
rect 182140 3516 182146 3528
rect 183738 3516 183744 3528
rect 182140 3488 183744 3516
rect 182140 3476 182146 3488
rect 183738 3476 183744 3488
rect 183796 3476 183802 3528
rect 190426 3488 191052 3516
rect 160738 3448 160744 3460
rect 158088 3420 160744 3448
rect 160738 3408 160744 3420
rect 160796 3408 160802 3460
rect 166074 3408 166080 3460
rect 166132 3448 166138 3460
rect 173158 3448 173164 3460
rect 166132 3420 173164 3448
rect 166132 3408 166138 3420
rect 173158 3408 173164 3420
rect 173216 3408 173222 3460
rect 181530 3408 181536 3460
rect 181588 3448 181594 3460
rect 190426 3448 190454 3488
rect 181588 3420 190454 3448
rect 191024 3448 191052 3488
rect 191098 3476 191104 3528
rect 191156 3516 191162 3528
rect 192018 3516 192024 3528
rect 191156 3488 192024 3516
rect 191156 3476 191162 3488
rect 192018 3476 192024 3488
rect 192076 3476 192082 3528
rect 193858 3476 193864 3528
rect 193916 3516 193922 3528
rect 195606 3516 195612 3528
rect 193916 3488 195612 3516
rect 193916 3476 193922 3488
rect 195606 3476 195612 3488
rect 195664 3476 195670 3528
rect 196618 3476 196624 3528
rect 196676 3516 196682 3528
rect 199102 3516 199108 3528
rect 196676 3488 199108 3516
rect 196676 3476 196682 3488
rect 199102 3476 199108 3488
rect 199160 3476 199166 3528
rect 199930 3476 199936 3528
rect 199988 3516 199994 3528
rect 468294 3516 468300 3528
rect 199988 3488 468300 3516
rect 199988 3476 199994 3488
rect 468294 3476 468300 3488
rect 468352 3476 468358 3528
rect 468478 3476 468484 3528
rect 468536 3516 468542 3528
rect 469858 3516 469864 3528
rect 468536 3488 469864 3516
rect 468536 3476 468542 3488
rect 469858 3476 469864 3488
rect 469916 3476 469922 3528
rect 472618 3476 472624 3528
rect 472676 3516 472682 3528
rect 473446 3516 473452 3528
rect 472676 3488 473452 3516
rect 472676 3476 472682 3488
rect 473446 3476 473452 3488
rect 473504 3476 473510 3528
rect 498194 3476 498200 3528
rect 498252 3516 498258 3528
rect 499022 3516 499028 3528
rect 498252 3488 499028 3516
rect 498252 3476 498258 3488
rect 499022 3476 499028 3488
rect 499080 3476 499086 3528
rect 520918 3476 520924 3528
rect 520976 3516 520982 3528
rect 521838 3516 521844 3528
rect 520976 3488 521844 3516
rect 520976 3476 520982 3488
rect 521838 3476 521844 3488
rect 521896 3476 521902 3528
rect 522298 3476 522304 3528
rect 522356 3516 522362 3528
rect 523034 3516 523040 3528
rect 522356 3488 523040 3516
rect 522356 3476 522362 3488
rect 523034 3476 523040 3488
rect 523092 3476 523098 3528
rect 564434 3476 564440 3528
rect 564492 3516 564498 3528
rect 565262 3516 565268 3528
rect 564492 3488 565268 3516
rect 564492 3476 564498 3488
rect 565262 3476 565268 3488
rect 565320 3476 565326 3528
rect 193214 3448 193220 3460
rect 191024 3420 193220 3448
rect 181588 3408 181594 3420
rect 193214 3408 193220 3420
rect 193272 3408 193278 3460
rect 200022 3408 200028 3460
rect 200080 3448 200086 3460
rect 472250 3448 472256 3460
rect 200080 3420 472256 3448
rect 200080 3408 200086 3420
rect 472250 3408 472256 3420
rect 472308 3408 472314 3460
rect 78582 3340 78588 3392
rect 78640 3380 78646 3392
rect 79318 3380 79324 3392
rect 78640 3352 79324 3380
rect 78640 3340 78646 3352
rect 79318 3340 79324 3352
rect 79376 3340 79382 3392
rect 110414 3340 110420 3392
rect 110472 3380 110478 3392
rect 111610 3380 111616 3392
rect 110472 3352 111616 3380
rect 110472 3340 110478 3352
rect 111610 3340 111616 3352
rect 111668 3340 111674 3392
rect 114002 3340 114008 3392
rect 114060 3380 114066 3392
rect 115198 3380 115204 3392
rect 114060 3352 115204 3380
rect 114060 3340 114066 3352
rect 115198 3340 115204 3352
rect 115256 3340 115262 3392
rect 118694 3340 118700 3392
rect 118752 3380 118758 3392
rect 119890 3380 119896 3392
rect 118752 3352 119896 3380
rect 118752 3340 118758 3352
rect 119890 3340 119896 3352
rect 119948 3340 119954 3392
rect 126974 3340 126980 3392
rect 127032 3380 127038 3392
rect 128998 3380 129004 3392
rect 127032 3352 129004 3380
rect 127032 3340 127038 3352
rect 128998 3340 129004 3352
rect 129056 3340 129062 3392
rect 149514 3340 149520 3392
rect 149572 3380 149578 3392
rect 151078 3380 151084 3392
rect 149572 3352 151084 3380
rect 149572 3340 149578 3352
rect 151078 3340 151084 3352
rect 151136 3340 151142 3392
rect 182818 3340 182824 3392
rect 182876 3380 182882 3392
rect 196802 3380 196808 3392
rect 182876 3352 196808 3380
rect 182876 3340 182882 3352
rect 196802 3340 196808 3352
rect 196860 3340 196866 3392
rect 239398 3340 239404 3392
rect 239456 3380 239462 3392
rect 253474 3380 253480 3392
rect 239456 3352 253480 3380
rect 239456 3340 239462 3352
rect 253474 3340 253480 3352
rect 253532 3340 253538 3392
rect 253566 3340 253572 3392
rect 253624 3380 253630 3392
rect 258258 3380 258264 3392
rect 253624 3352 258264 3380
rect 253624 3340 253630 3352
rect 258258 3340 258264 3352
rect 258316 3340 258322 3392
rect 264238 3340 264244 3392
rect 264296 3380 264302 3392
rect 271230 3380 271236 3392
rect 264296 3352 271236 3380
rect 264296 3340 264302 3352
rect 271230 3340 271236 3352
rect 271288 3340 271294 3392
rect 275278 3340 275284 3392
rect 275336 3380 275342 3392
rect 278314 3380 278320 3392
rect 275336 3352 278320 3380
rect 275336 3340 275342 3352
rect 278314 3340 278320 3352
rect 278372 3340 278378 3392
rect 307662 3340 307668 3392
rect 307720 3380 307726 3392
rect 315022 3380 315028 3392
rect 307720 3352 315028 3380
rect 307720 3340 307726 3352
rect 315022 3340 315028 3352
rect 315080 3340 315086 3392
rect 324406 3340 324412 3392
rect 324464 3380 324470 3392
rect 325602 3380 325608 3392
rect 324464 3352 325608 3380
rect 324464 3340 324470 3352
rect 325602 3340 325608 3352
rect 325660 3340 325666 3392
rect 327534 3340 327540 3392
rect 327592 3380 327598 3392
rect 335078 3380 335084 3392
rect 327592 3352 335084 3380
rect 327592 3340 327598 3352
rect 335078 3340 335084 3352
rect 335136 3340 335142 3392
rect 340966 3340 340972 3392
rect 341024 3380 341030 3392
rect 342162 3380 342168 3392
rect 341024 3352 342168 3380
rect 341024 3340 341030 3352
rect 342162 3340 342168 3352
rect 342220 3340 342226 3392
rect 349246 3340 349252 3392
rect 349304 3380 349310 3392
rect 350442 3380 350448 3392
rect 349304 3352 350448 3380
rect 349304 3340 349310 3352
rect 350442 3340 350448 3352
rect 350500 3340 350506 3392
rect 359458 3340 359464 3392
rect 359516 3380 359522 3392
rect 363506 3380 363512 3392
rect 359516 3352 363512 3380
rect 359516 3340 359522 3352
rect 363506 3340 363512 3352
rect 363564 3340 363570 3392
rect 374086 3340 374092 3392
rect 374144 3380 374150 3392
rect 375282 3380 375288 3392
rect 374144 3352 375288 3380
rect 374144 3340 374150 3352
rect 375282 3340 375288 3352
rect 375340 3340 375346 3392
rect 376110 3340 376116 3392
rect 376168 3380 376174 3392
rect 381170 3380 381176 3392
rect 376168 3352 381176 3380
rect 376168 3340 376174 3352
rect 381170 3340 381176 3352
rect 381228 3340 381234 3392
rect 390554 3340 390560 3392
rect 390612 3380 390618 3392
rect 391842 3380 391848 3392
rect 390612 3352 391848 3380
rect 390612 3340 390618 3352
rect 391842 3340 391848 3352
rect 391900 3340 391906 3392
rect 398926 3340 398932 3392
rect 398984 3380 398990 3392
rect 400122 3380 400128 3392
rect 398984 3352 400128 3380
rect 398984 3340 398990 3352
rect 400122 3340 400128 3352
rect 400180 3340 400186 3392
rect 407206 3340 407212 3392
rect 407264 3380 407270 3392
rect 408402 3380 408408 3392
rect 407264 3352 408408 3380
rect 407264 3340 407270 3352
rect 408402 3340 408408 3352
rect 408460 3340 408466 3392
rect 423766 3340 423772 3392
rect 423824 3380 423830 3392
rect 424962 3380 424968 3392
rect 423824 3352 424968 3380
rect 423824 3340 423830 3352
rect 424962 3340 424968 3352
rect 425020 3340 425026 3392
rect 570598 3340 570604 3392
rect 570656 3380 570662 3392
rect 577406 3380 577412 3392
rect 570656 3352 577412 3380
rect 570656 3340 570662 3352
rect 577406 3340 577412 3352
rect 577464 3340 577470 3392
rect 4062 3272 4068 3324
rect 4120 3312 4126 3324
rect 4798 3312 4804 3324
rect 4120 3284 4804 3312
rect 4120 3272 4126 3284
rect 4798 3272 4804 3284
rect 4856 3272 4862 3324
rect 24210 3272 24216 3324
rect 24268 3312 24274 3324
rect 25498 3312 25504 3324
rect 24268 3284 25504 3312
rect 24268 3272 24274 3284
rect 25498 3272 25504 3284
rect 25556 3272 25562 3324
rect 93946 3272 93952 3324
rect 94004 3312 94010 3324
rect 95878 3312 95884 3324
rect 94004 3284 95884 3312
rect 94004 3272 94010 3284
rect 95878 3272 95884 3284
rect 95936 3272 95942 3324
rect 162486 3272 162492 3324
rect 162544 3312 162550 3324
rect 166258 3312 166264 3324
rect 162544 3284 166264 3312
rect 162544 3272 162550 3284
rect 166258 3272 166264 3284
rect 166316 3272 166322 3324
rect 246298 3272 246304 3324
rect 246356 3312 246362 3324
rect 257062 3312 257068 3324
rect 246356 3284 257068 3312
rect 246356 3272 246362 3284
rect 257062 3272 257068 3284
rect 257120 3272 257126 3324
rect 265618 3272 265624 3324
rect 265676 3312 265682 3324
rect 266538 3312 266544 3324
rect 265676 3284 266544 3312
rect 265676 3272 265682 3284
rect 266538 3272 266544 3284
rect 266596 3272 266602 3324
rect 271138 3272 271144 3324
rect 271196 3312 271202 3324
rect 274818 3312 274824 3324
rect 271196 3284 274824 3312
rect 271196 3272 271202 3284
rect 274818 3272 274824 3284
rect 274876 3272 274882 3324
rect 571978 3272 571984 3324
rect 572036 3312 572042 3324
rect 572714 3312 572720 3324
rect 572036 3284 572720 3312
rect 572036 3272 572042 3284
rect 572714 3272 572720 3284
rect 572772 3272 572778 3324
rect 27706 3204 27712 3256
rect 27764 3244 27770 3256
rect 31018 3244 31024 3256
rect 27764 3216 31024 3244
rect 27764 3204 27770 3216
rect 31018 3204 31024 3216
rect 31076 3204 31082 3256
rect 31294 3204 31300 3256
rect 31352 3244 31358 3256
rect 36538 3244 36544 3256
rect 31352 3216 36544 3244
rect 31352 3204 31358 3216
rect 36538 3204 36544 3216
rect 36596 3204 36602 3256
rect 115198 3204 115204 3256
rect 115256 3244 115262 3256
rect 117958 3244 117964 3256
rect 115256 3216 117964 3244
rect 115256 3204 115262 3216
rect 117958 3204 117964 3216
rect 118016 3204 118022 3256
rect 160094 3204 160100 3256
rect 160152 3244 160158 3256
rect 161474 3244 161480 3256
rect 160152 3216 161480 3244
rect 160152 3204 160158 3216
rect 161474 3204 161480 3216
rect 161532 3204 161538 3256
rect 241238 3204 241244 3256
rect 241296 3244 241302 3256
rect 251174 3244 251180 3256
rect 241296 3216 251180 3244
rect 241296 3204 241302 3216
rect 251174 3204 251180 3216
rect 251232 3204 251238 3256
rect 253106 3204 253112 3256
rect 253164 3244 253170 3256
rect 253164 3216 254900 3244
rect 253164 3204 253170 3216
rect 249702 3136 249708 3188
rect 249760 3176 249766 3188
rect 254762 3176 254768 3188
rect 249760 3148 254768 3176
rect 249760 3136 249766 3148
rect 254762 3136 254768 3148
rect 254820 3136 254826 3188
rect 254872 3176 254900 3216
rect 309870 3204 309876 3256
rect 309928 3244 309934 3256
rect 313826 3244 313832 3256
rect 309928 3216 313832 3244
rect 309928 3204 309934 3216
rect 313826 3204 313832 3216
rect 313884 3204 313890 3256
rect 260650 3176 260656 3188
rect 254872 3148 260656 3176
rect 260650 3136 260656 3148
rect 260708 3136 260714 3188
rect 542998 3136 543004 3188
rect 543056 3176 543062 3188
rect 545482 3176 545488 3188
rect 543056 3148 545488 3176
rect 543056 3136 543062 3148
rect 545482 3136 545488 3148
rect 545540 3136 545546 3188
rect 552750 3136 552756 3188
rect 552808 3176 552814 3188
rect 556154 3176 556160 3188
rect 552808 3148 556160 3176
rect 552808 3136 552814 3148
rect 556154 3136 556160 3148
rect 556212 3136 556218 3188
rect 569218 3136 569224 3188
rect 569276 3176 569282 3188
rect 571518 3176 571524 3188
rect 569276 3148 571524 3176
rect 569276 3136 569282 3148
rect 571518 3136 571524 3148
rect 571576 3136 571582 3188
rect 189810 3068 189816 3120
rect 189868 3108 189874 3120
rect 190822 3108 190828 3120
rect 189868 3080 190828 3108
rect 189868 3068 189874 3080
rect 190822 3068 190828 3080
rect 190880 3068 190886 3120
rect 210418 3068 210424 3120
rect 210476 3108 210482 3120
rect 218054 3108 218060 3120
rect 210476 3080 218060 3108
rect 210476 3068 210482 3080
rect 218054 3068 218060 3080
rect 218112 3068 218118 3120
rect 287698 3068 287704 3120
rect 287756 3108 287762 3120
rect 290182 3108 290188 3120
rect 287756 3080 290188 3108
rect 287756 3068 287762 3080
rect 290182 3068 290188 3080
rect 290240 3068 290246 3120
rect 307110 3068 307116 3120
rect 307168 3108 307174 3120
rect 310238 3108 310244 3120
rect 307168 3080 310244 3108
rect 307168 3068 307174 3080
rect 310238 3068 310244 3080
rect 310296 3068 310302 3120
rect 471238 3068 471244 3120
rect 471296 3108 471302 3120
rect 474550 3108 474556 3120
rect 471296 3080 474556 3108
rect 471296 3068 471302 3080
rect 474550 3068 474556 3080
rect 474608 3068 474614 3120
rect 167178 3000 167184 3052
rect 167236 3040 167242 3052
rect 169018 3040 169024 3052
rect 167236 3012 169024 3040
rect 167236 3000 167242 3012
rect 169018 3000 169024 3012
rect 169076 3000 169082 3052
rect 184198 3000 184204 3052
rect 184256 3040 184262 3052
rect 186130 3040 186136 3052
rect 184256 3012 186136 3040
rect 184256 3000 184262 3012
rect 186130 3000 186136 3012
rect 186188 3000 186194 3052
rect 225598 3000 225604 3052
rect 225656 3040 225662 3052
rect 228726 3040 228732 3052
rect 225656 3012 228732 3040
rect 225656 3000 225662 3012
rect 228726 3000 228732 3012
rect 228784 3000 228790 3052
rect 278038 3000 278044 3052
rect 278096 3040 278102 3052
rect 281902 3040 281908 3052
rect 278096 3012 281908 3040
rect 278096 3000 278102 3012
rect 281902 3000 281908 3012
rect 281960 3000 281966 3052
rect 282178 3000 282184 3052
rect 282236 3040 282242 3052
rect 285398 3040 285404 3052
rect 282236 3012 285404 3040
rect 282236 3000 282242 3012
rect 285398 3000 285404 3012
rect 285456 3000 285462 3052
rect 289078 3000 289084 3052
rect 289136 3040 289142 3052
rect 296070 3040 296076 3052
rect 289136 3012 296076 3040
rect 289136 3000 289142 3012
rect 296070 3000 296076 3012
rect 296128 3000 296134 3052
rect 399478 3000 399484 3052
rect 399536 3040 399542 3052
rect 402514 3040 402520 3052
rect 399536 3012 402520 3040
rect 399536 3000 399542 3012
rect 402514 3000 402520 3012
rect 402572 3000 402578 3052
rect 422938 3000 422944 3052
rect 422996 3040 423002 3052
rect 423766 3040 423772 3052
rect 422996 3012 423772 3040
rect 422996 3000 423002 3012
rect 423766 3000 423772 3012
rect 423824 3000 423830 3052
rect 436738 3000 436744 3052
rect 436796 3040 436802 3052
rect 437934 3040 437940 3052
rect 436796 3012 437940 3040
rect 436796 3000 436802 3012
rect 437934 3000 437940 3012
rect 437992 3000 437998 3052
rect 514018 3000 514024 3052
rect 514076 3040 514082 3052
rect 515950 3040 515956 3052
rect 514076 3012 515956 3040
rect 514076 3000 514082 3012
rect 515950 3000 515956 3012
rect 516008 3000 516014 3052
rect 201402 2932 201408 2984
rect 201460 2972 201466 2984
rect 205082 2972 205088 2984
rect 201460 2944 205088 2972
rect 201460 2932 201466 2944
rect 205082 2932 205088 2944
rect 205140 2932 205146 2984
rect 240778 2932 240784 2984
rect 240836 2972 240842 2984
rect 247586 2972 247592 2984
rect 240836 2944 247592 2972
rect 240836 2932 240842 2944
rect 247586 2932 247592 2944
rect 247644 2932 247650 2984
rect 18230 2864 18236 2916
rect 18288 2904 18294 2916
rect 22738 2904 22744 2916
rect 18288 2876 22744 2904
rect 18288 2864 18294 2876
rect 22738 2864 22744 2876
rect 22796 2864 22802 2916
rect 242158 2864 242164 2916
rect 242216 2904 242222 2916
rect 244090 2904 244096 2916
rect 242216 2876 244096 2904
rect 242216 2864 242222 2876
rect 244090 2864 244096 2876
rect 244148 2864 244154 2916
rect 247678 2864 247684 2916
rect 247736 2904 247742 2916
rect 248782 2904 248788 2916
rect 247736 2876 248788 2904
rect 247736 2864 247742 2876
rect 248782 2864 248788 2876
rect 248840 2864 248846 2916
rect 291838 2864 291844 2916
rect 291896 2904 291902 2916
rect 293678 2904 293684 2916
rect 291896 2876 293684 2904
rect 291896 2864 291902 2876
rect 293678 2864 293684 2876
rect 293736 2864 293742 2916
rect 318150 2864 318156 2916
rect 318208 2904 318214 2916
rect 319714 2904 319720 2916
rect 318208 2876 319720 2904
rect 318208 2864 318214 2876
rect 319714 2864 319720 2876
rect 319772 2864 319778 2916
rect 448514 2456 448520 2508
rect 448572 2496 448578 2508
rect 449802 2496 449808 2508
rect 448572 2468 449808 2496
rect 448572 2456 448578 2468
rect 449802 2456 449808 2468
rect 449860 2456 449866 2508
rect 415394 2048 415400 2100
rect 415452 2088 415458 2100
rect 416682 2088 416688 2100
rect 415452 2060 416688 2088
rect 415452 2048 415458 2060
rect 416682 2048 416688 2060
rect 416740 2048 416746 2100
rect 440234 2048 440240 2100
rect 440292 2088 440298 2100
rect 441522 2088 441528 2100
rect 440292 2060 441528 2088
rect 440292 2048 440298 2060
rect 441522 2048 441528 2060
rect 441580 2048 441586 2100
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 348792 700340 348844 700392
rect 364340 700340 364392 700392
rect 8116 700272 8168 700324
rect 250444 700272 250496 700324
rect 332508 700272 332560 700324
rect 364432 700272 364484 700324
rect 218980 699660 219032 699712
rect 220084 699660 220136 699712
rect 396724 699660 396776 699712
rect 397460 699660 397512 699712
rect 363604 698640 363656 698692
rect 364984 698640 365036 698692
rect 266360 697552 266412 697604
rect 267648 697552 267700 697604
rect 378784 696940 378836 696992
rect 580172 696940 580224 696992
rect 3424 683136 3476 683188
rect 369860 683136 369912 683188
rect 3424 671032 3476 671084
rect 7564 671032 7616 671084
rect 359464 670692 359516 670744
rect 580172 670692 580224 670744
rect 2780 656956 2832 657008
rect 4804 656956 4856 657008
rect 359556 643084 359608 643136
rect 580172 643084 580224 643136
rect 3424 632068 3476 632120
rect 371424 632068 371476 632120
rect 359648 630640 359700 630692
rect 579988 630640 580040 630692
rect 382924 616836 382976 616888
rect 580172 616836 580224 616888
rect 3516 605820 3568 605872
rect 142804 605820 142856 605872
rect 367744 590656 367796 590708
rect 580172 590656 580224 590708
rect 3332 579640 3384 579692
rect 372620 579640 372672 579692
rect 358452 576852 358504 576904
rect 580172 576852 580224 576904
rect 3240 565836 3292 565888
rect 195244 565836 195296 565888
rect 376024 563048 376076 563100
rect 580172 563048 580224 563100
rect 3332 553392 3384 553444
rect 10324 553392 10376 553444
rect 377404 536800 377456 536852
rect 579896 536800 579948 536852
rect 2964 527144 3016 527196
rect 374000 527144 374052 527196
rect 392584 524424 392636 524476
rect 580172 524424 580224 524476
rect 3516 514768 3568 514820
rect 13084 514768 13136 514820
rect 360844 511232 360896 511284
rect 580264 511232 580316 511284
rect 3056 500964 3108 501016
rect 298744 500964 298796 501016
rect 355324 484372 355376 484424
rect 580172 484372 580224 484424
rect 3056 474716 3108 474768
rect 374092 474716 374144 474768
rect 363696 473968 363748 474020
rect 412640 473968 412692 474020
rect 356704 472608 356756 472660
rect 392584 472608 392636 472660
rect 367836 470568 367888 470620
rect 580080 470568 580132 470620
rect 360936 469820 360988 469872
rect 527180 469820 527232 469872
rect 358084 468460 358136 468512
rect 367744 468460 367796 468512
rect 40040 467100 40092 467152
rect 368572 467100 368624 467152
rect 104900 465672 104952 465724
rect 276020 465672 276072 465724
rect 362316 465672 362368 465724
rect 477500 465672 477552 465724
rect 276020 465060 276072 465112
rect 277308 465060 277360 465112
rect 368664 465060 368716 465112
rect 169760 464312 169812 464364
rect 273260 464312 273312 464364
rect 362224 464312 362276 464364
rect 542360 464312 542412 464364
rect 273260 463700 273312 463752
rect 274548 463700 274600 463752
rect 367100 463700 367152 463752
rect 356244 462952 356296 463004
rect 377404 462952 377456 463004
rect 3516 462544 3568 462596
rect 8944 462544 8996 462596
rect 234620 461592 234672 461644
rect 275284 461592 275336 461644
rect 363052 461592 363104 461644
rect 396724 461592 396776 461644
rect 275284 460912 275336 460964
rect 365812 460912 365864 460964
rect 357256 460232 357308 460284
rect 367836 460232 367888 460284
rect 363236 460164 363288 460216
rect 429200 460164 429252 460216
rect 360660 458804 360712 458856
rect 558920 458804 558972 458856
rect 334716 457104 334768 457156
rect 373540 457104 373592 457156
rect 334900 457036 334952 457088
rect 375748 457036 375800 457088
rect 333520 456968 333572 457020
rect 380164 456968 380216 457020
rect 332048 456900 332100 456952
rect 378232 456900 378284 456952
rect 320824 456832 320876 456884
rect 381268 456832 381320 456884
rect 355968 456764 356020 456816
rect 580172 456764 580224 456816
rect 358636 456084 358688 456136
rect 382924 456084 382976 456136
rect 362316 456016 362368 456068
rect 462320 456016 462372 456068
rect 359188 455880 359240 455932
rect 359648 455880 359700 455932
rect 363512 455880 363564 455932
rect 363696 455880 363748 455932
rect 336464 455812 336516 455864
rect 364432 455812 364484 455864
rect 327816 455744 327868 455796
rect 360476 455744 360528 455796
rect 324964 455676 325016 455728
rect 362500 455676 362552 455728
rect 322204 455608 322256 455660
rect 363512 455608 363564 455660
rect 301504 455540 301556 455592
rect 356704 455540 356756 455592
rect 356980 455540 357032 455592
rect 304264 455472 304316 455524
rect 364340 455472 364392 455524
rect 364708 455472 364760 455524
rect 298836 455404 298888 455456
rect 359188 455404 359240 455456
rect 278596 454928 278648 454980
rect 350724 454928 350776 454980
rect 307024 454860 307076 454912
rect 367192 454860 367244 454912
rect 278688 454792 278740 454844
rect 352104 454792 352156 454844
rect 358728 454792 358780 454844
rect 376024 454792 376076 454844
rect 337936 454724 337988 454776
rect 363236 454724 363288 454776
rect 338028 454656 338080 454708
rect 360660 454656 360712 454708
rect 361580 454656 361632 454708
rect 494060 454656 494112 454708
rect 334624 454588 334676 454640
rect 363328 454588 363380 454640
rect 289820 454520 289872 454572
rect 349988 454520 350040 454572
rect 317604 454452 317656 454504
rect 377588 454452 377640 454504
rect 322388 454384 322440 454436
rect 382464 454384 382516 454436
rect 316868 454316 316920 454368
rect 376944 454316 376996 454368
rect 319444 454248 319496 454300
rect 379796 454248 379848 454300
rect 340788 454180 340840 454232
rect 357624 454180 357676 454232
rect 358728 454180 358780 454232
rect 341524 454112 341576 454164
rect 360936 454112 360988 454164
rect 340512 454044 340564 454096
rect 361580 454044 361632 454096
rect 359096 453976 359148 454028
rect 359556 453976 359608 454028
rect 337844 453568 337896 453620
rect 358084 453568 358136 453620
rect 294604 453500 294656 453552
rect 355416 453500 355468 453552
rect 355968 453500 356020 453552
rect 335084 453432 335136 453484
rect 359096 453432 359148 453484
rect 360384 453432 360436 453484
rect 378784 453432 378836 453484
rect 299480 453364 299532 453416
rect 309048 453364 309100 453416
rect 357348 453296 357400 453348
rect 580356 453296 580408 453348
rect 327908 453228 327960 453280
rect 356060 453228 356112 453280
rect 357256 453228 357308 453280
rect 325056 453160 325108 453212
rect 371240 453160 371292 453212
rect 315304 453092 315356 453144
rect 369952 453092 370004 453144
rect 323676 453024 323728 453076
rect 382740 453024 382792 453076
rect 322296 452956 322348 453008
rect 381636 452956 381688 453008
rect 316776 452888 316828 452940
rect 376116 452888 376168 452940
rect 318064 452820 318116 452872
rect 377220 452820 377272 452872
rect 323584 452752 323636 452804
rect 383844 452752 383896 452804
rect 316684 452684 316736 452736
rect 376760 452684 376812 452736
rect 340696 452616 340748 452668
rect 356336 452616 356388 452668
rect 357348 452616 357400 452668
rect 281264 452140 281316 452192
rect 347412 452140 347464 452192
rect 294696 452072 294748 452124
rect 353668 452072 353720 452124
rect 340144 452004 340196 452056
rect 384580 452004 384632 452056
rect 279884 451936 279936 451988
rect 354864 451936 354916 451988
rect 291844 451868 291896 451920
rect 350540 451868 350592 451920
rect 371240 451868 371292 451920
rect 385040 451868 385092 451920
rect 341800 451800 341852 451852
rect 379060 451800 379112 451852
rect 337384 451732 337436 451784
rect 351460 451732 351512 451784
rect 338764 451664 338816 451716
rect 352564 451664 352616 451716
rect 334808 451596 334860 451648
rect 370228 451596 370280 451648
rect 340972 451528 341024 451580
rect 382556 451528 382608 451580
rect 341616 451460 341668 451512
rect 342260 451392 342312 451444
rect 340328 451256 340380 451308
rect 348148 451324 348200 451376
rect 365812 451392 365864 451444
rect 352196 451324 352248 451376
rect 362224 451324 362276 451376
rect 369124 451324 369176 451376
rect 341892 451256 341944 451308
rect 349252 451256 349304 451308
rect 358544 451256 358596 451308
rect 363972 451256 364024 451308
rect 369952 451256 370004 451308
rect 375380 451256 375432 451308
rect 297364 450848 297416 450900
rect 356244 450848 356296 450900
rect 266360 450780 266412 450832
rect 271328 450780 271380 450832
rect 365720 450780 365772 450832
rect 302884 450712 302936 450764
rect 362316 450712 362368 450764
rect 294788 450644 294840 450696
rect 353300 450644 353352 450696
rect 355232 450644 355284 450696
rect 356704 450644 356756 450696
rect 320916 450576 320968 450628
rect 380532 450576 380584 450628
rect 136640 450508 136692 450560
rect 356244 450508 356296 450560
rect 356612 450508 356664 450560
rect 356704 450508 356756 450560
rect 580264 450508 580316 450560
rect 307760 450440 307812 450492
rect 367652 450440 367704 450492
rect 295984 450372 296036 450424
rect 355324 450372 355376 450424
rect 355508 450372 355560 450424
rect 321008 450304 321060 450356
rect 380900 450304 380952 450356
rect 318156 450236 318208 450288
rect 378324 450236 378376 450288
rect 319536 450168 319588 450220
rect 379658 450168 379710 450220
rect 313924 450100 313976 450152
rect 374506 450100 374558 450152
rect 339316 450032 339368 450084
rect 366548 450032 366600 450084
rect 342168 449964 342220 450016
rect 351092 449964 351144 450016
rect 353300 449964 353352 450016
rect 354128 449964 354180 450016
rect 388444 449964 388496 450016
rect 332232 449896 332284 449948
rect 354772 449896 354824 449948
rect 389824 449896 389876 449948
rect 342352 449488 342404 449540
rect 349620 449488 349672 449540
rect 304356 449284 304408 449336
rect 358544 449420 358596 449472
rect 341708 449352 341760 449404
rect 344100 449352 344152 449404
rect 348516 449352 348568 449404
rect 365076 449420 365128 449472
rect 369860 449420 369912 449472
rect 370596 449420 370648 449472
rect 342444 449284 342496 449336
rect 305644 449216 305696 449268
rect 309048 449216 309100 449268
rect 362224 449352 362276 449404
rect 88340 449148 88392 449200
rect 309140 449148 309192 449200
rect 3056 448604 3108 448656
rect 281540 448604 281592 448656
rect 282828 448604 282880 448656
rect 342444 448604 342496 448656
rect 281172 448536 281224 448588
rect 342352 448536 342404 448588
rect 322480 445000 322532 445052
rect 340972 445000 341024 445052
rect 311164 443640 311216 443692
rect 340880 443640 340932 443692
rect 289728 438132 289780 438184
rect 340972 438132 341024 438184
rect 319628 436704 319680 436756
rect 340972 436704 341024 436756
rect 389824 431876 389876 431928
rect 580172 431876 580224 431928
rect 284944 428408 284996 428460
rect 340972 428408 341024 428460
rect 288348 424328 288400 424380
rect 340328 424328 340380 424380
rect 3516 422288 3568 422340
rect 315580 422288 315632 422340
rect 316776 422288 316828 422340
rect 8944 421540 8996 421592
rect 314660 421540 314712 421592
rect 314660 420860 314712 420912
rect 315396 420860 315448 420912
rect 334900 420860 334952 420912
rect 3424 420180 3476 420232
rect 311900 420180 311952 420232
rect 7564 419432 7616 419484
rect 311164 419432 311216 419484
rect 311900 419432 311952 419484
rect 312636 419432 312688 419484
rect 337660 419432 337712 419484
rect 310704 418140 310756 418192
rect 311164 418140 311216 418192
rect 10324 418072 10376 418124
rect 313556 418072 313608 418124
rect 313556 417664 313608 417716
rect 314016 417664 314068 417716
rect 142804 416032 142856 416084
rect 312728 416032 312780 416084
rect 4804 414672 4856 414724
rect 310520 414672 310572 414724
rect 310520 413924 310572 413976
rect 337476 413924 337528 413976
rect 71780 411884 71832 411936
rect 308128 411884 308180 411936
rect 308128 411204 308180 411256
rect 309048 411204 309100 411256
rect 340236 411204 340288 411256
rect 282920 409164 282972 409216
rect 305000 409164 305052 409216
rect 293224 409096 293276 409148
rect 338764 409096 338816 409148
rect 23480 407736 23532 407788
rect 310428 407736 310480 407788
rect 325148 407736 325200 407788
rect 340144 407736 340196 407788
rect 3424 407056 3476 407108
rect 316224 407056 316276 407108
rect 316868 407056 316920 407108
rect 309876 406988 309928 407040
rect 310428 406988 310480 407040
rect 334808 406988 334860 407040
rect 292028 406376 292080 406428
rect 337384 406376 337436 406428
rect 305000 405628 305052 405680
rect 305736 405628 305788 405680
rect 340972 405628 341024 405680
rect 388996 405628 389048 405680
rect 580172 405628 580224 405680
rect 195244 404948 195296 405000
rect 314016 404948 314068 405000
rect 281540 404268 281592 404320
rect 282000 404268 282052 404320
rect 315304 404268 315356 404320
rect 314016 404200 314068 404252
rect 334716 404200 334768 404252
rect 13084 403588 13136 403640
rect 220176 403588 220228 403640
rect 255964 403588 256016 403640
rect 282000 403588 282052 403640
rect 220176 402976 220228 403028
rect 315488 402976 315540 403028
rect 298744 402908 298796 402960
rect 313924 402908 313976 402960
rect 315580 402840 315632 402892
rect 316132 402840 316184 402892
rect 313372 402228 313424 402280
rect 313924 402228 313976 402280
rect 341892 400936 341944 400988
rect 333336 400528 333388 400580
rect 341708 400596 341760 400648
rect 336188 400460 336240 400512
rect 282092 400392 282144 400444
rect 333888 400392 333940 400444
rect 341800 400392 341852 400444
rect 342260 400392 342312 400444
rect 279976 400324 280028 400376
rect 274456 400256 274508 400308
rect 275836 400188 275888 400240
rect 342260 400188 342312 400240
rect 333888 400120 333940 400172
rect 342076 400052 342128 400104
rect 342260 400052 342312 400104
rect 273168 399644 273220 399696
rect 334348 399916 334400 399968
rect 327540 399848 327592 399900
rect 342858 399848 342910 399900
rect 343042 399848 343094 399900
rect 343318 399848 343370 399900
rect 335820 399780 335872 399832
rect 342950 399780 343002 399832
rect 334900 399712 334952 399764
rect 335636 399644 335688 399696
rect 343870 399848 343922 399900
rect 343962 399848 344014 399900
rect 344146 399848 344198 399900
rect 344330 399848 344382 399900
rect 344698 399848 344750 399900
rect 344882 399848 344934 399900
rect 345250 399848 345302 399900
rect 345526 399848 345578 399900
rect 345802 399848 345854 399900
rect 346078 399848 346130 399900
rect 346262 399848 346314 399900
rect 346446 399848 346498 399900
rect 346538 399848 346590 399900
rect 343502 399780 343554 399832
rect 343502 399644 343554 399696
rect 262128 399576 262180 399628
rect 342076 399576 342128 399628
rect 342260 399576 342312 399628
rect 343778 399780 343830 399832
rect 343686 399712 343738 399764
rect 311164 399508 311216 399560
rect 341892 399508 341944 399560
rect 341984 399508 342036 399560
rect 344054 399780 344106 399832
rect 343962 399712 344014 399764
rect 344284 399644 344336 399696
rect 344836 399644 344888 399696
rect 344008 399576 344060 399628
rect 344100 399576 344152 399628
rect 344744 399576 344796 399628
rect 345388 399576 345440 399628
rect 343916 399508 343968 399560
rect 344560 399508 344612 399560
rect 345710 399780 345762 399832
rect 346170 399780 346222 399832
rect 345756 399576 345808 399628
rect 345940 399576 345992 399628
rect 346124 399576 346176 399628
rect 346492 399712 346544 399764
rect 346308 399576 346360 399628
rect 346906 399848 346958 399900
rect 347458 399848 347510 399900
rect 347642 399848 347694 399900
rect 348010 399848 348062 399900
rect 348286 399848 348338 399900
rect 349574 399848 349626 399900
rect 349666 399848 349718 399900
rect 349758 399848 349810 399900
rect 349942 399848 349994 399900
rect 350310 399848 350362 399900
rect 350586 399848 350638 399900
rect 350770 399848 350822 399900
rect 351046 399848 351098 399900
rect 351138 399848 351190 399900
rect 351230 399848 351282 399900
rect 351414 399848 351466 399900
rect 351690 399848 351742 399900
rect 352058 399848 352110 399900
rect 352242 399848 352294 399900
rect 352426 399848 352478 399900
rect 352794 399848 352846 399900
rect 352978 399848 353030 399900
rect 353898 399848 353950 399900
rect 354082 399848 354134 399900
rect 354266 399848 354318 399900
rect 347274 399780 347326 399832
rect 347044 399644 347096 399696
rect 347504 399644 347556 399696
rect 346768 399576 346820 399628
rect 346952 399576 347004 399628
rect 347320 399576 347372 399628
rect 281448 399440 281500 399492
rect 347228 399440 347280 399492
rect 347872 399576 347924 399628
rect 348102 399780 348154 399832
rect 348194 399780 348246 399832
rect 348378 399780 348430 399832
rect 348240 399644 348292 399696
rect 348148 399576 348200 399628
rect 348056 399440 348108 399492
rect 349436 399508 349488 399560
rect 349804 399644 349856 399696
rect 350034 399780 350086 399832
rect 349620 399440 349672 399492
rect 349988 399440 350040 399492
rect 336280 399372 336332 399424
rect 341800 399372 341852 399424
rect 342260 399372 342312 399424
rect 346400 399372 346452 399424
rect 347688 399372 347740 399424
rect 349896 399372 349948 399424
rect 334716 399304 334768 399356
rect 345664 399304 345716 399356
rect 333796 399236 333848 399288
rect 340052 399168 340104 399220
rect 344560 399168 344612 399220
rect 348700 399304 348752 399356
rect 350402 399780 350454 399832
rect 350678 399780 350730 399832
rect 350954 399780 351006 399832
rect 350816 399712 350868 399764
rect 350724 399644 350776 399696
rect 350908 399644 350960 399696
rect 350448 399576 350500 399628
rect 350632 399576 350684 399628
rect 351184 399644 351236 399696
rect 351644 399712 351696 399764
rect 351276 399576 351328 399628
rect 351460 399576 351512 399628
rect 352380 399508 352432 399560
rect 353760 399644 353812 399696
rect 354404 399644 354456 399696
rect 352932 399576 352984 399628
rect 354036 399576 354088 399628
rect 355462 399848 355514 399900
rect 355738 399848 355790 399900
rect 356290 399848 356342 399900
rect 356474 399848 356526 399900
rect 356566 399848 356618 399900
rect 356750 399848 356802 399900
rect 357302 399848 357354 399900
rect 357394 399848 357446 399900
rect 356106 399780 356158 399832
rect 356520 399712 356572 399764
rect 356934 399780 356986 399832
rect 356152 399644 356204 399696
rect 356428 399644 356480 399696
rect 356796 399644 356848 399696
rect 355232 399508 355284 399560
rect 355416 399508 355468 399560
rect 355692 399508 355744 399560
rect 355968 399508 356020 399560
rect 357164 399576 357216 399628
rect 353576 399440 353628 399492
rect 350264 399372 350316 399424
rect 352104 399372 352156 399424
rect 352472 399372 352524 399424
rect 354220 399372 354272 399424
rect 354772 399372 354824 399424
rect 357256 399440 357308 399492
rect 357670 399848 357722 399900
rect 357946 399848 357998 399900
rect 358130 399848 358182 399900
rect 358682 399848 358734 399900
rect 358958 399848 359010 399900
rect 359142 399848 359194 399900
rect 359234 399848 359286 399900
rect 359878 399848 359930 399900
rect 359970 399848 360022 399900
rect 360246 399848 360298 399900
rect 360338 399848 360390 399900
rect 360430 399848 360482 399900
rect 360522 399848 360574 399900
rect 357532 399576 357584 399628
rect 357762 399780 357814 399832
rect 357808 399576 357860 399628
rect 358314 399780 358366 399832
rect 358360 399644 358412 399696
rect 358268 399576 358320 399628
rect 357624 399508 357676 399560
rect 359004 399576 359056 399628
rect 359694 399780 359746 399832
rect 359280 399576 359332 399628
rect 359188 399508 359240 399560
rect 359740 399576 359792 399628
rect 360016 399712 360068 399764
rect 360200 399576 360252 399628
rect 359924 399508 359976 399560
rect 360706 399780 360758 399832
rect 360476 399508 360528 399560
rect 358728 399440 358780 399492
rect 359648 399440 359700 399492
rect 360384 399440 360436 399492
rect 361074 399848 361126 399900
rect 361258 399848 361310 399900
rect 361350 399848 361402 399900
rect 361442 399848 361494 399900
rect 361626 399848 361678 399900
rect 361810 399848 361862 399900
rect 362454 399848 362506 399900
rect 362822 399848 362874 399900
rect 362914 399848 362966 399900
rect 363006 399848 363058 399900
rect 361120 399576 361172 399628
rect 361488 399712 361540 399764
rect 361396 399644 361448 399696
rect 361580 399644 361632 399696
rect 361764 399576 361816 399628
rect 362730 399780 362782 399832
rect 361304 399508 361356 399560
rect 362592 399508 362644 399560
rect 362960 399712 363012 399764
rect 362868 399644 362920 399696
rect 363190 399780 363242 399832
rect 363144 399644 363196 399696
rect 363236 399576 363288 399628
rect 363558 399848 363610 399900
rect 363742 399848 363794 399900
rect 363926 399848 363978 399900
rect 364110 399848 364162 399900
rect 364294 399848 364346 399900
rect 364386 399848 364438 399900
rect 364570 399848 364622 399900
rect 364846 399848 364898 399900
rect 363466 399780 363518 399832
rect 363834 399780 363886 399832
rect 363696 399712 363748 399764
rect 363604 399644 363656 399696
rect 364156 399712 364208 399764
rect 363880 399576 363932 399628
rect 363604 399508 363656 399560
rect 364340 399508 364392 399560
rect 364432 399508 364484 399560
rect 363788 399440 363840 399492
rect 364064 399440 364116 399492
rect 364800 399644 364852 399696
rect 364616 399508 364668 399560
rect 365582 399848 365634 399900
rect 365674 399848 365726 399900
rect 365766 399848 365818 399900
rect 366226 399848 366278 399900
rect 366410 399848 366462 399900
rect 365214 399780 365266 399832
rect 365398 399780 365450 399832
rect 365260 399644 365312 399696
rect 365858 399780 365910 399832
rect 365950 399780 366002 399832
rect 365812 399644 365864 399696
rect 365904 399644 365956 399696
rect 365720 399576 365772 399628
rect 365168 399508 365220 399560
rect 365352 399508 365404 399560
rect 366088 399644 366140 399696
rect 366180 399508 366232 399560
rect 366686 399848 366738 399900
rect 366778 399848 366830 399900
rect 366870 399848 366922 399900
rect 366824 399576 366876 399628
rect 366640 399440 366692 399492
rect 359556 399372 359608 399424
rect 365996 399372 366048 399424
rect 367054 399848 367106 399900
rect 367422 399848 367474 399900
rect 367790 399848 367842 399900
rect 367974 399848 368026 399900
rect 367514 399780 367566 399832
rect 367376 399644 367428 399696
rect 367468 399644 367520 399696
rect 367744 399644 367796 399696
rect 367192 399576 367244 399628
rect 368066 399780 368118 399832
rect 368158 399780 368210 399832
rect 368020 399644 368072 399696
rect 368112 399576 368164 399628
rect 368342 399848 368394 399900
rect 368618 399848 368670 399900
rect 367100 399508 367152 399560
rect 368434 399780 368486 399832
rect 368526 399780 368578 399832
rect 368296 399440 368348 399492
rect 368986 399848 369038 399900
rect 369446 399848 369498 399900
rect 369906 399848 369958 399900
rect 369998 399848 370050 399900
rect 370182 399848 370234 399900
rect 368848 399576 368900 399628
rect 368572 399508 368624 399560
rect 368480 399440 368532 399492
rect 368664 399440 368716 399492
rect 369216 399712 369268 399764
rect 369124 399576 369176 399628
rect 369814 399780 369866 399832
rect 369860 399576 369912 399628
rect 370090 399780 370142 399832
rect 369952 399508 370004 399560
rect 387524 400324 387576 400376
rect 371378 399848 371430 399900
rect 371930 399848 371982 399900
rect 372390 399848 372442 399900
rect 372574 399848 372626 399900
rect 372942 399848 372994 399900
rect 373494 399848 373546 399900
rect 373954 399848 374006 399900
rect 374046 399848 374098 399900
rect 374322 399848 374374 399900
rect 374598 399848 374650 399900
rect 374874 399848 374926 399900
rect 374966 399848 375018 399900
rect 375518 399848 375570 399900
rect 375610 399848 375662 399900
rect 375886 399848 375938 399900
rect 376070 399848 376122 399900
rect 370550 399780 370602 399832
rect 370596 399644 370648 399696
rect 370504 399576 370556 399628
rect 371976 399712 372028 399764
rect 372528 399644 372580 399696
rect 372620 399644 372672 399696
rect 370320 399508 370372 399560
rect 369676 399440 369728 399492
rect 370136 399440 370188 399492
rect 369400 399372 369452 399424
rect 350908 399304 350960 399356
rect 351184 399304 351236 399356
rect 351276 399304 351328 399356
rect 353208 399304 353260 399356
rect 360292 399304 360344 399356
rect 363052 399304 363104 399356
rect 363420 399304 363472 399356
rect 361028 399236 361080 399288
rect 351184 399168 351236 399220
rect 359556 399168 359608 399220
rect 370688 399304 370740 399356
rect 370964 399304 371016 399356
rect 371516 399304 371568 399356
rect 372804 399576 372856 399628
rect 373264 399508 373316 399560
rect 374368 399508 374420 399560
rect 374644 399508 374696 399560
rect 374736 399508 374788 399560
rect 375472 399712 375524 399764
rect 375012 399576 375064 399628
rect 375978 399780 376030 399832
rect 375932 399644 375984 399696
rect 376024 399576 376076 399628
rect 375932 399508 375984 399560
rect 373540 399440 373592 399492
rect 373724 399440 373776 399492
rect 374000 399440 374052 399492
rect 375656 399372 375708 399424
rect 376438 399848 376490 399900
rect 376622 399848 376674 399900
rect 376484 399712 376536 399764
rect 376898 399848 376950 399900
rect 377082 399848 377134 399900
rect 377266 399848 377318 399900
rect 377634 399848 377686 399900
rect 377818 399848 377870 399900
rect 377910 399848 377962 399900
rect 376944 399712 376996 399764
rect 376852 399508 376904 399560
rect 377680 399644 377732 399696
rect 377772 399644 377824 399696
rect 377864 399576 377916 399628
rect 378094 399848 378146 399900
rect 378278 399848 378330 399900
rect 378646 399848 378698 399900
rect 378922 399848 378974 399900
rect 379014 399848 379066 399900
rect 379106 399848 379158 399900
rect 379382 399848 379434 399900
rect 379842 399848 379894 399900
rect 380302 399848 380354 399900
rect 380486 399848 380538 399900
rect 380762 399848 380814 399900
rect 380946 399848 380998 399900
rect 381314 399848 381366 399900
rect 381406 399848 381458 399900
rect 381498 399848 381550 399900
rect 381682 399848 381734 399900
rect 377496 399508 377548 399560
rect 377956 399508 378008 399560
rect 377128 399440 377180 399492
rect 378692 399712 378744 399764
rect 378416 399576 378468 399628
rect 379566 399780 379618 399832
rect 379428 399712 379480 399764
rect 379060 399644 379112 399696
rect 379336 399508 379388 399560
rect 378508 399440 378560 399492
rect 379796 399712 379848 399764
rect 380532 399644 380584 399696
rect 380808 399644 380860 399696
rect 380256 399508 380308 399560
rect 381452 399644 381504 399696
rect 381544 399644 381596 399696
rect 392032 399984 392084 400036
rect 390560 399916 390612 399968
rect 381958 399848 382010 399900
rect 382142 399848 382194 399900
rect 382418 399848 382470 399900
rect 383062 399848 383114 399900
rect 383246 399848 383298 399900
rect 383706 399848 383758 399900
rect 383890 399848 383942 399900
rect 384258 399848 384310 399900
rect 384626 399848 384678 399900
rect 384810 399848 384862 399900
rect 385454 399848 385506 399900
rect 381820 399644 381872 399696
rect 381084 399576 381136 399628
rect 381268 399576 381320 399628
rect 382188 399644 382240 399696
rect 381176 399508 381228 399560
rect 379888 399440 379940 399492
rect 383108 399712 383160 399764
rect 382556 399508 382608 399560
rect 383936 399644 383988 399696
rect 384120 399644 384172 399696
rect 384580 399644 384632 399696
rect 384948 399644 385000 399696
rect 381176 399372 381228 399424
rect 381452 399372 381504 399424
rect 381636 399372 381688 399424
rect 382096 399372 382148 399424
rect 382280 399372 382332 399424
rect 382556 399372 382608 399424
rect 383568 399372 383620 399424
rect 385730 399848 385782 399900
rect 385914 399848 385966 399900
rect 386006 399848 386058 399900
rect 386190 399848 386242 399900
rect 386374 399848 386426 399900
rect 386926 399848 386978 399900
rect 387018 399848 387070 399900
rect 385868 399644 385920 399696
rect 386052 399644 386104 399696
rect 386466 399780 386518 399832
rect 386328 399712 386380 399764
rect 386788 399644 386840 399696
rect 386420 399576 386472 399628
rect 386972 399644 387024 399696
rect 385592 399508 385644 399560
rect 385684 399508 385736 399560
rect 387984 399440 388036 399492
rect 385684 399372 385736 399424
rect 371700 399304 371752 399356
rect 370228 399236 370280 399288
rect 376300 399236 376352 399288
rect 380164 399236 380216 399288
rect 338948 399100 339000 399152
rect 362960 399100 363012 399152
rect 364248 399100 364300 399152
rect 372712 399168 372764 399220
rect 373908 399168 373960 399220
rect 380256 399168 380308 399220
rect 384488 399168 384540 399220
rect 384948 399168 385000 399220
rect 385776 399168 385828 399220
rect 580264 399440 580316 399492
rect 379612 399100 379664 399152
rect 380532 399100 380584 399152
rect 382096 399100 382148 399152
rect 385868 399100 385920 399152
rect 281356 399032 281408 399084
rect 358176 399032 358228 399084
rect 276848 398964 276900 399016
rect 349160 398964 349212 399016
rect 276756 398896 276808 398948
rect 346216 398896 346268 398948
rect 346676 398896 346728 398948
rect 359740 398964 359792 399016
rect 360292 398964 360344 399016
rect 372252 399032 372304 399084
rect 373908 399032 373960 399084
rect 374276 399032 374328 399084
rect 381912 399032 381964 399084
rect 393320 399032 393372 399084
rect 357808 398896 357860 398948
rect 359004 398896 359056 398948
rect 359556 398896 359608 398948
rect 364248 398896 364300 398948
rect 337660 398828 337712 398880
rect 380624 398964 380676 399016
rect 385868 398964 385920 399016
rect 393504 398964 393556 399016
rect 372252 398896 372304 398948
rect 376300 398896 376352 398948
rect 379612 398896 379664 398948
rect 380808 398896 380860 398948
rect 387524 398896 387576 398948
rect 394976 398896 395028 398948
rect 368940 398828 368992 398880
rect 369308 398828 369360 398880
rect 373816 398828 373868 398880
rect 327724 398760 327776 398812
rect 344652 398760 344704 398812
rect 343456 398692 343508 398744
rect 346400 398760 346452 398812
rect 345112 398692 345164 398744
rect 360476 398760 360528 398812
rect 360844 398760 360896 398812
rect 366548 398760 366600 398812
rect 300400 398624 300452 398676
rect 344284 398624 344336 398676
rect 344468 398624 344520 398676
rect 345480 398624 345532 398676
rect 346216 398624 346268 398676
rect 350448 398624 350500 398676
rect 351828 398624 351880 398676
rect 360660 398692 360712 398744
rect 361488 398692 361540 398744
rect 366548 398624 366600 398676
rect 368940 398624 368992 398676
rect 329196 398556 329248 398608
rect 362408 398556 362460 398608
rect 362868 398556 362920 398608
rect 373908 398556 373960 398608
rect 309968 398488 310020 398540
rect 344468 398488 344520 398540
rect 305092 398420 305144 398472
rect 343640 398420 343692 398472
rect 305000 398352 305052 398404
rect 343824 398352 343876 398404
rect 354772 398488 354824 398540
rect 358176 398488 358228 398540
rect 362316 398488 362368 398540
rect 369768 398488 369820 398540
rect 373448 398488 373500 398540
rect 379888 398828 379940 398880
rect 393412 398828 393464 398880
rect 379796 398760 379848 398812
rect 379980 398760 380032 398812
rect 380164 398760 380216 398812
rect 385776 398760 385828 398812
rect 377956 398692 378008 398744
rect 379980 398624 380032 398676
rect 382648 398692 382700 398744
rect 389272 398692 389324 398744
rect 382832 398624 382884 398676
rect 383016 398624 383068 398676
rect 389180 398556 389232 398608
rect 380900 398488 380952 398540
rect 381452 398488 381504 398540
rect 392216 398488 392268 398540
rect 348332 398420 348384 398472
rect 357348 398420 357400 398472
rect 377588 398420 377640 398472
rect 377956 398420 378008 398472
rect 382372 398420 382424 398472
rect 389640 398420 389692 398472
rect 342076 398284 342128 398336
rect 349160 398352 349212 398404
rect 352196 398352 352248 398404
rect 357072 398352 357124 398404
rect 357624 398352 357676 398404
rect 357992 398352 358044 398404
rect 371148 398352 371200 398404
rect 373264 398352 373316 398404
rect 382832 398352 382884 398404
rect 383660 398352 383712 398404
rect 388168 398352 388220 398404
rect 344284 398284 344336 398336
rect 352012 398284 352064 398336
rect 360660 398284 360712 398336
rect 374552 398284 374604 398336
rect 282920 398216 282972 398268
rect 327540 398216 327592 398268
rect 344560 398216 344612 398268
rect 351184 398216 351236 398268
rect 352288 398216 352340 398268
rect 352656 398216 352708 398268
rect 353392 398216 353444 398268
rect 355324 398216 355376 398268
rect 357624 398216 357676 398268
rect 358820 398216 358872 398268
rect 362224 398216 362276 398268
rect 369676 398216 369728 398268
rect 372252 398216 372304 398268
rect 376760 398216 376812 398268
rect 377588 398216 377640 398268
rect 383660 398216 383712 398268
rect 276940 398148 276992 398200
rect 335636 398148 335688 398200
rect 342536 398148 342588 398200
rect 342720 398148 342772 398200
rect 344100 398148 344152 398200
rect 355416 398148 355468 398200
rect 377128 398148 377180 398200
rect 387800 398148 387852 398200
rect 341892 398080 341944 398132
rect 345112 398080 345164 398132
rect 346400 398080 346452 398132
rect 349160 398080 349212 398132
rect 358820 398080 358872 398132
rect 376760 398080 376812 398132
rect 347044 398012 347096 398064
rect 347688 398012 347740 398064
rect 352012 398012 352064 398064
rect 356244 398012 356296 398064
rect 357164 398012 357216 398064
rect 357348 398012 357400 398064
rect 372528 398012 372580 398064
rect 372712 398012 372764 398064
rect 373356 398012 373408 398064
rect 374000 398012 374052 398064
rect 382556 398012 382608 398064
rect 388076 398012 388128 398064
rect 324228 397944 324280 397996
rect 343916 397944 343968 397996
rect 352656 397944 352708 397996
rect 355600 397944 355652 397996
rect 375380 397944 375432 397996
rect 389364 398148 389416 398200
rect 345664 397876 345716 397928
rect 356520 397876 356572 397928
rect 367836 397876 367888 397928
rect 369032 397876 369084 397928
rect 376576 397876 376628 397928
rect 381452 397876 381504 397928
rect 383292 397876 383344 397928
rect 383568 397876 383620 397928
rect 383936 397876 383988 397928
rect 389456 397876 389508 397928
rect 343732 397808 343784 397860
rect 346584 397808 346636 397860
rect 352748 397808 352800 397860
rect 352932 397808 352984 397860
rect 337752 397740 337804 397792
rect 359372 397808 359424 397860
rect 362868 397808 362920 397860
rect 365812 397808 365864 397860
rect 376208 397808 376260 397860
rect 339132 397672 339184 397724
rect 345664 397672 345716 397724
rect 345848 397672 345900 397724
rect 346216 397672 346268 397724
rect 346584 397672 346636 397724
rect 362040 397740 362092 397792
rect 384488 397808 384540 397860
rect 390928 397808 390980 397860
rect 383568 397740 383620 397792
rect 384212 397740 384264 397792
rect 387892 397740 387944 397792
rect 356336 397672 356388 397724
rect 363696 397672 363748 397724
rect 364156 397672 364208 397724
rect 368664 397672 368716 397724
rect 384672 397672 384724 397724
rect 392308 397672 392360 397724
rect 278504 397604 278556 397656
rect 356612 397604 356664 397656
rect 356796 397604 356848 397656
rect 357164 397604 357216 397656
rect 366548 397604 366600 397656
rect 370412 397604 370464 397656
rect 386696 397604 386748 397656
rect 393136 397604 393188 397656
rect 343824 397536 343876 397588
rect 3424 397468 3476 397520
rect 256884 397468 256936 397520
rect 307668 397468 307720 397520
rect 347872 397536 347924 397588
rect 348884 397536 348936 397588
rect 350816 397536 350868 397588
rect 351276 397536 351328 397588
rect 351920 397536 351972 397588
rect 352196 397536 352248 397588
rect 356888 397536 356940 397588
rect 357348 397536 357400 397588
rect 365812 397536 365864 397588
rect 346584 397468 346636 397520
rect 348148 397468 348200 397520
rect 348608 397468 348660 397520
rect 351184 397468 351236 397520
rect 352380 397468 352432 397520
rect 352748 397468 352800 397520
rect 354588 397468 354640 397520
rect 356612 397468 356664 397520
rect 360200 397468 360252 397520
rect 386788 397536 386840 397588
rect 391940 397536 391992 397588
rect 369124 397468 369176 397520
rect 370780 397468 370832 397520
rect 372620 397468 372672 397520
rect 383660 397468 383712 397520
rect 384396 397468 384448 397520
rect 385868 397468 385920 397520
rect 390744 397468 390796 397520
rect 343088 397400 343140 397452
rect 346952 397400 347004 397452
rect 348516 397400 348568 397452
rect 348884 397400 348936 397452
rect 350172 397400 350224 397452
rect 360752 397400 360804 397452
rect 369492 397400 369544 397452
rect 374552 397400 374604 397452
rect 377312 397400 377364 397452
rect 386052 397400 386104 397452
rect 341156 397332 341208 397384
rect 344008 397332 344060 397384
rect 345664 397332 345716 397384
rect 356612 397332 356664 397384
rect 357348 397332 357400 397384
rect 358452 397332 358504 397384
rect 364984 397332 365036 397384
rect 366272 397332 366324 397384
rect 366456 397332 366508 397384
rect 366732 397332 366784 397384
rect 367008 397332 367060 397384
rect 369860 397332 369912 397384
rect 386696 397332 386748 397384
rect 387340 397332 387392 397384
rect 334808 397264 334860 397316
rect 356152 397264 356204 397316
rect 356796 397264 356848 397316
rect 359464 397264 359516 397316
rect 382280 397264 382332 397316
rect 383200 397264 383252 397316
rect 333428 397196 333480 397248
rect 358912 397196 358964 397248
rect 360476 397196 360528 397248
rect 361212 397196 361264 397248
rect 337476 397128 337528 397180
rect 364432 397128 364484 397180
rect 337568 397060 337620 397112
rect 370136 397060 370188 397112
rect 333244 396992 333296 397044
rect 366824 396992 366876 397044
rect 329104 396924 329156 396976
rect 368112 396924 368164 396976
rect 336648 396856 336700 396908
rect 381544 396924 381596 396976
rect 281540 396788 281592 396840
rect 295340 396788 295392 396840
rect 340420 396788 340472 396840
rect 385408 396788 385460 396840
rect 270132 396720 270184 396772
rect 346124 396720 346176 396772
rect 348516 396720 348568 396772
rect 349896 396720 349948 396772
rect 359464 396720 359516 396772
rect 362684 396720 362736 396772
rect 375564 396720 375616 396772
rect 376576 396720 376628 396772
rect 341984 396652 342036 396704
rect 357256 396652 357308 396704
rect 360292 396652 360344 396704
rect 361580 396652 361632 396704
rect 362040 396652 362092 396704
rect 362500 396652 362552 396704
rect 341708 396584 341760 396636
rect 350172 396584 350224 396636
rect 363604 396584 363656 396636
rect 364248 396584 364300 396636
rect 343364 396516 343416 396568
rect 345940 396516 345992 396568
rect 360568 396516 360620 396568
rect 361396 396516 361448 396568
rect 343640 396448 343692 396500
rect 346768 396448 346820 396500
rect 359740 396448 359792 396500
rect 360108 396448 360160 396500
rect 339040 396380 339092 396432
rect 357440 396380 357492 396432
rect 361672 396380 361724 396432
rect 362592 396380 362644 396432
rect 336372 396312 336424 396364
rect 356244 396312 356296 396364
rect 363696 396312 363748 396364
rect 365352 396312 365404 396364
rect 355508 396176 355560 396228
rect 358268 396176 358320 396228
rect 377312 396176 377364 396228
rect 378232 396176 378284 396228
rect 340236 396108 340288 396160
rect 345664 396108 345716 396160
rect 345848 396040 345900 396092
rect 346032 396040 346084 396092
rect 355600 396040 355652 396092
rect 356980 396040 357032 396092
rect 358268 396040 358320 396092
rect 359096 396040 359148 396092
rect 377404 396040 377456 396092
rect 384672 396040 384724 396092
rect 338764 395972 338816 396024
rect 362868 395972 362920 396024
rect 341800 395904 341852 395956
rect 343548 395904 343600 395956
rect 345848 395904 345900 395956
rect 364892 395904 364944 395956
rect 377864 395904 377916 395956
rect 384212 395904 384264 395956
rect 341340 395836 341392 395888
rect 370688 395836 370740 395888
rect 340328 395768 340380 395820
rect 370964 395768 371016 395820
rect 331864 395700 331916 395752
rect 360844 395700 360896 395752
rect 330944 395632 330996 395684
rect 368020 395632 368072 395684
rect 374736 395632 374788 395684
rect 378692 395632 378744 395684
rect 344192 395564 344244 395616
rect 345020 395564 345072 395616
rect 345296 395564 345348 395616
rect 345572 395564 345624 395616
rect 345664 395564 345716 395616
rect 385316 395564 385368 395616
rect 272984 395496 273036 395548
rect 334900 395496 334952 395548
rect 271604 395428 271656 395480
rect 343364 395428 343416 395480
rect 376392 395428 376444 395480
rect 378692 395428 378744 395480
rect 379060 395428 379112 395480
rect 379796 395428 379848 395480
rect 268476 395360 268528 395412
rect 334348 395360 334400 395412
rect 343916 395360 343968 395412
rect 344376 395360 344428 395412
rect 345204 395360 345256 395412
rect 345756 395360 345808 395412
rect 357716 395360 357768 395412
rect 357900 395360 357952 395412
rect 361120 395360 361172 395412
rect 369952 395360 370004 395412
rect 376668 395360 376720 395412
rect 376944 395360 376996 395412
rect 378324 395360 378376 395412
rect 380256 395360 380308 395412
rect 274364 395292 274416 395344
rect 367652 395292 367704 395344
rect 371792 395292 371844 395344
rect 376760 395292 376812 395344
rect 378508 395292 378560 395344
rect 379428 395292 379480 395344
rect 379796 395292 379848 395344
rect 380348 395292 380400 395344
rect 383292 395292 383344 395344
rect 394792 395292 394844 395344
rect 338672 395224 338724 395276
rect 345664 395224 345716 395276
rect 348240 395224 348292 395276
rect 348792 395224 348844 395276
rect 376392 395224 376444 395276
rect 378140 395224 378192 395276
rect 339960 395156 340012 395208
rect 353484 395156 353536 395208
rect 356796 395156 356848 395208
rect 358636 395156 358688 395208
rect 281632 395088 281684 395140
rect 282920 395088 282972 395140
rect 336096 395088 336148 395140
rect 353760 395088 353812 395140
rect 362132 395088 362184 395140
rect 365720 395088 365772 395140
rect 375656 395088 375708 395140
rect 378140 395088 378192 395140
rect 378784 395088 378836 395140
rect 336004 395020 336056 395072
rect 345848 395020 345900 395072
rect 346492 395020 346544 395072
rect 346676 395020 346728 395072
rect 346768 395020 346820 395072
rect 347596 395020 347648 395072
rect 345388 394952 345440 395004
rect 346308 394952 346360 395004
rect 375656 394884 375708 394936
rect 386328 394884 386380 394936
rect 394884 394884 394936 394936
rect 342904 394816 342956 394868
rect 349160 394816 349212 394868
rect 393136 394748 393188 394800
rect 394700 394748 394752 394800
rect 366456 394680 366508 394732
rect 367100 394680 367152 394732
rect 370504 394680 370556 394732
rect 371240 394680 371292 394732
rect 381544 394680 381596 394732
rect 384304 394680 384356 394732
rect 307668 394612 307720 394664
rect 316316 394612 316368 394664
rect 316684 394612 316736 394664
rect 363236 394612 363288 394664
rect 364708 394612 364760 394664
rect 342536 394544 342588 394596
rect 342996 394544 343048 394596
rect 363144 394544 363196 394596
rect 363328 394544 363380 394596
rect 355876 394408 355928 394460
rect 375288 394408 375340 394460
rect 347688 394340 347740 394392
rect 349068 394340 349120 394392
rect 350816 394340 350868 394392
rect 352840 394340 352892 394392
rect 353668 394340 353720 394392
rect 354496 394340 354548 394392
rect 354588 394340 354640 394392
rect 377036 394340 377088 394392
rect 340604 394272 340656 394324
rect 366732 394272 366784 394324
rect 374276 394272 374328 394324
rect 374644 394272 374696 394324
rect 332140 394204 332192 394256
rect 367928 394204 367980 394256
rect 371240 394204 371292 394256
rect 371516 394204 371568 394256
rect 374368 394204 374420 394256
rect 375288 394204 375340 394256
rect 321376 394136 321428 394188
rect 381084 394136 381136 394188
rect 383844 394136 383896 394188
rect 268844 394068 268896 394120
rect 350816 394068 350868 394120
rect 351000 394068 351052 394120
rect 351644 394068 351696 394120
rect 359556 394068 359608 394120
rect 383108 394068 383160 394120
rect 268752 394000 268804 394052
rect 358176 394000 358228 394052
rect 370228 394000 370280 394052
rect 370872 394000 370924 394052
rect 371516 394000 371568 394052
rect 371884 394000 371936 394052
rect 377220 394000 377272 394052
rect 377864 394000 377916 394052
rect 382556 394000 382608 394052
rect 383384 394000 383436 394052
rect 267372 393932 267424 393984
rect 343180 393864 343232 393916
rect 343456 393864 343508 393916
rect 350816 393932 350868 393984
rect 351368 393932 351420 393984
rect 353392 393932 353444 393984
rect 354128 393932 354180 393984
rect 355416 393932 355468 393984
rect 356060 393932 356112 393984
rect 365904 393932 365956 393984
rect 366272 393932 366324 393984
rect 367284 393932 367336 393984
rect 367928 393932 367980 393984
rect 368572 393932 368624 393984
rect 369124 393932 369176 393984
rect 370136 393932 370188 393984
rect 370596 393932 370648 393984
rect 371792 393932 371844 393984
rect 372344 393932 372396 393984
rect 377036 393932 377088 393984
rect 377772 393932 377824 393984
rect 381084 393932 381136 393984
rect 382004 393932 382056 393984
rect 385132 393932 385184 393984
rect 385316 393932 385368 393984
rect 386604 393932 386656 393984
rect 387340 393932 387392 393984
rect 359924 393864 359976 393916
rect 372712 393864 372764 393916
rect 372988 393864 373040 393916
rect 374368 393864 374420 393916
rect 375012 393864 375064 393916
rect 383844 393864 383896 393916
rect 347964 393796 348016 393848
rect 348332 393796 348384 393848
rect 351092 393796 351144 393848
rect 351644 393796 351696 393848
rect 358176 393796 358228 393848
rect 363512 393796 363564 393848
rect 370596 393796 370648 393848
rect 370780 393796 370832 393848
rect 382740 393796 382792 393848
rect 383292 393796 383344 393848
rect 383752 393796 383804 393848
rect 384764 393796 384816 393848
rect 385040 393796 385092 393848
rect 385776 393796 385828 393848
rect 350724 393728 350776 393780
rect 351736 393728 351788 393780
rect 357072 393728 357124 393780
rect 359556 393728 359608 393780
rect 360844 393728 360896 393780
rect 365628 393728 365680 393780
rect 372988 393728 373040 393780
rect 373540 393728 373592 393780
rect 347780 393660 347832 393712
rect 347964 393660 348016 393712
rect 351276 393660 351328 393712
rect 353576 393660 353628 393712
rect 363696 393660 363748 393712
rect 364156 393660 364208 393712
rect 366916 393660 366968 393712
rect 367468 393660 367520 393712
rect 374092 393660 374144 393712
rect 374828 393660 374880 393712
rect 344652 393592 344704 393644
rect 349436 393592 349488 393644
rect 352656 393592 352708 393644
rect 359648 393592 359700 393644
rect 367192 393592 367244 393644
rect 367560 393592 367612 393644
rect 384212 393524 384264 393576
rect 384672 393524 384724 393576
rect 342996 393456 343048 393508
rect 350632 393456 350684 393508
rect 363512 393456 363564 393508
rect 363972 393456 364024 393508
rect 321284 393388 321336 393440
rect 380900 393388 380952 393440
rect 267556 393320 267608 393372
rect 349344 393320 349396 393372
rect 349436 393320 349488 393372
rect 349620 393320 349672 393372
rect 353944 393320 353996 393372
rect 354588 393320 354640 393372
rect 355324 393320 355376 393372
rect 355876 393320 355928 393372
rect 338856 393048 338908 393100
rect 350448 393116 350500 393168
rect 343180 393048 343232 393100
rect 364248 392980 364300 393032
rect 333612 392912 333664 392964
rect 373724 392912 373776 392964
rect 332324 392844 332376 392896
rect 386420 392912 386472 392964
rect 381268 392844 381320 392896
rect 381728 392844 381780 392896
rect 302148 392776 302200 392828
rect 361580 392776 361632 392828
rect 375380 392776 375432 392828
rect 375932 392776 375984 392828
rect 379336 392776 379388 392828
rect 380072 392776 380124 392828
rect 303344 392708 303396 392760
rect 363144 392708 363196 392760
rect 280988 392640 281040 392692
rect 344928 392640 344980 392692
rect 359096 392640 359148 392692
rect 360016 392640 360068 392692
rect 374184 392640 374236 392692
rect 375104 392640 375156 392692
rect 269856 392572 269908 392624
rect 341156 392572 341208 392624
rect 352840 392572 352892 392624
rect 363052 392572 363104 392624
rect 343824 392504 343876 392556
rect 344560 392504 344612 392556
rect 367376 392504 367428 392556
rect 367744 392504 367796 392556
rect 374552 392504 374604 392556
rect 375196 392504 375248 392556
rect 344100 392436 344152 392488
rect 344744 392436 344796 392488
rect 346492 392368 346544 392420
rect 347136 392368 347188 392420
rect 314292 392096 314344 392148
rect 374000 392096 374052 392148
rect 268936 392028 268988 392080
rect 343088 392028 343140 392080
rect 345940 392028 345992 392080
rect 348700 392028 348752 392080
rect 277032 391960 277084 392012
rect 368480 391960 368532 392012
rect 307944 391892 307996 391944
rect 368204 391892 368256 391944
rect 379888 391824 379940 391876
rect 380716 391824 380768 391876
rect 337384 391756 337436 391808
rect 350356 391756 350408 391808
rect 345664 391688 345716 391740
rect 365536 391688 365588 391740
rect 338580 391620 338632 391672
rect 376116 391620 376168 391672
rect 329288 391552 329340 391604
rect 368572 391552 368624 391604
rect 314384 391484 314436 391536
rect 372620 391484 372672 391536
rect 313188 391416 313240 391468
rect 372712 391416 372764 391468
rect 311808 391348 311860 391400
rect 371240 391348 371292 391400
rect 315856 391280 315908 391332
rect 375472 391280 375524 391332
rect 311716 391212 311768 391264
rect 371332 391212 371384 391264
rect 354220 391144 354272 391196
rect 354404 391144 354456 391196
rect 356888 391144 356940 391196
rect 357348 391144 357400 391196
rect 344376 390736 344428 390788
rect 348976 390736 349028 390788
rect 360660 390736 360712 390788
rect 361304 390736 361356 390788
rect 368756 390736 368808 390788
rect 369584 390736 369636 390788
rect 386604 390736 386656 390788
rect 386880 390736 386932 390788
rect 386880 390600 386932 390652
rect 387432 390600 387484 390652
rect 349620 390464 349672 390516
rect 350080 390464 350132 390516
rect 354220 390192 354272 390244
rect 356336 390192 356388 390244
rect 319812 390056 319864 390108
rect 378140 390056 378192 390108
rect 319904 389988 319956 390040
rect 378968 389988 379020 390040
rect 318708 389920 318760 389972
rect 379428 389920 379480 389972
rect 281724 389852 281776 389904
rect 342444 389852 342496 389904
rect 345756 389852 345808 389904
rect 366180 389852 366232 389904
rect 265992 389784 266044 389836
rect 350540 389784 350592 389836
rect 354128 389784 354180 389836
rect 380992 389784 381044 389836
rect 377956 389716 378008 389768
rect 378140 389716 378192 389768
rect 377680 389648 377732 389700
rect 378048 389648 378100 389700
rect 340144 389104 340196 389156
rect 346768 389104 346820 389156
rect 328000 388968 328052 389020
rect 349712 388968 349764 389020
rect 344928 388900 344980 388952
rect 370136 388900 370188 388952
rect 335268 388832 335320 388884
rect 370228 388832 370280 388884
rect 324596 388764 324648 388816
rect 384856 388764 384908 388816
rect 279608 388696 279660 388748
rect 342536 388696 342588 388748
rect 343088 388696 343140 388748
rect 370044 388696 370096 388748
rect 271512 388628 271564 388680
rect 345296 388628 345348 388680
rect 347412 388628 347464 388680
rect 360568 388628 360620 388680
rect 261944 388560 261996 388612
rect 342260 388560 342312 388612
rect 347136 388560 347188 388612
rect 375380 388560 375432 388612
rect 267648 388492 267700 388544
rect 349344 388492 349396 388544
rect 263416 388424 263468 388476
rect 347872 388424 347924 388476
rect 351368 388424 351420 388476
rect 361212 388424 361264 388476
rect 351276 388152 351328 388204
rect 355048 388152 355100 388204
rect 357624 387472 357676 387524
rect 358544 387472 358596 387524
rect 263324 387336 263376 387388
rect 344836 387336 344888 387388
rect 347320 387336 347372 387388
rect 354956 387336 355008 387388
rect 330852 387268 330904 387320
rect 380256 387268 380308 387320
rect 278412 387200 278464 387252
rect 345204 387200 345256 387252
rect 346032 387200 346084 387252
rect 379888 387200 379940 387252
rect 344100 387132 344152 387184
rect 382280 387132 382332 387184
rect 264888 387064 264940 387116
rect 346400 387064 346452 387116
rect 349804 387064 349856 387116
rect 357716 387064 357768 387116
rect 350080 386520 350132 386572
rect 355692 386520 355744 386572
rect 320180 386316 320232 386368
rect 321008 386316 321060 386368
rect 322940 386316 322992 386368
rect 323768 386316 323820 386368
rect 330668 386112 330720 386164
rect 374736 386112 374788 386164
rect 329472 386044 329524 386096
rect 377956 386044 378008 386096
rect 333704 385976 333756 386028
rect 385960 385976 386012 386028
rect 282736 385908 282788 385960
rect 339960 385908 340012 385960
rect 265900 385840 265952 385892
rect 346676 385840 346728 385892
rect 276664 385772 276716 385824
rect 363512 385772 363564 385824
rect 280896 385704 280948 385756
rect 369768 385704 369820 385756
rect 273812 385636 273864 385688
rect 365904 385636 365956 385688
rect 271144 385160 271196 385212
rect 320180 385160 320232 385212
rect 262956 385092 263008 385144
rect 322940 385092 322992 385144
rect 264336 385024 264388 385076
rect 324596 385024 324648 385076
rect 319076 384956 319128 385008
rect 319720 384956 319772 385008
rect 321744 384956 321796 385008
rect 322388 384956 322440 385008
rect 259184 384276 259236 384328
rect 348240 384276 348292 384328
rect 265624 383800 265676 383852
rect 324320 383800 324372 383852
rect 261484 383732 261536 383784
rect 321744 383732 321796 383784
rect 258724 383664 258776 383716
rect 319076 383664 319128 383716
rect 343548 383460 343600 383512
rect 359096 383460 359148 383512
rect 343456 383392 343508 383444
rect 367744 383392 367796 383444
rect 331036 383324 331088 383376
rect 379796 383324 379848 383376
rect 332416 383256 332468 383308
rect 382556 383256 382608 383308
rect 274088 383188 274140 383240
rect 348608 383188 348660 383240
rect 349896 383188 349948 383240
rect 361856 383188 361908 383240
rect 277768 383120 277820 383172
rect 360476 383120 360528 383172
rect 269948 383052 270000 383104
rect 354496 383052 354548 383104
rect 263232 382984 263284 383036
rect 348148 382984 348200 383036
rect 348608 382984 348660 383036
rect 360200 382984 360252 383036
rect 280804 382916 280856 382968
rect 372988 382916 373040 382968
rect 321652 382644 321704 382696
rect 322480 382644 322532 382696
rect 271236 382372 271288 382424
rect 321652 382440 321704 382492
rect 318892 382372 318944 382424
rect 319628 382372 319680 382424
rect 260104 382304 260156 382356
rect 257344 382236 257396 382288
rect 318892 382236 318944 382288
rect 318984 382236 319036 382288
rect 319444 382236 319496 382288
rect 323032 381692 323084 381744
rect 323676 381692 323728 381744
rect 320272 381284 320324 381336
rect 320824 381284 320876 381336
rect 272616 381012 272668 381064
rect 320272 381012 320324 381064
rect 253848 380944 253900 380996
rect 313372 380944 313424 380996
rect 262864 380876 262916 380928
rect 323032 380876 323084 380928
rect 314844 380332 314896 380384
rect 315304 380332 315356 380384
rect 281816 380196 281868 380248
rect 342720 380196 342772 380248
rect 261852 380128 261904 380180
rect 348056 380128 348108 380180
rect 272708 379856 272760 379908
rect 314844 379856 314896 379908
rect 244924 379788 244976 379840
rect 303620 379788 303672 379840
rect 304264 379788 304316 379840
rect 249064 379720 249116 379772
rect 309140 379720 309192 379772
rect 264704 379652 264756 379704
rect 264428 379584 264480 379636
rect 324504 379584 324556 379636
rect 325148 379584 325200 379636
rect 259368 379516 259420 379568
rect 320916 379516 320968 379568
rect 324320 379516 324372 379568
rect 325056 379516 325108 379568
rect 345848 379516 345900 379568
rect 353576 379516 353628 379568
rect 254124 378292 254176 378344
rect 313924 378428 313976 378480
rect 259736 378224 259788 378276
rect 319536 378360 319588 378412
rect 313924 378224 313976 378276
rect 314200 378224 314252 378276
rect 263508 378156 263560 378208
rect 323860 378156 323912 378208
rect 348700 378020 348752 378072
rect 357256 378020 357308 378072
rect 348792 377544 348844 377596
rect 359004 377544 359056 377596
rect 350172 377476 350224 377528
rect 363236 377476 363288 377528
rect 281908 377408 281960 377460
rect 342628 377408 342680 377460
rect 348516 377408 348568 377460
rect 367376 377408 367428 377460
rect 264244 376932 264296 376984
rect 311992 376932 312044 376984
rect 312544 376932 312596 376984
rect 242164 376864 242216 376916
rect 301596 376864 301648 376916
rect 255504 376796 255556 376848
rect 316132 376796 316184 376848
rect 245016 376728 245068 376780
rect 307852 376728 307904 376780
rect 291292 376116 291344 376168
rect 291936 376116 291988 376168
rect 292304 376116 292356 376168
rect 275376 376048 275428 376100
rect 293040 376048 293092 376100
rect 274180 375980 274232 376032
rect 292212 375980 292264 376032
rect 275652 375912 275704 375964
rect 298560 375912 298612 375964
rect 274272 375844 274324 375896
rect 302608 375844 302660 375896
rect 279700 375776 279752 375828
rect 312912 375776 312964 375828
rect 264520 375708 264572 375760
rect 300216 375708 300268 375760
rect 267096 375640 267148 375692
rect 311072 375640 311124 375692
rect 232504 375572 232556 375624
rect 291292 375572 291344 375624
rect 298560 375572 298612 375624
rect 298928 375572 298980 375624
rect 236644 375504 236696 375556
rect 297456 375504 297508 375556
rect 301504 375504 301556 375556
rect 238668 375436 238720 375488
rect 298836 375436 298888 375488
rect 261300 375368 261352 375420
rect 321836 375368 321888 375420
rect 322296 375368 322348 375420
rect 268384 374756 268436 374808
rect 293316 374756 293368 374808
rect 294328 374756 294380 374808
rect 294788 374756 294840 374808
rect 318432 374756 318484 374808
rect 267188 374688 267240 374740
rect 275284 374688 275336 374740
rect 306196 374688 306248 374740
rect 318892 374688 318944 374740
rect 319168 374688 319220 374740
rect 320180 374688 320232 374740
rect 321008 374688 321060 374740
rect 324320 374756 324372 374808
rect 324964 374756 325016 374808
rect 332048 374688 332100 374740
rect 219256 374620 219308 374672
rect 282828 374620 282880 374672
rect 299388 374620 299440 374672
rect 340788 374620 340840 374672
rect 267280 374552 267332 374604
rect 295800 374552 295852 374604
rect 321652 374552 321704 374604
rect 322388 374552 322440 374604
rect 324504 374552 324556 374604
rect 324688 374552 324740 374604
rect 277308 374484 277360 374536
rect 308404 374484 308456 374536
rect 324412 374484 324464 374536
rect 325332 374484 325384 374536
rect 272340 374416 272392 374468
rect 303252 374416 303304 374468
rect 273076 374348 273128 374400
rect 304356 374348 304408 374400
rect 269764 374280 269816 374332
rect 305368 374280 305420 374332
rect 277860 374212 277912 374264
rect 317972 374212 318024 374264
rect 318432 374212 318484 374264
rect 245108 374144 245160 374196
rect 297088 374144 297140 374196
rect 238852 374076 238904 374128
rect 298836 374076 298888 374128
rect 219348 374008 219400 374060
rect 294328 374008 294380 374060
rect 153200 373940 153252 373992
rect 280160 373940 280212 373992
rect 220084 373872 220136 373924
rect 282276 373872 282328 373924
rect 297364 373872 297416 373924
rect 307116 373872 307168 373924
rect 314936 373600 314988 373652
rect 315488 373600 315540 373652
rect 304172 373464 304224 373516
rect 304356 373464 304408 373516
rect 300860 373396 300912 373448
rect 338028 373396 338080 373448
rect 294512 373328 294564 373380
rect 332232 373328 332284 373380
rect 220728 373260 220780 373312
rect 281264 373260 281316 373312
rect 287428 373260 287480 373312
rect 296628 373260 296680 373312
rect 340696 373260 340748 373312
rect 233884 373192 233936 373244
rect 294512 373192 294564 373244
rect 278136 373124 278188 373176
rect 294604 373124 294656 373176
rect 295340 373124 295392 373176
rect 275192 373056 275244 373108
rect 297824 373056 297876 373108
rect 299388 373056 299440 373108
rect 279056 372988 279108 373040
rect 299940 372988 299992 373040
rect 300308 372988 300360 373040
rect 313372 372988 313424 373040
rect 314660 372988 314712 373040
rect 322848 372988 322900 373040
rect 323032 372988 323084 373040
rect 275100 372920 275152 372972
rect 298744 372920 298796 372972
rect 275744 372852 275796 372904
rect 300860 372852 300912 372904
rect 277216 372784 277268 372836
rect 303528 372784 303580 372836
rect 272432 372716 272484 372768
rect 301044 372716 301096 372768
rect 274548 372648 274600 372700
rect 278228 372580 278280 372632
rect 296628 372580 296680 372632
rect 307300 372512 307352 372564
rect 314936 372512 314988 372564
rect 358360 372512 358412 372564
rect 298836 372444 298888 372496
rect 335084 372444 335136 372496
rect 303252 372376 303304 372428
rect 337936 372376 337988 372428
rect 303528 372308 303580 372360
rect 334624 372308 334676 372360
rect 278044 372240 278096 372292
rect 288256 372240 288308 372292
rect 280160 372104 280212 372156
rect 287704 372104 287756 372156
rect 288256 372104 288308 372156
rect 273904 372036 273956 372088
rect 282736 372036 282788 372088
rect 282920 372036 282972 372088
rect 288532 372036 288584 372088
rect 293868 372104 293920 372156
rect 294788 372104 294840 372156
rect 329656 372104 329708 372156
rect 328368 372036 328420 372088
rect 279884 371968 279936 372020
rect 294788 371968 294840 372020
rect 229744 371900 229796 371952
rect 281080 371900 281132 371952
rect 286324 371900 286376 371952
rect 220636 371832 220688 371884
rect 281172 371832 281224 371884
rect 282736 371832 282788 371884
rect 283656 371832 283708 371884
rect 287612 371832 287664 371884
rect 293868 371832 293920 371884
rect 282276 371764 282328 371816
rect 304080 371832 304132 371884
rect 322204 371832 322256 371884
rect 332784 371832 332836 371884
rect 346216 371832 346268 371884
rect 282184 371696 282236 371748
rect 305828 371696 305880 371748
rect 280712 371628 280764 371680
rect 285220 371628 285272 371680
rect 287704 371628 287756 371680
rect 308312 371696 308364 371748
rect 307760 371628 307812 371680
rect 318064 371628 318116 371680
rect 281264 371560 281316 371612
rect 312636 371560 312688 371612
rect 312820 371560 312872 371612
rect 316224 371560 316276 371612
rect 316868 371560 316920 371612
rect 280620 371492 280672 371544
rect 314016 371492 314068 371544
rect 277952 371424 278004 371476
rect 279884 371424 279936 371476
rect 280712 371424 280764 371476
rect 332600 371492 332652 371544
rect 333520 371492 333572 371544
rect 279240 371356 279292 371408
rect 315764 371356 315816 371408
rect 320640 371356 320692 371408
rect 332600 371356 332652 371408
rect 279516 371288 279568 371340
rect 287612 371288 287664 371340
rect 288348 371288 288400 371340
rect 291844 371288 291896 371340
rect 323584 371288 323636 371340
rect 333980 371288 334032 371340
rect 3424 371220 3476 371272
rect 257068 371220 257120 371272
rect 279332 371220 279384 371272
rect 287152 371220 287204 371272
rect 289728 371220 289780 371272
rect 290740 371220 290792 371272
rect 326252 371220 326304 371272
rect 332784 371220 332836 371272
rect 307760 371152 307812 371204
rect 278596 371084 278648 371136
rect 289728 371084 289780 371136
rect 233148 370676 233200 370728
rect 278688 371016 278740 371068
rect 288348 371016 288400 371068
rect 300308 370880 300360 370932
rect 327816 370880 327868 370932
rect 305092 370812 305144 370864
rect 336464 370812 336516 370864
rect 271328 370744 271380 370796
rect 305460 370744 305512 370796
rect 301504 370676 301556 370728
rect 341524 370676 341576 370728
rect 231768 370608 231820 370660
rect 278596 370608 278648 370660
rect 298100 370608 298152 370660
rect 337844 370608 337896 370660
rect 245752 370540 245804 370592
rect 271328 370540 271380 370592
rect 276572 370540 276624 370592
rect 333796 370540 333848 370592
rect 258816 370472 258868 370524
rect 318340 370472 318392 370524
rect 278320 370404 278372 370456
rect 285128 370404 285180 370456
rect 235264 370336 235316 370388
rect 295892 370336 295944 370388
rect 264612 370268 264664 370320
rect 300308 370268 300360 370320
rect 279884 370200 279936 370252
rect 306564 370200 306616 370252
rect 245200 370132 245252 370184
rect 305092 370132 305144 370184
rect 281080 370064 281132 370116
rect 317604 370064 317656 370116
rect 318984 370064 319036 370116
rect 320042 370064 320094 370116
rect 320272 370064 320324 370116
rect 321514 370064 321566 370116
rect 238024 369996 238076 370048
rect 298100 369996 298152 370048
rect 301044 369996 301096 370048
rect 301872 369996 301924 370048
rect 340512 369996 340564 370048
rect 293040 369928 293092 369980
rect 534724 369928 534776 369980
rect 292580 369860 292632 369912
rect 577596 369860 577648 369912
rect 291568 369792 291620 369844
rect 340880 369792 340932 369844
rect 304724 369724 304776 369776
rect 305092 369724 305144 369776
rect 317604 369724 317656 369776
rect 318064 369724 318116 369776
rect 291936 369588 291988 369640
rect 292212 369588 292264 369640
rect 233976 369112 234028 369164
rect 281448 369112 281500 369164
rect 229836 368636 229888 368688
rect 288992 369384 289044 369436
rect 291476 369384 291528 369436
rect 301412 369520 301464 369572
rect 296352 369452 296404 369504
rect 310612 369588 310664 369640
rect 310980 369588 311032 369640
rect 306932 369384 306984 369436
rect 231124 368568 231176 368620
rect 240140 368500 240192 368552
rect 340880 369180 340932 369232
rect 342168 369180 342220 369232
rect 580632 369180 580684 369232
rect 580356 369112 580408 369164
rect 327908 368568 327960 368620
rect 339316 368500 339368 368552
rect 201500 367752 201552 367804
rect 245660 367752 245712 367804
rect 245660 367004 245712 367056
rect 246304 367004 246356 367056
rect 279884 367004 279936 367056
rect 329748 366324 329800 366376
rect 384028 366324 384080 366376
rect 329656 365644 329708 365696
rect 580172 365644 580224 365696
rect 247040 365032 247092 365084
rect 274548 365032 274600 365084
rect 247684 364964 247736 365016
rect 280160 364964 280212 365016
rect 249156 363604 249208 363656
rect 277308 363604 277360 363656
rect 334992 362176 335044 362228
rect 350816 362176 350868 362228
rect 253388 360816 253440 360868
rect 280620 360816 280672 360868
rect 333520 359524 333572 359576
rect 352104 359524 352156 359576
rect 256792 359456 256844 359508
rect 280712 359456 280764 359508
rect 329656 359456 329708 359508
rect 385408 359456 385460 359508
rect 226984 358776 227036 358828
rect 277676 358776 277728 358828
rect 279424 358776 279476 358828
rect 271052 358708 271104 358760
rect 277860 358708 277912 358760
rect 3148 357416 3200 357468
rect 271052 357416 271104 357468
rect 253296 356668 253348 356720
rect 280712 356668 280764 356720
rect 333796 356668 333848 356720
rect 350724 356668 350776 356720
rect 256056 355308 256108 355360
rect 279240 355308 279292 355360
rect 227076 351160 227128 351212
rect 279332 351160 279384 351212
rect 383844 349052 383896 349104
rect 384396 349052 384448 349104
rect 384396 347760 384448 347812
rect 534080 347760 534132 347812
rect 332048 347012 332100 347064
rect 351552 347012 351604 347064
rect 255412 345652 255464 345704
rect 280712 345652 280764 345704
rect 3332 345040 3384 345092
rect 255412 345040 255464 345092
rect 332232 342864 332284 342916
rect 350264 342864 350316 342916
rect 332508 340144 332560 340196
rect 351644 340144 351696 340196
rect 329012 338716 329064 338768
rect 386972 338716 387024 338768
rect 350264 335996 350316 336048
rect 368756 335996 368808 336048
rect 336464 334568 336516 334620
rect 377036 334568 377088 334620
rect 385224 333956 385276 334008
rect 385684 333956 385736 334008
rect 552020 333956 552072 334008
rect 335176 333208 335228 333260
rect 371792 333208 371844 333260
rect 379704 331236 379756 331288
rect 481640 331236 481692 331288
rect 331128 329060 331180 329112
rect 345572 329060 345624 329112
rect 235356 327700 235408 327752
rect 277952 327700 278004 327752
rect 380900 327088 380952 327140
rect 381360 327088 381412 327140
rect 495440 327088 495492 327140
rect 336924 326340 336976 326392
rect 375656 326340 375708 326392
rect 577596 325456 577648 325508
rect 580724 325456 580776 325508
rect 234068 324912 234120 324964
rect 279516 324912 279568 324964
rect 385776 324300 385828 324352
rect 547972 324300 548024 324352
rect 339316 323620 339368 323672
rect 378416 323620 378468 323672
rect 335084 323552 335136 323604
rect 374368 323552 374420 323604
rect 380900 323008 380952 323060
rect 381268 323008 381320 323060
rect 381544 322940 381596 322992
rect 383384 322940 383436 322992
rect 506480 322940 506532 322992
rect 272248 322260 272300 322312
rect 273168 322260 273220 322312
rect 339960 322260 340012 322312
rect 363696 322260 363748 322312
rect 228456 322192 228508 322244
rect 278044 322192 278096 322244
rect 334072 322192 334124 322244
rect 380900 322192 380952 322244
rect 272524 322124 272576 322176
rect 273168 322124 273220 322176
rect 218704 321716 218756 321768
rect 268568 321716 268620 321768
rect 206744 321648 206796 321700
rect 272524 321648 272576 321700
rect 201408 321580 201460 321632
rect 269856 321580 269908 321632
rect 270316 321580 270368 321632
rect 327908 321376 327960 321428
rect 328184 321376 328236 321428
rect 271328 321104 271380 321156
rect 271604 321104 271656 321156
rect 327816 321104 327868 321156
rect 328092 321104 328144 321156
rect 271604 320968 271656 321020
rect 271788 320968 271840 321020
rect 272984 320900 273036 320952
rect 276756 321036 276808 321088
rect 337016 321036 337068 321088
rect 368664 321036 368716 321088
rect 299894 320696 299946 320748
rect 353392 320968 353444 321020
rect 333152 320900 333204 320952
rect 359556 320900 359608 320952
rect 217876 320492 217928 320544
rect 281632 320560 281684 320612
rect 282276 320560 282328 320612
rect 276848 320424 276900 320476
rect 282184 320424 282236 320476
rect 220544 320220 220596 320272
rect 282184 320152 282236 320204
rect 278504 320084 278556 320136
rect 279976 319948 280028 320000
rect 282184 319948 282236 320000
rect 278044 319880 278096 319932
rect 281908 319744 281960 319796
rect 282368 319744 282420 319796
rect 287152 319744 287204 319796
rect 216312 319540 216364 319592
rect 273904 319676 273956 319728
rect 289038 319880 289090 319932
rect 288808 319676 288860 319728
rect 293500 319744 293552 319796
rect 294512 319880 294564 319932
rect 295018 319880 295070 319932
rect 294788 319812 294840 319864
rect 295754 319880 295806 319932
rect 296858 319880 296910 319932
rect 357440 320832 357492 320884
rect 297088 319812 297140 319864
rect 333152 320696 333204 320748
rect 328460 320628 328512 320680
rect 327632 320492 327684 320544
rect 298790 319880 298842 319932
rect 300170 319880 300222 319932
rect 301550 319880 301602 319932
rect 298560 319812 298612 319864
rect 300538 319812 300590 319864
rect 300768 319812 300820 319864
rect 301320 319744 301372 319796
rect 302378 319880 302430 319932
rect 303022 319880 303074 319932
rect 303206 319880 303258 319932
rect 304034 319880 304086 319932
rect 304310 319880 304362 319932
rect 304402 319880 304454 319932
rect 305322 319880 305374 319932
rect 302148 319812 302200 319864
rect 280068 319608 280120 319660
rect 292488 319608 292540 319660
rect 292672 319608 292724 319660
rect 296904 319608 296956 319660
rect 299756 319608 299808 319660
rect 300860 319608 300912 319660
rect 301136 319608 301188 319660
rect 276572 319540 276624 319592
rect 300952 319540 301004 319592
rect 301504 319540 301556 319592
rect 302240 319744 302292 319796
rect 302240 319608 302292 319660
rect 302470 319812 302522 319864
rect 302332 319540 302384 319592
rect 302608 319540 302660 319592
rect 302792 319540 302844 319592
rect 303666 319812 303718 319864
rect 303620 319676 303672 319728
rect 303988 319676 304040 319728
rect 303344 319608 303396 319660
rect 304494 319812 304546 319864
rect 304862 319812 304914 319864
rect 303160 319540 303212 319592
rect 304356 319540 304408 319592
rect 304816 319608 304868 319660
rect 306242 319812 306294 319864
rect 305460 319676 305512 319728
rect 305828 319608 305880 319660
rect 211068 319404 211120 319456
rect 272892 319472 272944 319524
rect 293132 319472 293184 319524
rect 294604 319472 294656 319524
rect 294972 319472 295024 319524
rect 295892 319472 295944 319524
rect 296168 319472 296220 319524
rect 296904 319472 296956 319524
rect 298100 319472 298152 319524
rect 273812 319404 273864 319456
rect 304448 319472 304500 319524
rect 306794 319880 306846 319932
rect 307438 319880 307490 319932
rect 307530 319880 307582 319932
rect 306564 319676 306616 319728
rect 307484 319676 307536 319728
rect 335544 320356 335596 320408
rect 310244 319880 310296 319932
rect 310152 319812 310204 319864
rect 342352 320288 342404 320340
rect 328460 320220 328512 320272
rect 335452 320220 335504 320272
rect 311210 319880 311262 319932
rect 337016 320152 337068 320204
rect 328276 320084 328328 320136
rect 313142 319880 313194 319932
rect 311992 319812 312044 319864
rect 310520 319608 310572 319660
rect 310612 319608 310664 319660
rect 311900 319608 311952 319660
rect 310336 319540 310388 319592
rect 312268 319540 312320 319592
rect 313188 319540 313240 319592
rect 313786 319880 313838 319932
rect 314062 319880 314114 319932
rect 314614 319880 314666 319932
rect 314706 319880 314758 319932
rect 315350 319880 315402 319932
rect 315534 319880 315586 319932
rect 314568 319608 314620 319660
rect 313556 319540 313608 319592
rect 314384 319540 314436 319592
rect 315120 319608 315172 319660
rect 317282 319880 317334 319932
rect 317834 319880 317886 319932
rect 317926 319812 317978 319864
rect 317144 319744 317196 319796
rect 317236 319744 317288 319796
rect 317788 319744 317840 319796
rect 318248 319744 318300 319796
rect 317880 319676 317932 319728
rect 315580 319608 315632 319660
rect 317144 319608 317196 319660
rect 314844 319540 314896 319592
rect 315488 319540 315540 319592
rect 315672 319540 315724 319592
rect 320870 319880 320922 319932
rect 320962 319880 321014 319932
rect 319582 319812 319634 319864
rect 319858 319812 319910 319864
rect 320732 319744 320784 319796
rect 320916 319676 320968 319728
rect 321422 319880 321474 319932
rect 322158 319880 322210 319932
rect 322802 319880 322854 319932
rect 323998 319880 324050 319932
rect 319628 319608 319680 319660
rect 319904 319608 319956 319660
rect 321284 319608 321336 319660
rect 321698 319812 321750 319864
rect 322020 319744 322072 319796
rect 322710 319812 322762 319864
rect 321744 319608 321796 319660
rect 322020 319608 322072 319660
rect 322204 319608 322256 319660
rect 322480 319608 322532 319660
rect 309784 319404 309836 319456
rect 309968 319404 310020 319456
rect 312820 319472 312872 319524
rect 321560 319540 321612 319592
rect 321652 319540 321704 319592
rect 323492 319812 323544 319864
rect 322756 319676 322808 319728
rect 323400 319676 323452 319728
rect 323860 319676 323912 319728
rect 327632 320016 327684 320068
rect 325102 319880 325154 319932
rect 329932 319948 329984 320000
rect 326666 319880 326718 319932
rect 327126 319880 327178 319932
rect 327632 319880 327684 319932
rect 325286 319812 325338 319864
rect 325056 319676 325108 319728
rect 326436 319744 326488 319796
rect 325700 319676 325752 319728
rect 326758 319812 326810 319864
rect 327080 319744 327132 319796
rect 327172 319744 327224 319796
rect 335360 319744 335412 319796
rect 326620 319676 326672 319728
rect 326804 319676 326856 319728
rect 332324 319676 332376 319728
rect 323492 319608 323544 319660
rect 354864 319608 354916 319660
rect 318064 319472 318116 319524
rect 318248 319472 318300 319524
rect 318340 319472 318392 319524
rect 343364 319540 343416 319592
rect 326344 319472 326396 319524
rect 327172 319472 327224 319524
rect 327356 319472 327408 319524
rect 361764 319472 361816 319524
rect 323492 319404 323544 319456
rect 325056 319404 325108 319456
rect 325332 319404 325384 319456
rect 329932 319404 329984 319456
rect 330116 319404 330168 319456
rect 371700 319404 371752 319456
rect 282920 319336 282972 319388
rect 283104 319336 283156 319388
rect 283380 319336 283432 319388
rect 283564 319336 283616 319388
rect 285220 319336 285272 319388
rect 285680 319336 285732 319388
rect 287520 319336 287572 319388
rect 287980 319336 288032 319388
rect 288900 319336 288952 319388
rect 289820 319336 289872 319388
rect 291292 319336 291344 319388
rect 292028 319336 292080 319388
rect 206652 319268 206704 319320
rect 276480 319200 276532 319252
rect 279976 319200 280028 319252
rect 278320 319132 278372 319184
rect 280068 319132 280120 319184
rect 3424 318792 3476 318844
rect 197360 318792 197412 318844
rect 258264 319064 258316 319116
rect 258816 319064 258868 319116
rect 275928 319064 275980 319116
rect 283104 319064 283156 319116
rect 285036 319268 285088 319320
rect 285588 319268 285640 319320
rect 290004 319268 290056 319320
rect 290372 319268 290424 319320
rect 345940 319336 345992 319388
rect 292764 319268 292816 319320
rect 352932 319268 352984 319320
rect 284484 319200 284536 319252
rect 343916 319200 343968 319252
rect 287152 319132 287204 319184
rect 346492 319132 346544 319184
rect 288992 319064 289044 319116
rect 347964 319064 348016 319116
rect 224316 318996 224368 319048
rect 292764 318996 292816 319048
rect 292948 318996 293000 319048
rect 294420 318996 294472 319048
rect 294788 318996 294840 319048
rect 298560 318996 298612 319048
rect 301136 318996 301188 319048
rect 301688 318996 301740 319048
rect 302516 318996 302568 319048
rect 303160 318996 303212 319048
rect 303712 318996 303764 319048
rect 352472 318996 352524 319048
rect 208216 318928 208268 318980
rect 286968 318928 287020 318980
rect 206560 318860 206612 318912
rect 278044 318860 278096 318912
rect 279516 318860 279568 318912
rect 295984 318860 296036 318912
rect 346584 318928 346636 318980
rect 313464 318860 313516 318912
rect 314568 318860 314620 318912
rect 317972 318860 318024 318912
rect 318340 318860 318392 318912
rect 319536 318860 319588 318912
rect 319720 318860 319772 318912
rect 320088 318860 320140 318912
rect 379060 318860 379112 318912
rect 275560 318792 275612 318844
rect 276848 318792 276900 318844
rect 277676 318792 277728 318844
rect 278504 318792 278556 318844
rect 279792 318792 279844 318844
rect 281448 318792 281500 318844
rect 281908 318792 281960 318844
rect 282184 318792 282236 318844
rect 292948 318792 293000 318844
rect 293592 318792 293644 318844
rect 303712 318792 303764 318844
rect 320180 318792 320232 318844
rect 322940 318792 322992 318844
rect 325424 318792 325476 318844
rect 327356 318792 327408 318844
rect 335360 318792 335412 318844
rect 336464 318792 336516 318844
rect 282092 318724 282144 318776
rect 282460 318724 282512 318776
rect 285312 318724 285364 318776
rect 291660 318724 291712 318776
rect 291936 318724 291988 318776
rect 295984 318724 296036 318776
rect 296444 318724 296496 318776
rect 297272 318724 297324 318776
rect 297456 318724 297508 318776
rect 310980 318724 311032 318776
rect 314568 318724 314620 318776
rect 317788 318724 317840 318776
rect 322480 318724 322532 318776
rect 325884 318724 325936 318776
rect 329656 318724 329708 318776
rect 331772 318724 331824 318776
rect 357072 318724 357124 318776
rect 269304 318656 269356 318708
rect 274088 318656 274140 318708
rect 288164 318656 288216 318708
rect 290464 318656 290516 318708
rect 276940 318588 276992 318640
rect 284208 318588 284260 318640
rect 290648 318588 290700 318640
rect 270224 318520 270276 318572
rect 278044 318520 278096 318572
rect 270040 318452 270092 318504
rect 274456 318452 274508 318504
rect 292304 318520 292356 318572
rect 300860 318656 300912 318708
rect 302424 318656 302476 318708
rect 324780 318656 324832 318708
rect 329564 318656 329616 318708
rect 298100 318588 298152 318640
rect 303988 318588 304040 318640
rect 314752 318588 314804 318640
rect 329472 318588 329524 318640
rect 290372 318452 290424 318504
rect 290648 318452 290700 318504
rect 291752 318452 291804 318504
rect 291936 318452 291988 318504
rect 332232 318520 332284 318572
rect 297732 318452 297784 318504
rect 301504 318452 301556 318504
rect 302700 318452 302752 318504
rect 303988 318452 304040 318504
rect 304632 318452 304684 318504
rect 309508 318452 309560 318504
rect 310244 318452 310296 318504
rect 317696 318452 317748 318504
rect 324780 318452 324832 318504
rect 269396 318384 269448 318436
rect 269948 318384 270000 318436
rect 270316 318384 270368 318436
rect 284760 318384 284812 318436
rect 271696 318316 271748 318368
rect 286140 318316 286192 318368
rect 242532 318248 242584 318300
rect 278044 318248 278096 318300
rect 288072 318248 288124 318300
rect 281540 318180 281592 318232
rect 282736 318180 282788 318232
rect 238760 318112 238812 318164
rect 213828 318044 213880 318096
rect 271328 318044 271380 318096
rect 271696 318044 271748 318096
rect 281632 318112 281684 318164
rect 289912 318180 289964 318232
rect 282276 318044 282328 318096
rect 275836 317976 275888 318028
rect 295892 318384 295944 318436
rect 296444 318384 296496 318436
rect 297180 318384 297232 318436
rect 291292 318316 291344 318368
rect 291752 318316 291804 318368
rect 333520 318384 333572 318436
rect 291476 318248 291528 318300
rect 292488 318248 292540 318300
rect 332048 318316 332100 318368
rect 297732 318248 297784 318300
rect 328092 318248 328144 318300
rect 328736 318248 328788 318300
rect 359464 318248 359516 318300
rect 315028 318180 315080 318232
rect 328184 318180 328236 318232
rect 328828 318180 328880 318232
rect 360936 318180 360988 318232
rect 290556 318112 290608 318164
rect 291108 318112 291160 318164
rect 297272 318112 297324 318164
rect 299296 318112 299348 318164
rect 300492 318112 300544 318164
rect 304632 318112 304684 318164
rect 304908 318112 304960 318164
rect 309876 318112 309928 318164
rect 310152 318112 310204 318164
rect 322296 318112 322348 318164
rect 324044 318112 324096 318164
rect 328644 318112 328696 318164
rect 364524 318112 364576 318164
rect 292120 318044 292172 318096
rect 292580 318044 292632 318096
rect 317512 318044 317564 318096
rect 323124 318044 323176 318096
rect 331404 318044 331456 318096
rect 331772 318044 331824 318096
rect 332324 318044 332376 318096
rect 388260 318044 388312 318096
rect 303160 317976 303212 318028
rect 305000 317976 305052 318028
rect 328460 317976 328512 318028
rect 354220 317976 354272 318028
rect 259184 317908 259236 317960
rect 288532 317908 288584 317960
rect 294512 317908 294564 317960
rect 295064 317908 295116 317960
rect 302608 317908 302660 317960
rect 307392 317908 307444 317960
rect 309876 317908 309928 317960
rect 310428 317908 310480 317960
rect 325700 317908 325752 317960
rect 326988 317908 327040 317960
rect 328552 317908 328604 317960
rect 338580 317908 338632 317960
rect 268568 317840 268620 317892
rect 282920 317840 282972 317892
rect 286048 317840 286100 317892
rect 331128 317840 331180 317892
rect 298100 317772 298152 317824
rect 302608 317772 302660 317824
rect 303436 317772 303488 317824
rect 303712 317772 303764 317824
rect 305368 317772 305420 317824
rect 306840 317772 306892 317824
rect 318064 317772 318116 317824
rect 327172 317772 327224 317824
rect 327448 317772 327500 317824
rect 275468 317704 275520 317756
rect 276664 317704 276716 317756
rect 282920 317704 282972 317756
rect 283104 317704 283156 317756
rect 249800 317636 249852 317688
rect 286048 317704 286100 317756
rect 287336 317704 287388 317756
rect 288256 317704 288308 317756
rect 284116 317636 284168 317688
rect 290188 317636 290240 317688
rect 290280 317636 290332 317688
rect 291108 317636 291160 317688
rect 291200 317636 291252 317688
rect 292304 317636 292356 317688
rect 334992 317704 335044 317756
rect 293500 317636 293552 317688
rect 294236 317636 294288 317688
rect 297272 317636 297324 317688
rect 332508 317636 332560 317688
rect 269396 317568 269448 317620
rect 293684 317568 293736 317620
rect 295064 317568 295116 317620
rect 296628 317568 296680 317620
rect 296720 317568 296772 317620
rect 298284 317568 298336 317620
rect 303436 317568 303488 317620
rect 304816 317568 304868 317620
rect 304908 317568 304960 317620
rect 306472 317568 306524 317620
rect 307392 317568 307444 317620
rect 313648 317568 313700 317620
rect 286324 317500 286376 317552
rect 290832 317500 290884 317552
rect 291200 317500 291252 317552
rect 291936 317500 291988 317552
rect 320640 317568 320692 317620
rect 324780 317568 324832 317620
rect 325332 317568 325384 317620
rect 326988 317568 327040 317620
rect 333796 317500 333848 317552
rect 274548 317432 274600 317484
rect 276940 317432 276992 317484
rect 287152 317432 287204 317484
rect 291016 317432 291068 317484
rect 291108 317432 291160 317484
rect 306840 317432 306892 317484
rect 309324 317432 309376 317484
rect 310520 317432 310572 317484
rect 313648 317432 313700 317484
rect 325424 317432 325476 317484
rect 327540 317432 327592 317484
rect 328184 317432 328236 317484
rect 328368 317432 328420 317484
rect 329564 317432 329616 317484
rect 280160 317364 280212 317416
rect 280988 317364 281040 317416
rect 284944 317364 284996 317416
rect 289728 317364 289780 317416
rect 290096 317364 290148 317416
rect 295340 317364 295392 317416
rect 320364 317364 320416 317416
rect 331036 317364 331088 317416
rect 334992 317364 335044 317416
rect 338672 317364 338724 317416
rect 280804 317296 280856 317348
rect 297272 317296 297324 317348
rect 303252 317296 303304 317348
rect 308220 317296 308272 317348
rect 316684 317296 316736 317348
rect 332140 317296 332192 317348
rect 278688 317228 278740 317280
rect 308404 317228 308456 317280
rect 315948 317228 316000 317280
rect 375564 317228 375616 317280
rect 376668 317228 376720 317280
rect 265900 317160 265952 317212
rect 286416 317160 286468 317212
rect 295616 317160 295668 317212
rect 296352 317160 296404 317212
rect 296996 317160 297048 317212
rect 330760 317160 330812 317212
rect 331680 317160 331732 317212
rect 389640 317160 389692 317212
rect 209596 317024 209648 317076
rect 266360 317024 266412 317076
rect 201316 316956 201368 317008
rect 260656 316956 260708 317008
rect 283840 317092 283892 317144
rect 284300 317092 284352 317144
rect 284484 317092 284536 317144
rect 295524 317092 295576 317144
rect 350080 317092 350132 317144
rect 274456 317024 274508 317076
rect 303804 317024 303856 317076
rect 328460 317024 328512 317076
rect 270960 316956 271012 317008
rect 209044 316888 209096 316940
rect 280160 316888 280212 316940
rect 308220 316956 308272 317008
rect 316684 316956 316736 317008
rect 317052 316956 317104 317008
rect 328552 316956 328604 317008
rect 310704 316888 310756 316940
rect 324044 316888 324096 316940
rect 219072 316820 219124 316872
rect 294420 316820 294472 316872
rect 297272 316820 297324 316872
rect 302240 316820 302292 316872
rect 303344 316820 303396 316872
rect 314568 316820 314620 316872
rect 327264 316820 327316 316872
rect 341340 316820 341392 316872
rect 215116 316752 215168 316804
rect 295524 316752 295576 316804
rect 317880 316752 317932 316804
rect 345940 316752 345992 316804
rect 378048 316752 378100 316804
rect 295984 316684 296036 316736
rect 309876 316684 309928 316736
rect 360200 316684 360252 316736
rect 376668 316684 376720 316736
rect 429844 316684 429896 316736
rect 212264 316616 212316 316668
rect 296996 316616 297048 316668
rect 314752 316616 314804 316668
rect 315396 316616 315448 316668
rect 322664 316616 322716 316668
rect 393504 316616 393556 316668
rect 308404 316548 308456 316600
rect 329288 316548 329340 316600
rect 329380 316548 329432 316600
rect 336556 316548 336608 316600
rect 303344 316480 303396 316532
rect 329104 316480 329156 316532
rect 284668 316412 284720 316464
rect 285312 316412 285364 316464
rect 324596 316412 324648 316464
rect 392308 316412 392360 316464
rect 294328 316344 294380 316396
rect 294880 316344 294932 316396
rect 295616 316344 295668 316396
rect 295800 316344 295852 316396
rect 315396 316344 315448 316396
rect 315948 316344 316000 316396
rect 329196 316344 329248 316396
rect 336648 316344 336700 316396
rect 284668 316276 284720 316328
rect 285128 316276 285180 316328
rect 287060 316276 287112 316328
rect 287520 316276 287572 316328
rect 287796 316276 287848 316328
rect 287980 316276 288032 316328
rect 292764 316276 292816 316328
rect 299204 316276 299256 316328
rect 331680 316276 331732 316328
rect 332048 316276 332100 316328
rect 282276 316208 282328 316260
rect 300860 316208 300912 316260
rect 301688 316208 301740 316260
rect 302148 316208 302200 316260
rect 302424 316208 302476 316260
rect 303528 316208 303580 316260
rect 305276 316208 305328 316260
rect 305552 316208 305604 316260
rect 312084 316208 312136 316260
rect 312820 316208 312872 316260
rect 323032 316208 323084 316260
rect 323492 316208 323544 316260
rect 276756 316140 276808 316192
rect 303160 316140 303212 316192
rect 303344 316140 303396 316192
rect 307852 316140 307904 316192
rect 308036 316140 308088 316192
rect 320916 316140 320968 316192
rect 321284 316140 321336 316192
rect 322940 316140 322992 316192
rect 324136 316140 324188 316192
rect 271328 316072 271380 316124
rect 303712 316072 303764 316124
rect 303804 316072 303856 316124
rect 304356 316072 304408 316124
rect 317696 316072 317748 316124
rect 318340 316072 318392 316124
rect 323308 316072 323360 316124
rect 324228 316072 324280 316124
rect 325056 316072 325108 316124
rect 325424 316072 325476 316124
rect 325884 316072 325936 316124
rect 326252 316072 326304 316124
rect 360200 316072 360252 316124
rect 361396 316072 361448 316124
rect 217692 316004 217744 316056
rect 292764 316004 292816 316056
rect 294328 316004 294380 316056
rect 295156 316004 295208 316056
rect 297272 316004 297324 316056
rect 297640 316004 297692 316056
rect 299848 316004 299900 316056
rect 300584 316004 300636 316056
rect 301044 316004 301096 316056
rect 302056 316004 302108 316056
rect 302240 316004 302292 316056
rect 302976 316004 303028 316056
rect 305460 316004 305512 316056
rect 305920 316004 305972 316056
rect 306748 316004 306800 316056
rect 307300 316004 307352 316056
rect 308036 316004 308088 316056
rect 308496 316004 308548 316056
rect 308588 316004 308640 316056
rect 308956 316004 309008 316056
rect 310888 316004 310940 316056
rect 311716 316004 311768 316056
rect 315028 316004 315080 316056
rect 315488 316004 315540 316056
rect 316132 316004 316184 316056
rect 316500 316004 316552 316056
rect 317512 316004 317564 316056
rect 318248 316004 318300 316056
rect 320456 316004 320508 316056
rect 321284 316004 321336 316056
rect 321560 316004 321612 316056
rect 322848 316004 322900 316056
rect 323032 316004 323084 316056
rect 323676 316004 323728 316056
rect 324412 316004 324464 316056
rect 325608 316004 325660 316056
rect 325976 316004 326028 316056
rect 326436 316004 326488 316056
rect 274364 315936 274416 315988
rect 278780 315868 278832 315920
rect 279148 315868 279200 315920
rect 270408 315800 270460 315852
rect 214840 315460 214892 315512
rect 268660 315732 268712 315784
rect 285772 315732 285824 315784
rect 286140 315732 286192 315784
rect 286692 315732 286744 315784
rect 287336 315732 287388 315784
rect 287704 315732 287756 315784
rect 287796 315732 287848 315784
rect 288348 315732 288400 315784
rect 289268 315732 289320 315784
rect 289728 315732 289780 315784
rect 290280 315732 290332 315784
rect 290648 315732 290700 315784
rect 291292 315732 291344 315784
rect 291568 315732 291620 315784
rect 294236 315800 294288 315852
rect 295248 315800 295300 315852
rect 295708 315800 295760 315852
rect 296536 315800 296588 315852
rect 297364 315800 297416 315852
rect 297916 315800 297968 315852
rect 298192 315800 298244 315852
rect 299112 315800 299164 315852
rect 300032 315800 300084 315852
rect 300400 315800 300452 315852
rect 301136 315800 301188 315852
rect 301780 315800 301832 315852
rect 294420 315732 294472 315784
rect 298284 315732 298336 315784
rect 299388 315732 299440 315784
rect 299940 315732 299992 315784
rect 300216 315732 300268 315784
rect 268752 315664 268804 315716
rect 263324 315596 263376 315648
rect 284852 315596 284904 315648
rect 286048 315664 286100 315716
rect 286784 315664 286836 315716
rect 287244 315664 287296 315716
rect 287888 315664 287940 315716
rect 291476 315664 291528 315716
rect 292396 315664 292448 315716
rect 296812 315664 296864 315716
rect 297916 315664 297968 315716
rect 287428 315596 287480 315648
rect 288072 315596 288124 315648
rect 291568 315596 291620 315648
rect 292212 315596 292264 315648
rect 293224 315596 293276 315648
rect 293776 315596 293828 315648
rect 291200 315528 291252 315580
rect 306840 315936 306892 315988
rect 307024 315936 307076 315988
rect 308220 315936 308272 315988
rect 309048 315936 309100 315988
rect 309784 315936 309836 315988
rect 310244 315936 310296 315988
rect 310704 315936 310756 315988
rect 311440 315936 311492 315988
rect 311532 315936 311584 315988
rect 311808 315936 311860 315988
rect 312176 315936 312228 315988
rect 312636 315936 312688 315988
rect 314936 315936 314988 315988
rect 315672 315936 315724 315988
rect 316224 315936 316276 315988
rect 316960 315936 317012 315988
rect 317880 315936 317932 315988
rect 318524 315936 318576 315988
rect 304172 315868 304224 315920
rect 304724 315868 304776 315920
rect 306656 315868 306708 315920
rect 307668 315868 307720 315920
rect 308128 315868 308180 315920
rect 308680 315868 308732 315920
rect 315212 315868 315264 315920
rect 315948 315868 316000 315920
rect 305184 315800 305236 315852
rect 305736 315800 305788 315852
rect 307024 315800 307076 315852
rect 307576 315800 307628 315852
rect 309692 315800 309744 315852
rect 310244 315800 310296 315852
rect 314936 315800 314988 315852
rect 315856 315800 315908 315852
rect 306472 315732 306524 315784
rect 307760 315732 307812 315784
rect 313096 315732 313148 315784
rect 313924 315664 313976 315716
rect 314384 315664 314436 315716
rect 317604 315732 317656 315784
rect 318616 315732 318668 315784
rect 320180 315936 320232 315988
rect 320732 315936 320784 315988
rect 341432 315936 341484 315988
rect 361396 315936 361448 315988
rect 366548 315936 366600 315988
rect 320456 315868 320508 315920
rect 372896 315868 372948 315920
rect 319260 315800 319312 315852
rect 372804 315800 372856 315852
rect 374184 315732 374236 315784
rect 320456 315664 320508 315716
rect 320548 315664 320600 315716
rect 321100 315664 321152 315716
rect 321744 315664 321796 315716
rect 322572 315664 322624 315716
rect 324044 315664 324096 315716
rect 344928 315664 344980 315716
rect 303344 315596 303396 315648
rect 328644 315596 328696 315648
rect 310980 315528 311032 315580
rect 316776 315528 316828 315580
rect 338304 315528 338356 315580
rect 354128 315528 354180 315580
rect 276664 315460 276716 315512
rect 293684 315460 293736 315512
rect 293776 315460 293828 315512
rect 306380 315460 306432 315512
rect 314660 315460 314712 315512
rect 348884 315460 348936 315512
rect 374276 315460 374328 315512
rect 214932 315392 214984 315444
rect 270408 315392 270460 315444
rect 273996 315392 274048 315444
rect 294144 315392 294196 315444
rect 295156 315392 295208 315444
rect 309600 315392 309652 315444
rect 316408 315392 316460 315444
rect 351460 315392 351512 315444
rect 383476 315392 383528 315444
rect 209688 315324 209740 315376
rect 268752 315324 268804 315376
rect 285772 315324 285824 315376
rect 292028 315324 292080 315376
rect 293132 315324 293184 315376
rect 293960 315324 294012 315376
rect 312452 315324 312504 315376
rect 347596 315324 347648 315376
rect 384580 315324 384632 315376
rect 216404 315256 216456 315308
rect 278780 315256 278832 315308
rect 292764 315256 292816 315308
rect 293316 315256 293368 315308
rect 313740 315256 313792 315308
rect 328644 315256 328696 315308
rect 382832 315256 382884 315308
rect 398932 315256 398984 315308
rect 278504 315188 278556 315240
rect 320088 315188 320140 315240
rect 325516 315188 325568 315240
rect 333888 315188 333940 315240
rect 312452 315120 312504 315172
rect 313004 315120 313056 315172
rect 313924 315120 313976 315172
rect 379980 315120 380032 315172
rect 280896 315052 280948 315104
rect 319812 315052 319864 315104
rect 324872 315052 324924 315104
rect 325608 315052 325660 315104
rect 300860 314984 300912 315036
rect 328736 314984 328788 315036
rect 313004 314916 313056 314968
rect 319260 314916 319312 314968
rect 324596 314916 324648 314968
rect 325516 314916 325568 314968
rect 208308 314644 208360 314696
rect 267372 314644 267424 314696
rect 271512 314576 271564 314628
rect 278412 314576 278464 314628
rect 284760 314576 284812 314628
rect 285588 314576 285640 314628
rect 304908 314576 304960 314628
rect 340604 314576 340656 314628
rect 284484 314508 284536 314560
rect 285220 314508 285272 314560
rect 299204 314508 299256 314560
rect 337752 314508 337804 314560
rect 277124 314440 277176 314492
rect 280160 314440 280212 314492
rect 318156 314440 318208 314492
rect 318616 314440 318668 314492
rect 384672 314440 384724 314492
rect 319076 314372 319128 314424
rect 320088 314372 320140 314424
rect 380072 314372 380124 314424
rect 285956 314304 286008 314356
rect 286508 314304 286560 314356
rect 316868 314304 316920 314356
rect 376852 314304 376904 314356
rect 288716 314236 288768 314288
rect 289084 314236 289136 314288
rect 318708 314236 318760 314288
rect 378324 314236 378376 314288
rect 280160 314168 280212 314220
rect 293500 314168 293552 314220
rect 296444 314168 296496 314220
rect 356612 314168 356664 314220
rect 282184 314100 282236 314152
rect 304080 314100 304132 314152
rect 363880 314100 363932 314152
rect 271420 314032 271472 314084
rect 295984 314032 296036 314084
rect 311900 314032 311952 314084
rect 312084 314032 312136 314084
rect 319168 314032 319220 314084
rect 319996 314032 320048 314084
rect 379244 314032 379296 314084
rect 216220 313964 216272 314016
rect 292580 313964 292632 314016
rect 300952 313964 301004 314016
rect 301320 313964 301372 314016
rect 351368 313964 351420 314016
rect 220452 313896 220504 313948
rect 314200 313896 314252 313948
rect 322388 313896 322440 313948
rect 322756 313896 322808 313948
rect 324780 313896 324832 313948
rect 330024 313896 330076 313948
rect 337660 313896 337712 313948
rect 378324 313896 378376 313948
rect 466460 313896 466512 313948
rect 300952 313828 301004 313880
rect 301596 313828 301648 313880
rect 310980 313828 311032 313880
rect 329932 313828 329984 313880
rect 312084 313760 312136 313812
rect 312728 313760 312780 313812
rect 318156 313760 318208 313812
rect 318708 313760 318760 313812
rect 317328 313692 317380 313744
rect 386052 313760 386104 313812
rect 322756 313692 322808 313744
rect 389548 313692 389600 313744
rect 329932 313624 329984 313676
rect 330116 313624 330168 313676
rect 293684 313488 293736 313540
rect 300860 313488 300912 313540
rect 275836 313420 275888 313472
rect 293868 313420 293920 313472
rect 327448 313420 327500 313472
rect 328276 313420 328328 313472
rect 215208 313352 215260 313404
rect 298100 313352 298152 313404
rect 212448 313284 212500 313336
rect 293684 313284 293736 313336
rect 293868 313284 293920 313336
rect 299848 313284 299900 313336
rect 311900 313284 311952 313336
rect 319628 313284 319680 313336
rect 263232 313216 263284 313268
rect 287060 313216 287112 313268
rect 308312 313216 308364 313268
rect 309048 313216 309100 313268
rect 309876 313216 309928 313268
rect 310060 313216 310112 313268
rect 277032 313148 277084 313200
rect 278872 313148 278924 313200
rect 307760 313148 307812 313200
rect 327080 313216 327132 313268
rect 327816 313216 327868 313268
rect 330208 313216 330260 313268
rect 333520 313216 333572 313268
rect 333888 313216 333940 313268
rect 340420 313216 340472 313268
rect 534724 313216 534776 313268
rect 579620 313216 579672 313268
rect 309048 313080 309100 313132
rect 329012 313148 329064 313200
rect 311624 313080 311676 313132
rect 371608 313080 371660 313132
rect 317144 313012 317196 313064
rect 377680 313012 377732 313064
rect 303712 312944 303764 312996
rect 365168 312944 365220 312996
rect 310336 312876 310388 312928
rect 370320 312876 370372 312928
rect 298100 312808 298152 312860
rect 298652 312808 298704 312860
rect 358728 312808 358780 312860
rect 209504 312740 209556 312792
rect 263232 312740 263284 312792
rect 210884 312672 210936 312724
rect 265900 312672 265952 312724
rect 277952 312672 278004 312724
rect 294604 312740 294656 312792
rect 342076 312740 342128 312792
rect 303620 312672 303672 312724
rect 350172 312672 350224 312724
rect 205456 312604 205508 312656
rect 288256 312604 288308 312656
rect 309876 312604 309928 312656
rect 328828 312604 328880 312656
rect 334256 312604 334308 312656
rect 390652 312604 390704 312656
rect 219164 312536 219216 312588
rect 310980 312536 311032 312588
rect 320640 312536 320692 312588
rect 321192 312536 321244 312588
rect 323952 312536 324004 312588
rect 330116 312536 330168 312588
rect 389456 312536 389508 312588
rect 300124 312468 300176 312520
rect 343548 312468 343600 312520
rect 319812 312400 319864 312452
rect 320732 312400 320784 312452
rect 320824 312332 320876 312384
rect 321376 312332 321428 312384
rect 392216 312332 392268 312384
rect 498200 312536 498252 312588
rect 322112 312264 322164 312316
rect 388076 312264 388128 312316
rect 313188 312196 313240 312248
rect 323124 312196 323176 312248
rect 278872 311992 278924 312044
rect 309140 311992 309192 312044
rect 282736 311924 282788 311976
rect 319812 311924 319864 311976
rect 278596 311856 278648 311908
rect 320640 311856 320692 311908
rect 202604 311448 202656 311500
rect 259276 311788 259328 311840
rect 288532 311788 288584 311840
rect 312452 311788 312504 311840
rect 313188 311788 313240 311840
rect 313556 311788 313608 311840
rect 314568 311788 314620 311840
rect 375288 311788 375340 311840
rect 263048 311720 263100 311772
rect 263416 311720 263468 311772
rect 288624 311720 288676 311772
rect 310980 311720 311032 311772
rect 311808 311720 311860 311772
rect 371424 311720 371476 311772
rect 297272 311652 297324 311704
rect 356980 311652 357032 311704
rect 294696 311584 294748 311636
rect 300216 311584 300268 311636
rect 313280 311584 313332 311636
rect 313648 311584 313700 311636
rect 373356 311584 373408 311636
rect 298928 311516 298980 311568
rect 358176 311516 358228 311568
rect 289268 311448 289320 311500
rect 302884 311448 302936 311500
rect 361672 311448 361724 311500
rect 208124 311380 208176 311432
rect 270132 311380 270184 311432
rect 297364 311380 297416 311432
rect 355508 311380 355560 311432
rect 200028 311312 200080 311364
rect 263048 311312 263100 311364
rect 267648 311312 267700 311364
rect 271880 311312 271932 311364
rect 286324 311312 286376 311364
rect 286416 311312 286468 311364
rect 309968 311312 310020 311364
rect 362224 311312 362276 311364
rect 214748 311244 214800 311296
rect 281632 311244 281684 311296
rect 283748 311244 283800 311296
rect 313280 311244 313332 311296
rect 323124 311244 323176 311296
rect 371516 311244 371568 311296
rect 211988 311176 212040 311228
rect 284852 311176 284904 311228
rect 295708 311176 295760 311228
rect 295984 311176 296036 311228
rect 339132 311176 339184 311228
rect 204168 311108 204220 311160
rect 284392 311108 284444 311160
rect 293224 311108 293276 311160
rect 333336 311108 333388 311160
rect 308220 311040 308272 311092
rect 342260 311108 342312 311160
rect 343456 311108 343508 311160
rect 296720 310972 296772 311024
rect 297456 310972 297508 311024
rect 331956 310972 332008 311024
rect 310796 310904 310848 310956
rect 311164 310904 311216 310956
rect 340328 310904 340380 310956
rect 212172 310428 212224 310480
rect 298560 310428 298612 310480
rect 299112 310428 299164 310480
rect 313464 310428 313516 310480
rect 314200 310428 314252 310480
rect 374920 310428 374972 310480
rect 375288 310428 375340 310480
rect 287888 310360 287940 310412
rect 303620 310360 303672 310412
rect 312268 310360 312320 310412
rect 312912 310360 312964 310412
rect 373632 310360 373684 310412
rect 296720 310292 296772 310344
rect 282368 310224 282420 310276
rect 298836 310224 298888 310276
rect 282828 310156 282880 310208
rect 291844 310156 291896 310208
rect 265992 310020 266044 310072
rect 273352 310020 273404 310072
rect 287060 310088 287112 310140
rect 279976 310020 280028 310072
rect 296076 310156 296128 310208
rect 355416 310292 355468 310344
rect 317512 310224 317564 310276
rect 318616 310224 318668 310276
rect 376300 310224 376352 310276
rect 299112 310156 299164 310208
rect 356888 310156 356940 310208
rect 294328 310088 294380 310140
rect 294972 310088 295024 310140
rect 344744 310088 344796 310140
rect 298836 310020 298888 310072
rect 301320 310020 301372 310072
rect 222200 309952 222252 310004
rect 282644 309952 282696 310004
rect 283656 309952 283708 310004
rect 302148 309952 302200 310004
rect 347412 310020 347464 310072
rect 308128 309952 308180 310004
rect 354036 309952 354088 310004
rect 265716 309884 265768 309936
rect 332784 309884 332836 309936
rect 260196 309816 260248 309868
rect 332600 309816 332652 309868
rect 291844 309748 291896 309800
rect 298008 309748 298060 309800
rect 341984 309748 342036 309800
rect 375288 309748 375340 309800
rect 414020 309748 414072 309800
rect 305000 309680 305052 309732
rect 305644 309680 305696 309732
rect 347504 309680 347556 309732
rect 298744 309612 298796 309664
rect 300492 309612 300544 309664
rect 333428 309612 333480 309664
rect 321284 309544 321336 309596
rect 346032 309544 346084 309596
rect 328460 309476 328512 309528
rect 328644 309476 328696 309528
rect 296076 309136 296128 309188
rect 307024 309136 307076 309188
rect 307484 309136 307536 309188
rect 270408 309068 270460 309120
rect 292764 309068 292816 309120
rect 302516 309068 302568 309120
rect 303068 309068 303120 309120
rect 277124 308796 277176 308848
rect 303988 309000 304040 309052
rect 334900 309068 334952 309120
rect 306840 309000 306892 309052
rect 307208 309000 307260 309052
rect 309784 309000 309836 309052
rect 337568 309000 337620 309052
rect 307484 308932 307536 308984
rect 368296 308932 368348 308984
rect 307208 308864 307260 308916
rect 366456 308864 366508 308916
rect 305460 308796 305512 308848
rect 306104 308796 306156 308848
rect 363604 308796 363656 308848
rect 293408 308728 293460 308780
rect 310520 308728 310572 308780
rect 365812 308728 365864 308780
rect 300400 308660 300452 308712
rect 305552 308660 305604 308712
rect 360844 308660 360896 308712
rect 303068 308592 303120 308644
rect 352840 308592 352892 308644
rect 296996 308524 297048 308576
rect 339040 308524 339092 308576
rect 213552 308456 213604 308508
rect 269580 308456 269632 308508
rect 270408 308456 270460 308508
rect 302608 308456 302660 308508
rect 343180 308456 343232 308508
rect 221924 308388 221976 308440
rect 301412 308388 301464 308440
rect 303620 308388 303672 308440
rect 364892 308388 364944 308440
rect 286784 308320 286836 308372
rect 327540 308320 327592 308372
rect 296996 308252 297048 308304
rect 297456 308252 297508 308304
rect 307484 308252 307536 308304
rect 367928 308252 367980 308304
rect 315120 308184 315172 308236
rect 315488 308184 315540 308236
rect 389364 308184 389416 308236
rect 284024 307844 284076 307896
rect 308588 307844 308640 307896
rect 308956 307844 309008 307896
rect 210608 307776 210660 307828
rect 296168 307776 296220 307828
rect 304448 307776 304500 307828
rect 306748 307776 306800 307828
rect 307484 307776 307536 307828
rect 261944 307708 261996 307760
rect 287796 307708 287848 307760
rect 298376 307708 298428 307760
rect 299204 307708 299256 307760
rect 299572 307708 299624 307760
rect 300492 307708 300544 307760
rect 301044 307708 301096 307760
rect 301596 307708 301648 307760
rect 304264 307708 304316 307760
rect 305828 307708 305880 307760
rect 314292 307708 314344 307760
rect 394976 307708 395028 307760
rect 395988 307708 396040 307760
rect 280988 307640 281040 307692
rect 301780 307640 301832 307692
rect 360660 307640 360712 307692
rect 260748 307572 260800 307624
rect 283196 307572 283248 307624
rect 303528 307572 303580 307624
rect 304540 307572 304592 307624
rect 301504 307504 301556 307556
rect 302424 307504 302476 307556
rect 363788 307572 363840 307624
rect 320640 307504 320692 307556
rect 381728 307504 381780 307556
rect 299204 307436 299256 307488
rect 356796 307436 356848 307488
rect 274364 307368 274416 307420
rect 302240 307368 302292 307420
rect 312176 307368 312228 307420
rect 370596 307368 370648 307420
rect 275928 307300 275980 307352
rect 303896 307300 303948 307352
rect 358084 307300 358136 307352
rect 300308 307232 300360 307284
rect 301136 307232 301188 307284
rect 301596 307232 301648 307284
rect 344560 307232 344612 307284
rect 202512 307164 202564 307216
rect 261944 307164 261996 307216
rect 300492 307164 300544 307216
rect 341892 307164 341944 307216
rect 217600 307096 217652 307148
rect 300032 307096 300084 307148
rect 209412 307028 209464 307080
rect 297732 307028 297784 307080
rect 305368 307096 305420 307148
rect 345756 307096 345808 307148
rect 301136 307028 301188 307080
rect 336188 307028 336240 307080
rect 395988 307028 396040 307080
rect 409880 307028 409932 307080
rect 329380 306960 329432 307012
rect 332784 306960 332836 307012
rect 302240 306892 302292 306944
rect 338948 306892 339000 306944
rect 336280 306824 336332 306876
rect 280068 306348 280120 306400
rect 303528 306348 303580 306400
rect 266084 306280 266136 306332
rect 285956 306280 286008 306332
rect 297824 306280 297876 306332
rect 359188 306280 359240 306332
rect 291568 306212 291620 306264
rect 351184 306212 351236 306264
rect 295616 306144 295668 306196
rect 355784 306144 355836 306196
rect 294788 306076 294840 306128
rect 352748 306076 352800 306128
rect 295064 306008 295116 306060
rect 348424 306008 348476 306060
rect 294420 305940 294472 305992
rect 347320 305940 347372 305992
rect 210332 305872 210384 305924
rect 266084 305872 266136 305924
rect 217416 305804 217468 305856
rect 291568 305804 291620 305856
rect 217508 305736 217560 305788
rect 295064 305872 295116 305924
rect 296904 305872 296956 305924
rect 349804 305872 349856 305924
rect 214472 305668 214524 305720
rect 294788 305668 294840 305720
rect 214656 305600 214708 305652
rect 304356 305804 304408 305856
rect 316224 305804 316276 305856
rect 316960 305804 317012 305856
rect 319628 305804 319680 305856
rect 372160 305804 372212 305856
rect 296168 305736 296220 305788
rect 336372 305736 336424 305788
rect 300860 305600 300912 305652
rect 340236 305600 340288 305652
rect 285036 305532 285088 305584
rect 327724 305532 327776 305584
rect 287520 305464 287572 305516
rect 330484 305464 330536 305516
rect 316960 305396 317012 305448
rect 353944 305396 353996 305448
rect 263876 305260 263928 305312
rect 264704 305260 264756 305312
rect 291476 305260 291528 305312
rect 292028 305260 292080 305312
rect 330576 305328 330628 305380
rect 209228 305124 209280 305176
rect 267004 305124 267056 305176
rect 205548 305056 205600 305108
rect 265716 305056 265768 305108
rect 204076 304988 204128 305040
rect 263876 304988 263928 305040
rect 287520 304988 287572 305040
rect 287796 304988 287848 305040
rect 291936 304988 291988 305040
rect 295616 304988 295668 305040
rect 297364 304988 297416 305040
rect 297824 304988 297876 305040
rect 299940 304988 299992 305040
rect 300860 304988 300912 305040
rect 285864 304920 285916 304972
rect 317604 304920 317656 304972
rect 330668 304920 330720 304972
rect 281080 304852 281132 304904
rect 294052 304852 294104 304904
rect 354404 304852 354456 304904
rect 303160 304784 303212 304836
rect 314660 304784 314712 304836
rect 315028 304784 315080 304836
rect 319812 304784 319864 304836
rect 381820 304784 381872 304836
rect 311992 304716 312044 304768
rect 373448 304716 373500 304768
rect 301780 304648 301832 304700
rect 310612 304648 310664 304700
rect 370504 304648 370556 304700
rect 295340 304580 295392 304632
rect 295524 304580 295576 304632
rect 355140 304580 355192 304632
rect 282644 304444 282696 304496
rect 294880 304444 294932 304496
rect 341616 304512 341668 304564
rect 288164 304376 288216 304428
rect 296444 304376 296496 304428
rect 334808 304444 334860 304496
rect 309508 304376 309560 304428
rect 343088 304376 343140 304428
rect 294788 304308 294840 304360
rect 311992 304308 312044 304360
rect 314936 304308 314988 304360
rect 315304 304308 315356 304360
rect 347136 304308 347188 304360
rect 286692 304240 286744 304292
rect 317604 304240 317656 304292
rect 320732 304240 320784 304292
rect 321284 304240 321336 304292
rect 314660 304172 314712 304224
rect 387800 304172 387852 304224
rect 309508 303764 309560 303816
rect 309968 303764 310020 303816
rect 270316 303628 270368 303680
rect 313280 303628 313332 303680
rect 269028 303560 269080 303612
rect 287428 303560 287480 303612
rect 303436 303560 303488 303612
rect 369032 303560 369084 303612
rect 365720 303492 365772 303544
rect 286324 303424 286376 303476
rect 301964 303424 302016 303476
rect 302792 303424 302844 303476
rect 364708 303424 364760 303476
rect 299388 303356 299440 303408
rect 359372 303356 359424 303408
rect 288072 303288 288124 303340
rect 300952 303288 301004 303340
rect 307668 303288 307720 303340
rect 331864 303288 331916 303340
rect 288348 303220 288400 303272
rect 300768 303220 300820 303272
rect 360384 303220 360436 303272
rect 298284 303152 298336 303204
rect 356704 303152 356756 303204
rect 279332 303084 279384 303136
rect 299848 303084 299900 303136
rect 334716 303084 334768 303136
rect 299664 303016 299716 303068
rect 352656 303016 352708 303068
rect 205364 302948 205416 303000
rect 269028 302948 269080 303000
rect 301136 302948 301188 303000
rect 349896 302948 349948 303000
rect 220268 302880 220320 302932
rect 298192 302880 298244 302932
rect 299388 302880 299440 302932
rect 300952 302880 301004 302932
rect 348608 302880 348660 302932
rect 395988 302880 396040 302932
rect 565820 302880 565872 302932
rect 299756 302812 299808 302864
rect 341708 302812 341760 302864
rect 303804 302744 303856 302796
rect 304540 302744 304592 302796
rect 337476 302744 337528 302796
rect 321652 302676 321704 302728
rect 322480 302676 322532 302728
rect 383292 302676 383344 302728
rect 213276 302268 213328 302320
rect 259552 302268 259604 302320
rect 260196 302268 260248 302320
rect 202696 302200 202748 302252
rect 262496 302200 262548 302252
rect 262956 302200 263008 302252
rect 299664 302200 299716 302252
rect 300216 302200 300268 302252
rect 302792 302200 302844 302252
rect 303252 302200 303304 302252
rect 264980 302132 265032 302184
rect 266268 302132 266320 302184
rect 287336 302132 287388 302184
rect 321652 302132 321704 302184
rect 394792 302132 394844 302184
rect 296168 302064 296220 302116
rect 296628 302064 296680 302116
rect 358452 302064 358504 302116
rect 300676 301996 300728 302048
rect 360752 301996 360804 302048
rect 300584 301928 300636 301980
rect 359280 301928 359332 301980
rect 312820 301860 312872 301912
rect 313004 301860 313056 301912
rect 372068 301860 372120 301912
rect 293960 301792 294012 301844
rect 294512 301792 294564 301844
rect 351276 301792 351328 301844
rect 295340 301724 295392 301776
rect 295892 301724 295944 301776
rect 352564 301724 352616 301776
rect 262128 301520 262180 301572
rect 275008 301520 275060 301572
rect 286600 301588 286652 301640
rect 288808 301588 288860 301640
rect 289636 301588 289688 301640
rect 344376 301656 344428 301708
rect 297916 301588 297968 301640
rect 348700 301588 348752 301640
rect 283932 301520 283984 301572
rect 293132 301520 293184 301572
rect 207848 301452 207900 301504
rect 264980 301452 265032 301504
rect 299480 301520 299532 301572
rect 300584 301520 300636 301572
rect 348792 301520 348844 301572
rect 321560 301452 321612 301504
rect 322664 301452 322716 301504
rect 381544 301452 381596 301504
rect 336096 301384 336148 301436
rect 255412 301316 255464 301368
rect 256148 301316 256200 301368
rect 263692 301316 263744 301368
rect 264336 301316 264388 301368
rect 197452 300976 197504 301028
rect 255412 300976 255464 301028
rect 202144 300908 202196 300960
rect 261484 300908 261536 300960
rect 204444 300840 204496 300892
rect 263692 300840 263744 300892
rect 255412 300772 255464 300824
rect 255964 300772 256016 300824
rect 262128 300772 262180 300824
rect 286140 300772 286192 300824
rect 291108 300772 291160 300824
rect 367560 300772 367612 300824
rect 265072 300704 265124 300756
rect 265624 300704 265676 300756
rect 306564 300704 306616 300756
rect 307024 300704 307076 300756
rect 305644 300636 305696 300688
rect 307668 300636 307720 300688
rect 303712 300568 303764 300620
rect 304632 300568 304684 300620
rect 336004 300704 336056 300756
rect 307116 300500 307168 300552
rect 307668 300500 307720 300552
rect 369952 300636 370004 300688
rect 314752 300568 314804 300620
rect 315856 300568 315908 300620
rect 376576 300568 376628 300620
rect 311348 300500 311400 300552
rect 367652 300500 367704 300552
rect 283104 300432 283156 300484
rect 341800 300432 341852 300484
rect 302240 300364 302292 300416
rect 362040 300364 362092 300416
rect 305276 300296 305328 300348
rect 305552 300296 305604 300348
rect 345664 300296 345716 300348
rect 304264 300228 304316 300280
rect 343272 300228 343324 300280
rect 205272 300160 205324 300212
rect 262128 300160 262180 300212
rect 307760 300160 307812 300212
rect 344652 300160 344704 300212
rect 193220 300092 193272 300144
rect 254032 300092 254084 300144
rect 286968 300092 287020 300144
rect 303712 300092 303764 300144
rect 305184 300092 305236 300144
rect 306196 300092 306248 300144
rect 338764 300092 338816 300144
rect 308036 300024 308088 300076
rect 336188 300024 336240 300076
rect 307024 299956 307076 300008
rect 311348 299956 311400 300008
rect 306932 299888 306984 299940
rect 333244 299956 333296 300008
rect 309416 299820 309468 299872
rect 374644 299888 374696 299940
rect 216036 299616 216088 299668
rect 259828 299616 259880 299668
rect 260104 299616 260156 299668
rect 204352 299548 204404 299600
rect 265072 299548 265124 299600
rect 194600 299480 194652 299532
rect 255412 299480 255464 299532
rect 4160 299412 4212 299464
rect 221740 299412 221792 299464
rect 256700 299412 256752 299464
rect 257344 299412 257396 299464
rect 288716 299412 288768 299464
rect 289360 299412 289412 299464
rect 316132 299412 316184 299464
rect 316776 299412 316828 299464
rect 378600 299412 378652 299464
rect 288256 299344 288308 299396
rect 348332 299344 348384 299396
rect 316040 299276 316092 299328
rect 316868 299276 316920 299328
rect 376484 299276 376536 299328
rect 289452 299208 289504 299260
rect 348976 299208 349028 299260
rect 289360 299140 289412 299192
rect 347228 299140 347280 299192
rect 287704 299072 287756 299124
rect 290924 299072 290976 299124
rect 345848 299072 345900 299124
rect 284116 299004 284168 299056
rect 290096 299004 290148 299056
rect 344468 299004 344520 299056
rect 207756 298800 207808 298852
rect 290832 298800 290884 298852
rect 338856 298936 338908 298988
rect 311532 298868 311584 298920
rect 349988 298868 350040 298920
rect 336188 298800 336240 298852
rect 369124 298800 369176 298852
rect 233148 298732 233200 298784
rect 580172 298732 580224 298784
rect 218796 298256 218848 298308
rect 264428 298256 264480 298308
rect 193404 298188 193456 298240
rect 253204 298188 253256 298240
rect 193312 298120 193364 298172
rect 253388 298120 253440 298172
rect 244556 298052 244608 298104
rect 245200 298052 245252 298104
rect 250076 298052 250128 298104
rect 250536 298052 250588 298104
rect 283840 298052 283892 298104
rect 284208 298052 284260 298104
rect 288624 298052 288676 298104
rect 289728 298052 289780 298104
rect 291292 298052 291344 298104
rect 292304 298052 292356 298104
rect 293776 298052 293828 298104
rect 366088 298052 366140 298104
rect 305092 297984 305144 298036
rect 305460 297984 305512 298036
rect 368940 297984 368992 298036
rect 309324 297916 309376 297968
rect 310060 297916 310112 297968
rect 319352 297916 319404 297968
rect 319628 297916 319680 297968
rect 382648 297916 382700 297968
rect 373172 297848 373224 297900
rect 308680 297780 308732 297832
rect 369308 297780 369360 297832
rect 307576 297712 307628 297764
rect 367468 297712 367520 297764
rect 289544 297644 289596 297696
rect 306288 297644 306340 297696
rect 364984 297644 365036 297696
rect 263508 297576 263560 297628
rect 264060 297576 264112 297628
rect 303528 297576 303580 297628
rect 363420 297576 363472 297628
rect 283840 297508 283892 297560
rect 337384 297508 337436 297560
rect 230480 297440 230532 297492
rect 242256 297440 242308 297492
rect 292304 297440 292356 297492
rect 342996 297440 343048 297492
rect 203064 297372 203116 297424
rect 263508 297372 263560 297424
rect 271696 297372 271748 297424
rect 315672 297372 315724 297424
rect 335084 297372 335136 297424
rect 307944 297304 307996 297356
rect 348516 297304 348568 297356
rect 178684 297236 178736 297288
rect 234068 297236 234120 297288
rect 187700 297168 187752 297220
rect 245016 297168 245068 297220
rect 202972 297100 203024 297152
rect 262864 297100 262916 297152
rect 176660 297032 176712 297084
rect 236644 297032 236696 297084
rect 293316 297032 293368 297084
rect 293776 297032 293828 297084
rect 195980 296964 196032 297016
rect 256884 296964 256936 297016
rect 173900 296896 173952 296948
rect 235356 296896 235408 296948
rect 189080 296828 189132 296880
rect 250076 296828 250128 296880
rect 183560 296760 183612 296812
rect 244556 296760 244608 296812
rect 203984 296692 204036 296744
rect 288624 296692 288676 296744
rect 305920 296692 305972 296744
rect 306932 296692 306984 296744
rect 287980 296624 288032 296676
rect 346952 296624 347004 296676
rect 236828 296080 236880 296132
rect 245108 296080 245160 296132
rect 169760 296012 169812 296064
rect 230480 296012 230532 296064
rect 210516 295944 210568 295996
rect 235172 295944 235224 295996
rect 212908 295876 212960 295928
rect 240140 296012 240192 296064
rect 264520 296012 264572 296064
rect 213184 295808 213236 295860
rect 243084 295808 243136 295860
rect 272340 295944 272392 295996
rect 213000 295740 213052 295792
rect 248604 295740 248656 295792
rect 249156 295740 249208 295792
rect 176752 295672 176804 295724
rect 236828 295672 236880 295724
rect 173992 295604 174044 295656
rect 233884 295604 233936 295656
rect 171140 295536 171192 295588
rect 232412 295536 232464 295588
rect 172520 295468 172572 295520
rect 233976 295468 234028 295520
rect 190460 295400 190512 295452
rect 251180 295400 251232 295452
rect 297732 295400 297784 295452
rect 305552 295400 305604 295452
rect 230940 295332 230992 295384
rect 231676 295332 231728 295384
rect 233884 295332 233936 295384
rect 234528 295332 234580 295384
rect 577596 295332 577648 295384
rect 288900 295264 288952 295316
rect 347044 295264 347096 295316
rect 288624 295196 288676 295248
rect 342904 295196 342956 295248
rect 287612 295128 287664 295180
rect 340144 295128 340196 295180
rect 291660 295060 291712 295112
rect 344284 295060 344336 295112
rect 167000 294788 167052 294840
rect 228272 294788 228324 294840
rect 242808 294788 242860 294840
rect 272432 294788 272484 294840
rect 168380 294720 168432 294772
rect 229100 294720 229152 294772
rect 229836 294720 229888 294772
rect 235724 294720 235776 294772
rect 267280 294720 267332 294772
rect 222476 294652 222528 294704
rect 283012 294652 283064 294704
rect 164240 294584 164292 294636
rect 224868 294584 224920 294636
rect 237472 294584 237524 294636
rect 275100 294584 275152 294636
rect 213736 294516 213788 294568
rect 232044 294516 232096 294568
rect 233148 294516 233200 294568
rect 171232 294448 171284 294500
rect 231124 294448 231176 294500
rect 165896 294380 165948 294432
rect 225604 294380 225656 294432
rect 169852 294312 169904 294364
rect 229928 294312 229980 294364
rect 230204 294312 230256 294364
rect 287612 294312 287664 294364
rect 288256 294312 288308 294364
rect 182180 294244 182232 294296
rect 242716 294244 242768 294296
rect 176844 294176 176896 294228
rect 237932 294176 237984 294228
rect 165712 294108 165764 294160
rect 226892 294108 226944 294160
rect 225604 294040 225656 294092
rect 225788 294040 225840 294092
rect 216496 293972 216548 294024
rect 241980 293972 242032 294024
rect 242808 293972 242860 294024
rect 226340 293904 226392 293956
rect 229744 293904 229796 293956
rect 198740 293428 198792 293480
rect 253112 293428 253164 293480
rect 237380 293360 237432 293412
rect 275192 293360 275244 293412
rect 164884 293292 164936 293344
rect 225696 293292 225748 293344
rect 236092 293292 236144 293344
rect 278228 293292 278280 293344
rect 157800 293224 157852 293276
rect 226340 293224 226392 293276
rect 235356 293224 235408 293276
rect 278136 293224 278188 293276
rect 188344 293156 188396 293208
rect 237472 293156 237524 293208
rect 238484 293156 238536 293208
rect 172704 293088 172756 293140
rect 233148 293088 233200 293140
rect 164332 293020 164384 293072
rect 224224 293020 224276 293072
rect 224684 293020 224736 293072
rect 254032 293020 254084 293072
rect 254308 293020 254360 293072
rect 259552 293020 259604 293072
rect 260196 293020 260248 293072
rect 262496 293020 262548 293072
rect 263140 293020 263192 293072
rect 263692 293020 263744 293072
rect 264244 293020 264296 293072
rect 179420 292952 179472 293004
rect 239772 292952 239824 293004
rect 263876 292952 263928 293004
rect 264612 292952 264664 293004
rect 176936 292884 176988 292936
rect 237380 292884 237432 292936
rect 172612 292816 172664 292868
rect 232780 292816 232832 292868
rect 175280 292748 175332 292800
rect 236092 292748 236144 292800
rect 236460 292748 236512 292800
rect 216588 292680 216640 292732
rect 235356 292680 235408 292732
rect 210700 292612 210752 292664
rect 3424 292544 3476 292596
rect 198740 292544 198792 292596
rect 219256 292544 219308 292596
rect 228732 292544 228784 292596
rect 235172 292476 235224 292528
rect 236092 292476 236144 292528
rect 237472 292476 237524 292528
rect 238576 292476 238628 292528
rect 239404 292476 239456 292528
rect 242256 292476 242308 292528
rect 261484 292476 261536 292528
rect 262220 292476 262272 292528
rect 264428 292476 264480 292528
rect 264980 292476 265032 292528
rect 311624 292476 311676 292528
rect 376760 292476 376812 292528
rect 378140 292476 378192 292528
rect 240876 292408 240928 292460
rect 275744 292408 275796 292460
rect 218888 292340 218940 292392
rect 255964 292340 256016 292392
rect 246672 292272 246724 292324
rect 267188 292272 267240 292324
rect 240508 292204 240560 292256
rect 264520 292204 264572 292256
rect 245292 292136 245344 292188
rect 269764 292136 269816 292188
rect 221464 292068 221516 292120
rect 237380 292068 237432 292120
rect 252836 292068 252888 292120
rect 279700 292068 279752 292120
rect 307116 292068 307168 292120
rect 311624 292068 311676 292120
rect 220820 292000 220872 292052
rect 237472 292000 237524 292052
rect 244188 292000 244240 292052
rect 273076 292000 273128 292052
rect 218612 291932 218664 291984
rect 220176 291932 220228 291984
rect 254860 291932 254912 291984
rect 218520 291864 218572 291916
rect 222108 291864 222160 291916
rect 224408 291864 224460 291916
rect 237380 291864 237432 291916
rect 238300 291864 238352 291916
rect 275652 291864 275704 291916
rect 215944 291796 215996 291848
rect 221740 291796 221792 291848
rect 258172 291796 258224 291848
rect 271052 291796 271104 291848
rect 272156 291796 272208 291848
rect 272340 291796 272392 291848
rect 334164 291796 334216 291848
rect 219900 291728 219952 291780
rect 249064 291728 249116 291780
rect 251916 291728 251968 291780
rect 264152 291728 264204 291780
rect 217232 291660 217284 291712
rect 229468 291660 229520 291712
rect 230020 291660 230072 291712
rect 232780 291660 232832 291712
rect 275376 291660 275428 291712
rect 221280 291592 221332 291644
rect 241888 291592 241940 291644
rect 255044 291592 255096 291644
rect 272708 291592 272760 291644
rect 221372 291524 221424 291576
rect 243636 291524 243688 291576
rect 253112 291524 253164 291576
rect 258724 291524 258776 291576
rect 271972 291524 272024 291576
rect 272616 291524 272668 291576
rect 220084 291456 220136 291508
rect 244924 291456 244976 291508
rect 256700 291456 256752 291508
rect 259276 291456 259328 291508
rect 220912 291388 220964 291440
rect 246396 291388 246448 291440
rect 263692 291388 263744 291440
rect 272064 291388 272116 291440
rect 272340 291388 272392 291440
rect 219808 291320 219860 291372
rect 247408 291320 247460 291372
rect 262588 291320 262640 291372
rect 270500 291320 270552 291372
rect 271236 291320 271288 291372
rect 217324 291252 217376 291304
rect 227168 291252 227220 291304
rect 227720 291252 227772 291304
rect 234252 291252 234304 291304
rect 244280 291252 244332 291304
rect 246304 291252 246356 291304
rect 246764 291252 246816 291304
rect 246948 291252 247000 291304
rect 249708 291252 249760 291304
rect 256148 291252 256200 291304
rect 257804 291252 257856 291304
rect 261116 291252 261168 291304
rect 270776 291252 270828 291304
rect 271144 291252 271196 291304
rect 227812 291184 227864 291236
rect 229836 291184 229888 291236
rect 245016 291184 245068 291236
rect 247868 291184 247920 291236
rect 259368 291184 259420 291236
rect 260748 291184 260800 291236
rect 261484 291184 261536 291236
rect 271972 291184 272024 291236
rect 239772 291116 239824 291168
rect 279056 291116 279108 291168
rect 325700 291116 325752 291168
rect 327540 291116 327592 291168
rect 233148 291048 233200 291100
rect 268384 291048 268436 291100
rect 169944 290776 169996 290828
rect 230940 290776 230992 290828
rect 173808 290708 173860 290760
rect 220636 290708 220688 290760
rect 227812 290708 227864 290760
rect 168288 290640 168340 290692
rect 220728 290640 220780 290692
rect 243452 290640 243504 290692
rect 277216 290640 277268 290692
rect 200764 290572 200816 290624
rect 259368 290572 259420 290624
rect 194692 290504 194744 290556
rect 255044 290504 255096 290556
rect 191932 290436 191984 290488
rect 252836 290436 252888 290488
rect 327540 290436 327592 290488
rect 394700 290436 394752 290488
rect 569960 290436 570012 290488
rect 182272 290368 182324 290420
rect 243452 290368 243504 290420
rect 221556 290300 221608 290352
rect 254124 290300 254176 290352
rect 221648 290232 221700 290284
rect 256792 290232 256844 290284
rect 257068 290232 257120 290284
rect 220360 290164 220412 290216
rect 259644 290164 259696 290216
rect 197544 290096 197596 290148
rect 257252 290096 257304 290148
rect 257436 290096 257488 290148
rect 196072 290028 196124 290080
rect 255504 290028 255556 290080
rect 256148 290028 256200 290080
rect 201500 289960 201552 290012
rect 261668 289960 261720 290012
rect 221740 289892 221792 289944
rect 240416 289892 240468 289944
rect 178040 289824 178092 289876
rect 238852 289824 238904 289876
rect 219716 289756 219768 289808
rect 223580 289756 223632 289808
rect 244832 289756 244884 289808
rect 246212 289756 246264 289808
rect 300584 289552 300636 289604
rect 306196 289552 306248 289604
rect 242624 289416 242676 289468
rect 174084 289280 174136 289332
rect 218060 289280 218112 289332
rect 180064 289212 180116 289264
rect 235540 289348 235592 289400
rect 183652 289144 183704 289196
rect 244004 289348 244056 289400
rect 245568 289348 245620 289400
rect 184940 289076 184992 289128
rect 274272 288396 274324 288448
rect 269028 287648 269080 287700
rect 319720 287648 319772 287700
rect 349252 286492 349304 286544
rect 350264 286492 350316 286544
rect 169668 286288 169720 286340
rect 219256 286288 219308 286340
rect 310244 286288 310296 286340
rect 349252 286288 349304 286340
rect 310060 285676 310112 285728
rect 310244 285676 310296 285728
rect 268936 285064 268988 285116
rect 315488 284996 315540 285048
rect 185124 284928 185176 284980
rect 220912 284928 220964 284980
rect 268936 284928 268988 284980
rect 326712 284928 326764 284980
rect 180800 283568 180852 283620
rect 220912 283568 220964 283620
rect 269764 283568 269816 283620
rect 325240 283568 325292 283620
rect 183744 282140 183796 282192
rect 220912 282140 220964 282192
rect 179512 280780 179564 280832
rect 220820 280780 220872 280832
rect 271144 280780 271196 280832
rect 291200 280780 291252 280832
rect 178132 279420 178184 279472
rect 220912 279420 220964 279472
rect 271236 279420 271288 279472
rect 291752 279420 291804 279472
rect 186412 273912 186464 273964
rect 219808 273912 219860 273964
rect 322940 273912 322992 273964
rect 324044 273912 324096 273964
rect 531320 273912 531372 273964
rect 189264 272484 189316 272536
rect 219900 272484 219952 272536
rect 315488 272484 315540 272536
rect 348884 272484 348936 272536
rect 416780 272484 416832 272536
rect 194784 271124 194836 271176
rect 218612 271124 218664 271176
rect 289636 271124 289688 271176
rect 318340 271124 318392 271176
rect 196164 269764 196216 269816
rect 218888 269764 218940 269816
rect 323676 268200 323728 268252
rect 324136 268200 324188 268252
rect 323676 267724 323728 267776
rect 523132 267724 523184 267776
rect 3056 266364 3108 266416
rect 14464 266364 14516 266416
rect 269120 265616 269172 265668
rect 322664 265616 322716 265668
rect 311348 262148 311400 262200
rect 311716 262148 311768 262200
rect 275376 261468 275428 261520
rect 307208 261468 307260 261520
rect 311348 260924 311400 260976
rect 374092 260924 374144 260976
rect 318524 260856 318576 260908
rect 463700 260856 463752 260908
rect 312912 259428 312964 259480
rect 396080 259428 396132 259480
rect 310336 258068 310388 258120
rect 357440 258068 357492 258120
rect 269120 257388 269172 257440
rect 290740 257388 290792 257440
rect 269580 257320 269632 257372
rect 318616 257320 318668 257372
rect 459560 257320 459612 257372
rect 273812 256708 273864 256760
rect 274640 256708 274692 256760
rect 312912 256708 312964 256760
rect 313096 256708 313148 256760
rect 389180 256776 389232 256828
rect 318156 256708 318208 256760
rect 318708 256708 318760 256760
rect 456800 256708 456852 256760
rect 311532 255348 311584 255400
rect 371240 255348 371292 255400
rect 316960 255280 317012 255332
rect 445760 255280 445812 255332
rect 284208 254532 284260 254584
rect 308496 254532 308548 254584
rect 3424 253920 3476 253972
rect 199936 253920 199988 253972
rect 312728 253920 312780 253972
rect 313188 253920 313240 253972
rect 391940 253920 391992 253972
rect 213276 253852 213328 253904
rect 270408 253308 270460 253360
rect 292488 253308 292540 253360
rect 289728 253240 289780 253292
rect 322388 253240 322440 253292
rect 286876 253172 286928 253224
rect 311440 253172 311492 253224
rect 312820 253172 312872 253224
rect 347596 253172 347648 253224
rect 385040 253172 385092 253224
rect 319720 253036 319772 253088
rect 319996 253036 320048 253088
rect 319720 252628 319772 252680
rect 471244 252628 471296 252680
rect 321468 252560 321520 252612
rect 491300 252560 491352 252612
rect 316776 251812 316828 251864
rect 351460 251812 351512 251864
rect 434720 251812 434772 251864
rect 313004 251268 313056 251320
rect 382280 251268 382332 251320
rect 323768 251200 323820 251252
rect 324228 251200 324280 251252
rect 538220 251200 538272 251252
rect 319812 251132 319864 251184
rect 320088 251132 320140 251184
rect 309048 250452 309100 250504
rect 332600 250452 332652 250504
rect 319812 249772 319864 249824
rect 470600 249772 470652 249824
rect 314568 248548 314620 248600
rect 407120 248548 407172 248600
rect 316040 248480 316092 248532
rect 317144 248480 317196 248532
rect 441620 248480 441672 248532
rect 320088 248412 320140 248464
rect 484400 248412 484452 248464
rect 271052 247868 271104 247920
rect 319904 247868 319956 247920
rect 275744 247800 275796 247852
rect 303252 247800 303304 247852
rect 307668 247800 307720 247852
rect 317420 247800 317472 247852
rect 272248 247732 272300 247784
rect 316040 247732 316092 247784
rect 168564 247664 168616 247716
rect 217232 247664 217284 247716
rect 318248 247664 318300 247716
rect 345940 247664 345992 247716
rect 452660 247664 452712 247716
rect 315396 247052 315448 247104
rect 315856 247052 315908 247104
rect 423772 247052 423824 247104
rect 269764 246372 269816 246424
rect 292212 246372 292264 246424
rect 198832 246304 198884 246356
rect 215944 246304 215996 246356
rect 288992 246304 289044 246356
rect 315304 246304 315356 246356
rect 270868 245692 270920 245744
rect 271512 245692 271564 245744
rect 316684 245624 316736 245676
rect 317236 245624 317288 245676
rect 438860 245624 438912 245676
rect 577596 245556 577648 245608
rect 579620 245556 579672 245608
rect 268936 244944 268988 244996
rect 271236 244944 271288 244996
rect 167092 244876 167144 244928
rect 217324 244876 217376 244928
rect 283472 244876 283524 244928
rect 304540 244876 304592 244928
rect 317328 244468 317380 244520
rect 448520 244468 448572 244520
rect 322388 244400 322440 244452
rect 322848 244400 322900 244452
rect 516140 244400 516192 244452
rect 325148 244332 325200 244384
rect 325516 244332 325568 244384
rect 540980 244332 541032 244384
rect 316868 244264 316920 244316
rect 317328 244264 317380 244316
rect 326344 244264 326396 244316
rect 326988 244264 327040 244316
rect 558920 244264 558972 244316
rect 206468 243584 206520 243636
rect 206652 243584 206704 243636
rect 271788 243516 271840 243568
rect 285036 243516 285088 243568
rect 315304 243040 315356 243092
rect 315948 243040 316000 243092
rect 420920 243040 420972 243092
rect 325056 242972 325108 243024
rect 325608 242972 325660 243024
rect 543004 242972 543056 243024
rect 326252 242904 326304 242956
rect 326896 242904 326948 242956
rect 563060 242904 563112 242956
rect 321468 242836 321520 242888
rect 322296 242836 322348 242888
rect 276204 242292 276256 242344
rect 320916 242292 320968 242344
rect 187884 242224 187936 242276
rect 219992 242224 220044 242276
rect 278780 242224 278832 242276
rect 326252 242224 326304 242276
rect 154396 242156 154448 242208
rect 277860 242156 277912 242208
rect 324964 242156 325016 242208
rect 211988 242020 212040 242072
rect 221096 242020 221148 242072
rect 221188 242020 221240 242072
rect 222476 242020 222528 242072
rect 269028 241612 269080 241664
rect 271144 241612 271196 241664
rect 160008 241544 160060 241596
rect 204904 241544 204956 241596
rect 154488 241476 154540 241528
rect 209044 241476 209096 241528
rect 277400 241476 277452 241528
rect 321468 241476 321520 241528
rect 215760 241408 215812 241460
rect 216312 241408 216364 241460
rect 288440 241408 288492 241460
rect 289636 241408 289688 241460
rect 267556 241340 267608 241392
rect 271144 241340 271196 241392
rect 270592 241272 270644 241324
rect 270960 241272 271012 241324
rect 217600 241204 217652 241256
rect 210424 241136 210476 241188
rect 217692 241136 217744 241188
rect 212264 241000 212316 241052
rect 214932 240864 214984 240916
rect 153108 240796 153160 240848
rect 207756 240796 207808 240848
rect 218612 240796 218664 240848
rect 14464 240728 14516 240780
rect 199384 240728 199436 240780
rect 213368 240388 213420 240440
rect 220544 240592 220596 240644
rect 219164 240456 219216 240508
rect 222200 240456 222252 240508
rect 214840 240320 214892 240372
rect 221096 240320 221148 240372
rect 222200 240320 222252 240372
rect 222292 240320 222344 240372
rect 218612 240252 218664 240304
rect 199936 240184 199988 240236
rect 200304 240184 200356 240236
rect 221372 240184 221424 240236
rect 155684 240116 155736 240168
rect 218704 240116 218756 240168
rect 222200 240116 222252 240168
rect 221280 240048 221332 240100
rect 221464 239980 221516 240032
rect 218704 239912 218756 239964
rect 223074 239912 223126 239964
rect 223350 239912 223402 239964
rect 223718 239912 223770 239964
rect 223902 239912 223954 239964
rect 224086 239912 224138 239964
rect 224178 239912 224230 239964
rect 224546 239912 224598 239964
rect 224822 239912 224874 239964
rect 222292 239844 222344 239896
rect 222798 239844 222850 239896
rect 222890 239844 222942 239896
rect 223166 239844 223218 239896
rect 214564 239776 214616 239828
rect 217600 239776 217652 239828
rect 221096 239776 221148 239828
rect 222706 239776 222758 239828
rect 213092 239708 213144 239760
rect 156512 239640 156564 239692
rect 219992 239640 220044 239692
rect 220084 239640 220136 239692
rect 222752 239640 222804 239692
rect 185216 239572 185268 239624
rect 222292 239572 222344 239624
rect 223120 239640 223172 239692
rect 223212 239572 223264 239624
rect 223442 239844 223494 239896
rect 223626 239844 223678 239896
rect 223672 239708 223724 239760
rect 224270 239844 224322 239896
rect 224132 239776 224184 239828
rect 223948 239708 224000 239760
rect 224224 239708 224276 239760
rect 223856 239640 223908 239692
rect 224040 239640 224092 239692
rect 225282 239912 225334 239964
rect 225466 239912 225518 239964
rect 225558 239912 225610 239964
rect 224684 239640 224736 239692
rect 224868 239640 224920 239692
rect 225742 239912 225794 239964
rect 225834 239912 225886 239964
rect 226018 239912 226070 239964
rect 226294 239912 226346 239964
rect 223488 239572 223540 239624
rect 223580 239572 223632 239624
rect 224316 239572 224368 239624
rect 158444 239504 158496 239556
rect 215024 239504 215076 239556
rect 218888 239504 218940 239556
rect 219072 239504 219124 239556
rect 220636 239504 220688 239556
rect 220728 239504 220780 239556
rect 222752 239504 222804 239556
rect 223856 239504 223908 239556
rect 225052 239504 225104 239556
rect 225236 239572 225288 239624
rect 225788 239572 225840 239624
rect 225512 239504 225564 239556
rect 225696 239504 225748 239556
rect 226478 239844 226530 239896
rect 226846 239912 226898 239964
rect 226662 239844 226714 239896
rect 226432 239708 226484 239760
rect 226570 239708 226622 239760
rect 158536 239436 158588 239488
rect 216312 239436 216364 239488
rect 218612 239436 218664 239488
rect 218704 239436 218756 239488
rect 219348 239436 219400 239488
rect 220912 239436 220964 239488
rect 227398 239912 227450 239964
rect 227582 239912 227634 239964
rect 227950 239912 228002 239964
rect 228042 239912 228094 239964
rect 227444 239640 227496 239692
rect 226984 239572 227036 239624
rect 228226 239912 228278 239964
rect 228088 239640 228140 239692
rect 227628 239572 227680 239624
rect 227076 239436 227128 239488
rect 227444 239436 227496 239488
rect 228410 239912 228462 239964
rect 228502 239912 228554 239964
rect 228594 239844 228646 239896
rect 228686 239844 228738 239896
rect 228778 239844 228830 239896
rect 228640 239708 228692 239760
rect 228364 239504 228416 239556
rect 228088 239436 228140 239488
rect 228548 239572 228600 239624
rect 3332 239368 3384 239420
rect 198924 239368 198976 239420
rect 216036 239368 216088 239420
rect 217416 239368 217468 239420
rect 217600 239368 217652 239420
rect 213644 239300 213696 239352
rect 217876 239300 217928 239352
rect 226432 239368 226484 239420
rect 227904 239368 227956 239420
rect 228640 239436 228692 239488
rect 229054 239912 229106 239964
rect 229146 239912 229198 239964
rect 229422 239912 229474 239964
rect 229514 239912 229566 239964
rect 229606 239912 229658 239964
rect 229974 239912 230026 239964
rect 230250 239912 230302 239964
rect 230526 239912 230578 239964
rect 231262 239912 231314 239964
rect 229100 239708 229152 239760
rect 229468 239776 229520 239828
rect 229192 239640 229244 239692
rect 229284 239640 229336 239692
rect 229882 239844 229934 239896
rect 229744 239708 229796 239760
rect 229836 239640 229888 239692
rect 229928 239640 229980 239692
rect 230802 239844 230854 239896
rect 230894 239844 230946 239896
rect 230986 239844 231038 239896
rect 231078 239844 231130 239896
rect 230388 239708 230440 239760
rect 230848 239708 230900 239760
rect 229652 239572 229704 239624
rect 230296 239572 230348 239624
rect 229284 239504 229336 239556
rect 230204 239504 230256 239556
rect 230848 239572 230900 239624
rect 231216 239708 231268 239760
rect 231446 239912 231498 239964
rect 231538 239912 231590 239964
rect 231722 239912 231774 239964
rect 231308 239640 231360 239692
rect 231124 239572 231176 239624
rect 231492 239572 231544 239624
rect 231998 239912 232050 239964
rect 232090 239912 232142 239964
rect 232274 239912 232326 239964
rect 232366 239912 232418 239964
rect 232734 239912 232786 239964
rect 232826 239912 232878 239964
rect 232044 239776 232096 239828
rect 232320 239776 232372 239828
rect 232136 239708 232188 239760
rect 231768 239572 231820 239624
rect 232596 239572 232648 239624
rect 230664 239504 230716 239556
rect 230296 239436 230348 239488
rect 231860 239436 231912 239488
rect 267556 241136 267608 241188
rect 233102 239912 233154 239964
rect 233378 239912 233430 239964
rect 233470 239912 233522 239964
rect 233654 239912 233706 239964
rect 233746 239912 233798 239964
rect 234022 239912 234074 239964
rect 234206 239912 234258 239964
rect 234574 239912 234626 239964
rect 233424 239776 233476 239828
rect 233930 239844 233982 239896
rect 233700 239776 233752 239828
rect 234390 239844 234442 239896
rect 234252 239708 234304 239760
rect 233976 239640 234028 239692
rect 234344 239640 234396 239692
rect 233056 239572 233108 239624
rect 233240 239572 233292 239624
rect 234160 239572 234212 239624
rect 234436 239572 234488 239624
rect 234758 239912 234810 239964
rect 235034 239912 235086 239964
rect 235218 239912 235270 239964
rect 235402 239912 235454 239964
rect 235586 239912 235638 239964
rect 235678 239912 235730 239964
rect 235770 239912 235822 239964
rect 235954 239912 236006 239964
rect 234896 239572 234948 239624
rect 233424 239504 233476 239556
rect 235264 239708 235316 239760
rect 235448 239640 235500 239692
rect 235172 239572 235224 239624
rect 235540 239504 235592 239556
rect 236046 239844 236098 239896
rect 236000 239708 236052 239760
rect 236092 239572 236144 239624
rect 236598 239912 236650 239964
rect 236690 239844 236742 239896
rect 236000 239436 236052 239488
rect 228732 239368 228784 239420
rect 229008 239368 229060 239420
rect 229100 239368 229152 239420
rect 233424 239368 233476 239420
rect 233792 239368 233844 239420
rect 235540 239368 235592 239420
rect 235724 239368 235776 239420
rect 236460 239504 236512 239556
rect 222016 239300 222068 239352
rect 223396 239300 223448 239352
rect 232780 239300 232832 239352
rect 236874 239912 236926 239964
rect 237058 239912 237110 239964
rect 237012 239776 237064 239828
rect 236920 239708 236972 239760
rect 236828 239572 236880 239624
rect 236920 239572 236972 239624
rect 237012 239504 237064 239556
rect 237426 239912 237478 239964
rect 237518 239912 237570 239964
rect 237794 239912 237846 239964
rect 238162 239912 238214 239964
rect 238254 239912 238306 239964
rect 238438 239912 238490 239964
rect 238622 239912 238674 239964
rect 237610 239844 237662 239896
rect 237564 239640 237616 239692
rect 237472 239572 237524 239624
rect 237886 239844 237938 239896
rect 237978 239844 238030 239896
rect 237932 239640 237984 239692
rect 238024 239640 238076 239692
rect 237840 239572 237892 239624
rect 237012 239300 237064 239352
rect 237656 239504 237708 239556
rect 238300 239640 238352 239692
rect 238116 239436 238168 239488
rect 237288 239368 237340 239420
rect 237380 239300 237432 239352
rect 238300 239300 238352 239352
rect 238530 239844 238582 239896
rect 238714 239844 238766 239896
rect 238484 239708 238536 239760
rect 238668 239640 238720 239692
rect 238576 239572 238628 239624
rect 239266 239912 239318 239964
rect 239358 239912 239410 239964
rect 239450 239912 239502 239964
rect 239818 239912 239870 239964
rect 240002 239912 240054 239964
rect 240186 239912 240238 239964
rect 240462 239912 240514 239964
rect 240738 239912 240790 239964
rect 240922 239912 240974 239964
rect 241014 239912 241066 239964
rect 239082 239844 239134 239896
rect 239220 239776 239272 239828
rect 239312 239708 239364 239760
rect 239220 239640 239272 239692
rect 239588 239572 239640 239624
rect 238944 239436 238996 239488
rect 239312 239436 239364 239488
rect 240646 239844 240698 239896
rect 240324 239708 240376 239760
rect 240968 239776 241020 239828
rect 240784 239708 240836 239760
rect 240876 239708 240928 239760
rect 241474 239912 241526 239964
rect 241566 239912 241618 239964
rect 241658 239912 241710 239964
rect 241750 239912 241802 239964
rect 241934 239912 241986 239964
rect 242302 239912 242354 239964
rect 242394 239912 242446 239964
rect 242486 239912 242538 239964
rect 242854 239912 242906 239964
rect 243038 239912 243090 239964
rect 243314 239912 243366 239964
rect 243498 239912 243550 239964
rect 244142 239912 244194 239964
rect 241290 239844 241342 239896
rect 240048 239640 240100 239692
rect 240692 239640 240744 239692
rect 241244 239640 241296 239692
rect 240600 239436 240652 239488
rect 241796 239708 241848 239760
rect 241520 239640 241572 239692
rect 241612 239640 241664 239692
rect 241980 239504 242032 239556
rect 238760 239368 238812 239420
rect 242348 239504 242400 239556
rect 243176 239640 243228 239692
rect 243268 239572 243320 239624
rect 242808 239504 242860 239556
rect 242900 239504 242952 239556
rect 243682 239844 243734 239896
rect 243636 239708 243688 239760
rect 244418 239912 244470 239964
rect 244602 239912 244654 239964
rect 244694 239912 244746 239964
rect 244786 239912 244838 239964
rect 245062 239912 245114 239964
rect 242440 239436 242492 239488
rect 244004 239436 244056 239488
rect 242716 239368 242768 239420
rect 242992 239368 243044 239420
rect 238668 239300 238720 239352
rect 239036 239300 239088 239352
rect 218980 239232 219032 239284
rect 241520 239300 241572 239352
rect 243268 239300 243320 239352
rect 244556 239708 244608 239760
rect 244740 239776 244792 239828
rect 244970 239776 245022 239828
rect 269212 241068 269264 241120
rect 245338 239912 245390 239964
rect 245430 239912 245482 239964
rect 245706 239912 245758 239964
rect 245982 239912 246034 239964
rect 246166 239912 246218 239964
rect 244648 239640 244700 239692
rect 244924 239640 244976 239692
rect 245292 239572 245344 239624
rect 245798 239844 245850 239896
rect 245752 239708 245804 239760
rect 245844 239708 245896 239760
rect 246120 239708 246172 239760
rect 246626 239912 246678 239964
rect 246718 239912 246770 239964
rect 247362 239912 247414 239964
rect 247730 239912 247782 239964
rect 247822 239912 247874 239964
rect 247914 239912 247966 239964
rect 248282 239912 248334 239964
rect 248466 239912 248518 239964
rect 246442 239844 246494 239896
rect 246396 239708 246448 239760
rect 246304 239640 246356 239692
rect 245476 239572 245528 239624
rect 245384 239504 245436 239556
rect 246488 239504 246540 239556
rect 246396 239436 246448 239488
rect 246948 239368 247000 239420
rect 247638 239844 247690 239896
rect 247500 239504 247552 239556
rect 247684 239504 247736 239556
rect 248006 239844 248058 239896
rect 248098 239844 248150 239896
rect 247914 239708 247966 239760
rect 248834 239912 248886 239964
rect 249202 239912 249254 239964
rect 249386 239912 249438 239964
rect 249938 239912 249990 239964
rect 248926 239844 248978 239896
rect 249018 239844 249070 239896
rect 249064 239708 249116 239760
rect 248144 239640 248196 239692
rect 248328 239640 248380 239692
rect 248604 239640 248656 239692
rect 248880 239640 248932 239692
rect 248972 239640 249024 239692
rect 247960 239572 248012 239624
rect 249340 239640 249392 239692
rect 249570 239844 249622 239896
rect 249662 239844 249714 239896
rect 249846 239844 249898 239896
rect 247868 239504 247920 239556
rect 249340 239504 249392 239556
rect 248696 239436 248748 239488
rect 249800 239708 249852 239760
rect 249892 239708 249944 239760
rect 249708 239504 249760 239556
rect 249616 239436 249668 239488
rect 250582 239912 250634 239964
rect 250674 239912 250726 239964
rect 251226 239912 251278 239964
rect 251318 239912 251370 239964
rect 251410 239912 251462 239964
rect 251502 239912 251554 239964
rect 251686 239912 251738 239964
rect 251778 239912 251830 239964
rect 251870 239912 251922 239964
rect 251042 239844 251094 239896
rect 250720 239708 250772 239760
rect 250996 239572 251048 239624
rect 250536 239504 250588 239556
rect 251272 239572 251324 239624
rect 251180 239436 251232 239488
rect 248788 239368 248840 239420
rect 249064 239368 249116 239420
rect 249248 239368 249300 239420
rect 250168 239368 250220 239420
rect 250812 239368 250864 239420
rect 251548 239708 251600 239760
rect 251732 239776 251784 239828
rect 251824 239708 251876 239760
rect 252054 239844 252106 239896
rect 251916 239572 251968 239624
rect 251640 239504 251692 239556
rect 251824 239504 251876 239556
rect 252008 239436 252060 239488
rect 252238 239912 252290 239964
rect 252422 239844 252474 239896
rect 252376 239708 252428 239760
rect 252698 239912 252750 239964
rect 252882 239912 252934 239964
rect 252974 239912 253026 239964
rect 253250 239912 253302 239964
rect 252836 239640 252888 239692
rect 252744 239572 252796 239624
rect 252560 239504 252612 239556
rect 252928 239436 252980 239488
rect 245108 239300 245160 239352
rect 247040 239300 247092 239352
rect 251548 239300 251600 239352
rect 252560 239300 252612 239352
rect 253526 239844 253578 239896
rect 253618 239844 253670 239896
rect 253572 239708 253624 239760
rect 253388 239572 253440 239624
rect 253894 239912 253946 239964
rect 254262 239912 254314 239964
rect 254170 239844 254222 239896
rect 253848 239504 253900 239556
rect 254538 239912 254590 239964
rect 254400 239708 254452 239760
rect 272248 241000 272300 241052
rect 273444 241000 273496 241052
rect 274456 241000 274508 241052
rect 267556 240932 267608 240984
rect 270684 240932 270736 240984
rect 283012 240932 283064 240984
rect 308404 240932 308456 240984
rect 267464 240864 267516 240916
rect 267740 240864 267792 240916
rect 268844 240796 268896 240848
rect 271604 240864 271656 240916
rect 278136 240864 278188 240916
rect 306104 240864 306156 240916
rect 254676 239640 254728 239692
rect 254308 239436 254360 239488
rect 254032 239368 254084 239420
rect 255182 239912 255234 239964
rect 255458 239912 255510 239964
rect 255826 239912 255878 239964
rect 256378 239912 256430 239964
rect 256654 239912 256706 239964
rect 256746 239912 256798 239964
rect 256838 239912 256890 239964
rect 257114 239912 257166 239964
rect 257482 239912 257534 239964
rect 257758 239912 257810 239964
rect 257942 239912 257994 239964
rect 254998 239844 255050 239896
rect 255136 239776 255188 239828
rect 255642 239844 255694 239896
rect 255320 239572 255372 239624
rect 253848 239300 253900 239352
rect 254952 239300 255004 239352
rect 255596 239640 255648 239692
rect 255688 239640 255740 239692
rect 256010 239844 256062 239896
rect 256056 239708 256108 239760
rect 255964 239640 256016 239692
rect 257022 239844 257074 239896
rect 256700 239776 256752 239828
rect 256792 239776 256844 239828
rect 256240 239504 256292 239556
rect 257390 239844 257442 239896
rect 258034 239844 258086 239896
rect 257896 239708 257948 239760
rect 257436 239640 257488 239692
rect 257620 239640 257672 239692
rect 257068 239572 257120 239624
rect 257252 239572 257304 239624
rect 258402 239912 258454 239964
rect 258770 239912 258822 239964
rect 258862 239912 258914 239964
rect 259138 239912 259190 239964
rect 258310 239844 258362 239896
rect 258172 239572 258224 239624
rect 257712 239504 257764 239556
rect 257988 239504 258040 239556
rect 258586 239844 258638 239896
rect 258678 239844 258730 239896
rect 258540 239640 258592 239692
rect 258724 239708 258776 239760
rect 258724 239572 258776 239624
rect 259046 239844 259098 239896
rect 259000 239708 259052 239760
rect 259414 239844 259466 239896
rect 259506 239844 259558 239896
rect 259690 239912 259742 239964
rect 259874 239912 259926 239964
rect 259966 239912 260018 239964
rect 260150 239912 260202 239964
rect 259460 239708 259512 239760
rect 259092 239572 259144 239624
rect 259368 239572 259420 239624
rect 259552 239572 259604 239624
rect 256792 239436 256844 239488
rect 258356 239436 258408 239488
rect 260012 239640 260064 239692
rect 260426 239912 260478 239964
rect 260610 239844 260662 239896
rect 260472 239708 260524 239760
rect 260012 239504 260064 239556
rect 260288 239436 260340 239488
rect 258448 239368 258500 239420
rect 259644 239368 259696 239420
rect 260656 239572 260708 239624
rect 260886 239912 260938 239964
rect 261162 239912 261214 239964
rect 261254 239912 261306 239964
rect 269488 240796 269540 240848
rect 271144 240796 271196 240848
rect 287704 240796 287756 240848
rect 287980 240796 288032 240848
rect 312544 240796 312596 240848
rect 269212 240728 269264 240780
rect 299204 240728 299256 240780
rect 261024 239640 261076 239692
rect 261300 239572 261352 239624
rect 269120 240660 269172 240712
rect 274732 240660 274784 240712
rect 269580 240592 269632 240644
rect 267924 240524 267976 240576
rect 269212 240524 269264 240576
rect 278780 240524 278832 240576
rect 278964 240524 279016 240576
rect 261806 239912 261858 239964
rect 261990 239912 262042 239964
rect 262174 239912 262226 239964
rect 261622 239844 261674 239896
rect 262358 239844 262410 239896
rect 262312 239708 262364 239760
rect 261852 239640 261904 239692
rect 261668 239572 261720 239624
rect 262726 239912 262778 239964
rect 270132 240456 270184 240508
rect 287796 240456 287848 240508
rect 287980 240456 288032 240508
rect 268292 240388 268344 240440
rect 268200 240320 268252 240372
rect 268844 240320 268896 240372
rect 283012 240320 283064 240372
rect 262910 239912 262962 239964
rect 263002 239912 263054 239964
rect 263094 239912 263146 239964
rect 263278 239912 263330 239964
rect 263462 239912 263514 239964
rect 262542 239844 262594 239896
rect 262956 239776 263008 239828
rect 263048 239776 263100 239828
rect 263416 239708 263468 239760
rect 263738 239912 263790 239964
rect 264014 239912 264066 239964
rect 263830 239844 263882 239896
rect 263876 239708 263928 239760
rect 263140 239640 263192 239692
rect 263600 239640 263652 239692
rect 263784 239640 263836 239692
rect 264382 239912 264434 239964
rect 267924 240252 267976 240304
rect 288440 240252 288492 240304
rect 270132 240184 270184 240236
rect 270684 240184 270736 240236
rect 278136 240184 278188 240236
rect 269488 240116 269540 240168
rect 267556 240048 267608 240100
rect 268200 240048 268252 240100
rect 285772 240048 285824 240100
rect 286784 240048 286836 240100
rect 264842 239912 264894 239964
rect 264934 239912 264986 239964
rect 265578 239912 265630 239964
rect 265670 239912 265722 239964
rect 266774 239912 266826 239964
rect 264796 239640 264848 239692
rect 264060 239572 264112 239624
rect 264152 239572 264204 239624
rect 264520 239572 264572 239624
rect 265118 239844 265170 239896
rect 265486 239844 265538 239896
rect 265624 239776 265676 239828
rect 265532 239708 265584 239760
rect 266038 239844 266090 239896
rect 266222 239844 266274 239896
rect 265440 239640 265492 239692
rect 265900 239572 265952 239624
rect 261024 239436 261076 239488
rect 261208 239436 261260 239488
rect 262128 239504 262180 239556
rect 262496 239504 262548 239556
rect 267050 239912 267102 239964
rect 267234 239912 267286 239964
rect 268108 239912 268160 239964
rect 267740 239776 267792 239828
rect 299112 239776 299164 239828
rect 267096 239708 267148 239760
rect 267188 239708 267240 239760
rect 268476 239708 268528 239760
rect 271236 239708 271288 239760
rect 293592 239708 293644 239760
rect 268016 239640 268068 239692
rect 266958 239572 267010 239624
rect 270868 239572 270920 239624
rect 262588 239436 262640 239488
rect 269212 239504 269264 239556
rect 263140 239368 263192 239420
rect 263600 239368 263652 239420
rect 264704 239368 264756 239420
rect 265900 239368 265952 239420
rect 259736 239300 259788 239352
rect 260288 239300 260340 239352
rect 264888 239300 264940 239352
rect 267188 239436 267240 239488
rect 267280 239436 267332 239488
rect 267740 239436 267792 239488
rect 268752 239436 268804 239488
rect 266636 239368 266688 239420
rect 267556 239368 267608 239420
rect 269488 239368 269540 239420
rect 278688 239640 278740 239692
rect 271512 239572 271564 239624
rect 297824 239572 297876 239624
rect 273260 239504 273312 239556
rect 311256 239504 311308 239556
rect 271604 239436 271656 239488
rect 320824 239436 320876 239488
rect 274272 239368 274324 239420
rect 293868 239368 293920 239420
rect 527180 239368 527232 239420
rect 269948 239300 270000 239352
rect 270684 239300 270736 239352
rect 285772 239300 285824 239352
rect 241428 239232 241480 239284
rect 269396 239232 269448 239284
rect 214748 239164 214800 239216
rect 221096 239164 221148 239216
rect 223396 239164 223448 239216
rect 223488 239164 223540 239216
rect 223856 239164 223908 239216
rect 224960 239164 225012 239216
rect 225696 239164 225748 239216
rect 227904 239164 227956 239216
rect 228180 239164 228232 239216
rect 233424 239164 233476 239216
rect 241152 239164 241204 239216
rect 245660 239164 245712 239216
rect 270040 239164 270092 239216
rect 215760 239096 215812 239148
rect 225972 239096 226024 239148
rect 221188 239028 221240 239080
rect 223120 239028 223172 239080
rect 228088 239028 228140 239080
rect 228824 239028 228876 239080
rect 211988 238960 212040 239012
rect 212264 238960 212316 239012
rect 213276 238960 213328 239012
rect 236184 239096 236236 239148
rect 236920 239096 236972 239148
rect 237840 239096 237892 239148
rect 238116 239096 238168 239148
rect 238576 239096 238628 239148
rect 229836 239028 229888 239080
rect 242256 239096 242308 239148
rect 242532 239096 242584 239148
rect 246304 239096 246356 239148
rect 247776 239096 247828 239148
rect 269856 239096 269908 239148
rect 229468 238960 229520 239012
rect 154304 238892 154356 238944
rect 223764 238892 223816 238944
rect 223856 238892 223908 238944
rect 227720 238892 227772 238944
rect 227996 238892 228048 238944
rect 231124 238892 231176 238944
rect 231584 238892 231636 238944
rect 235540 238892 235592 238944
rect 215944 238824 215996 238876
rect 238484 238824 238536 238876
rect 151544 238756 151596 238808
rect 221280 238756 221332 238808
rect 221464 238756 221516 238808
rect 223856 238756 223908 238808
rect 218980 238688 219032 238740
rect 219440 238688 219492 238740
rect 191656 238620 191708 238672
rect 222384 238620 222436 238672
rect 223120 238620 223172 238672
rect 232320 238756 232372 238808
rect 232412 238756 232464 238808
rect 239036 238756 239088 238808
rect 226432 238688 226484 238740
rect 235540 238688 235592 238740
rect 236000 238688 236052 238740
rect 225972 238620 226024 238672
rect 233516 238620 233568 238672
rect 233792 238620 233844 238672
rect 234436 238620 234488 238672
rect 234620 238620 234672 238672
rect 236368 238620 236420 238672
rect 237840 238688 237892 238740
rect 238024 238688 238076 238740
rect 242900 239028 242952 239080
rect 297640 239028 297692 239080
rect 242532 238960 242584 239012
rect 297548 238960 297600 239012
rect 241152 238892 241204 238944
rect 289360 238892 289412 238944
rect 247776 238824 247828 238876
rect 250168 238824 250220 238876
rect 255136 238824 255188 238876
rect 255688 238824 255740 238876
rect 255964 238824 256016 238876
rect 257528 238824 257580 238876
rect 258080 238824 258132 238876
rect 261116 238824 261168 238876
rect 261392 238824 261444 238876
rect 246856 238756 246908 238808
rect 248972 238756 249024 238808
rect 249156 238756 249208 238808
rect 241428 238688 241480 238740
rect 207664 238552 207716 238604
rect 232136 238552 232188 238604
rect 232320 238552 232372 238604
rect 235264 238552 235316 238604
rect 235540 238552 235592 238604
rect 238852 238552 238904 238604
rect 242900 238620 242952 238672
rect 260564 238756 260616 238808
rect 273260 238824 273312 238876
rect 251732 238688 251784 238740
rect 256516 238688 256568 238740
rect 258172 238688 258224 238740
rect 258816 238688 258868 238740
rect 252928 238620 252980 238672
rect 261576 238756 261628 238808
rect 266360 238756 266412 238808
rect 266544 238756 266596 238808
rect 267832 238756 267884 238808
rect 295248 238756 295300 238808
rect 488540 238756 488592 238808
rect 261300 238688 261352 238740
rect 262680 238688 262732 238740
rect 263692 238688 263744 238740
rect 266636 238688 266688 238740
rect 267280 238688 267332 238740
rect 271512 238688 271564 238740
rect 246672 238552 246724 238604
rect 255228 238552 255280 238604
rect 257160 238552 257212 238604
rect 257988 238552 258040 238604
rect 259736 238552 259788 238604
rect 270684 238620 270736 238672
rect 263968 238552 264020 238604
rect 264980 238552 265032 238604
rect 265072 238552 265124 238604
rect 278136 238552 278188 238604
rect 209044 238484 209096 238536
rect 221372 238484 221424 238536
rect 224868 238484 224920 238536
rect 226984 238484 227036 238536
rect 209136 238416 209188 238468
rect 229284 238416 229336 238468
rect 193772 238348 193824 238400
rect 224316 238348 224368 238400
rect 240784 238484 240836 238536
rect 241520 238484 241572 238536
rect 245660 238484 245712 238536
rect 246856 238484 246908 238536
rect 250168 238484 250220 238536
rect 250996 238484 251048 238536
rect 251180 238484 251232 238536
rect 255136 238484 255188 238536
rect 256700 238484 256752 238536
rect 259552 238484 259604 238536
rect 269120 238484 269172 238536
rect 296260 238484 296312 238536
rect 230848 238416 230900 238468
rect 161112 238280 161164 238332
rect 210608 238280 210660 238332
rect 219716 238280 219768 238332
rect 220544 238280 220596 238332
rect 222752 238280 222804 238332
rect 232596 238348 232648 238400
rect 236644 238348 236696 238400
rect 239036 238348 239088 238400
rect 241520 238348 241572 238400
rect 227904 238280 227956 238332
rect 228088 238280 228140 238332
rect 228916 238280 228968 238332
rect 240508 238280 240560 238332
rect 243728 238280 243780 238332
rect 268568 238416 268620 238468
rect 273536 238416 273588 238468
rect 295248 238416 295300 238468
rect 192484 238212 192536 238264
rect 219900 238212 219952 238264
rect 222936 238212 222988 238264
rect 230388 238212 230440 238264
rect 210240 238144 210292 238196
rect 231768 238212 231820 238264
rect 234896 238212 234948 238264
rect 237656 238212 237708 238264
rect 261576 238348 261628 238400
rect 248880 238280 248932 238332
rect 259736 238280 259788 238332
rect 262220 238280 262272 238332
rect 263600 238280 263652 238332
rect 255228 238212 255280 238264
rect 263048 238212 263100 238264
rect 231584 238144 231636 238196
rect 243728 238144 243780 238196
rect 259368 238144 259420 238196
rect 302976 238348 303028 238400
rect 265072 238280 265124 238332
rect 265440 238280 265492 238332
rect 266452 238280 266504 238332
rect 266820 238280 266872 238332
rect 267464 238280 267516 238332
rect 268200 238280 268252 238332
rect 268476 238280 268528 238332
rect 310244 238280 310296 238332
rect 269120 238212 269172 238264
rect 316960 238212 317012 238264
rect 264428 238144 264480 238196
rect 265808 238144 265860 238196
rect 267004 238144 267056 238196
rect 315396 238144 315448 238196
rect 161204 238076 161256 238128
rect 212356 238076 212408 238128
rect 220544 238076 220596 238128
rect 230664 238076 230716 238128
rect 231308 238076 231360 238128
rect 231492 238076 231544 238128
rect 239312 238076 239364 238128
rect 239496 238076 239548 238128
rect 248144 238076 248196 238128
rect 249340 238076 249392 238128
rect 260288 238076 260340 238128
rect 260380 238076 260432 238128
rect 266820 238076 266872 238128
rect 161296 238008 161348 238060
rect 237748 238008 237800 238060
rect 242532 238008 242584 238060
rect 245476 238008 245528 238060
rect 251732 238008 251784 238060
rect 255412 238008 255464 238060
rect 268200 238008 268252 238060
rect 217968 237940 218020 237992
rect 218888 237940 218940 237992
rect 223212 237940 223264 237992
rect 225604 237940 225656 237992
rect 234436 237940 234488 237992
rect 235448 237940 235500 237992
rect 236092 237940 236144 237992
rect 236644 237940 236696 237992
rect 210608 237872 210660 237924
rect 234620 237872 234672 237924
rect 237012 237872 237064 237924
rect 237656 237872 237708 237924
rect 238024 237872 238076 237924
rect 240232 237872 240284 237924
rect 240508 237872 240560 237924
rect 249064 237872 249116 237924
rect 251456 237940 251508 237992
rect 252836 237940 252888 237992
rect 254676 237940 254728 237992
rect 261300 237940 261352 237992
rect 266728 237940 266780 237992
rect 269764 238076 269816 238128
rect 269856 238076 269908 238128
rect 318340 238076 318392 238128
rect 268660 238008 268712 238060
rect 338396 238008 338448 238060
rect 268384 237940 268436 237992
rect 273536 237940 273588 237992
rect 258448 237872 258500 237924
rect 263416 237872 263468 237924
rect 274272 237872 274324 237924
rect 212356 237804 212408 237856
rect 236276 237804 236328 237856
rect 239220 237804 239272 237856
rect 208860 237736 208912 237788
rect 226616 237736 226668 237788
rect 226708 237736 226760 237788
rect 227076 237736 227128 237788
rect 227444 237736 227496 237788
rect 236920 237736 236972 237788
rect 240232 237736 240284 237788
rect 251456 237804 251508 237856
rect 251640 237804 251692 237856
rect 261576 237804 261628 237856
rect 268936 237804 268988 237856
rect 269028 237736 269080 237788
rect 161940 237464 161992 237516
rect 225420 237464 225472 237516
rect 161388 237396 161440 237448
rect 238392 237668 238444 237720
rect 232136 237600 232188 237652
rect 240140 237668 240192 237720
rect 241704 237668 241756 237720
rect 243728 237668 243780 237720
rect 270408 237668 270460 237720
rect 261576 237600 261628 237652
rect 263692 237600 263744 237652
rect 264704 237600 264756 237652
rect 265072 237600 265124 237652
rect 265348 237600 265400 237652
rect 265532 237600 265584 237652
rect 266176 237600 266228 237652
rect 226616 237532 226668 237584
rect 226892 237532 226944 237584
rect 231676 237532 231728 237584
rect 239220 237532 239272 237584
rect 225420 237328 225472 237380
rect 236000 237464 236052 237516
rect 239312 237464 239364 237516
rect 257804 237532 257856 237584
rect 263508 237532 263560 237584
rect 264244 237532 264296 237584
rect 272708 237532 272760 237584
rect 266728 237464 266780 237516
rect 266820 237464 266872 237516
rect 229376 237396 229428 237448
rect 230112 237396 230164 237448
rect 239036 237396 239088 237448
rect 244188 237396 244240 237448
rect 253572 237396 253624 237448
rect 254676 237396 254728 237448
rect 229284 237328 229336 237380
rect 230204 237328 230256 237380
rect 230756 237328 230808 237380
rect 231768 237328 231820 237380
rect 215852 237260 215904 237312
rect 220268 237260 220320 237312
rect 239128 237328 239180 237380
rect 258632 237328 258684 237380
rect 259276 237328 259328 237380
rect 261024 237328 261076 237380
rect 264980 237396 265032 237448
rect 267280 237328 267332 237380
rect 288532 237396 288584 237448
rect 288992 237396 289044 237448
rect 299020 237396 299072 237448
rect 301688 237396 301740 237448
rect 268844 237328 268896 237380
rect 235356 237260 235408 237312
rect 235724 237260 235776 237312
rect 243728 237260 243780 237312
rect 244004 237260 244056 237312
rect 251180 237260 251232 237312
rect 251456 237260 251508 237312
rect 253572 237260 253624 237312
rect 268476 237260 268528 237312
rect 275928 237328 275980 237380
rect 276296 237328 276348 237380
rect 330116 237260 330168 237312
rect 208400 237192 208452 237244
rect 209228 237192 209280 237244
rect 226248 237192 226300 237244
rect 226524 237192 226576 237244
rect 226800 237192 226852 237244
rect 234160 237192 234212 237244
rect 234344 237192 234396 237244
rect 240600 237192 240652 237244
rect 248420 237192 248472 237244
rect 256516 237192 256568 237244
rect 286876 237192 286928 237244
rect 214472 237124 214524 237176
rect 207848 237056 207900 237108
rect 222568 237056 222620 237108
rect 226984 237124 227036 237176
rect 229100 237124 229152 237176
rect 243820 237124 243872 237176
rect 275928 237124 275980 237176
rect 234712 237056 234764 237108
rect 244372 237056 244424 237108
rect 245108 237056 245160 237108
rect 247868 237056 247920 237108
rect 248236 237056 248288 237108
rect 208032 236988 208084 237040
rect 222476 236988 222528 237040
rect 222844 236988 222896 237040
rect 230020 236988 230072 237040
rect 236184 236988 236236 237040
rect 237472 236988 237524 237040
rect 244740 236988 244792 237040
rect 244924 236988 244976 237040
rect 211804 236920 211856 236972
rect 249248 236920 249300 236972
rect 253572 237056 253624 237108
rect 254400 237056 254452 237108
rect 261024 237056 261076 237108
rect 262864 237056 262916 237108
rect 289728 237056 289780 237108
rect 251548 236988 251600 237040
rect 274824 236988 274876 237040
rect 275376 236988 275428 237040
rect 251732 236920 251784 236972
rect 261024 236920 261076 236972
rect 262312 236920 262364 236972
rect 284392 236920 284444 236972
rect 284760 236920 284812 236972
rect 213092 236852 213144 236904
rect 254400 236852 254452 236904
rect 257344 236852 257396 236904
rect 259276 236852 259328 236904
rect 262588 236852 262640 236904
rect 274640 236852 274692 236904
rect 275652 236852 275704 236904
rect 197268 236784 197320 236836
rect 255688 236784 255740 236836
rect 257712 236784 257764 236836
rect 258264 236784 258316 236836
rect 261760 236784 261812 236836
rect 266912 236784 266964 236836
rect 159916 236716 159968 236768
rect 218888 236716 218940 236768
rect 218980 236716 219032 236768
rect 238576 236716 238628 236768
rect 241704 236716 241756 236768
rect 242256 236716 242308 236768
rect 244924 236716 244976 236768
rect 245200 236716 245252 236768
rect 268660 236716 268712 236768
rect 269580 236716 269632 236768
rect 295340 236716 295392 236768
rect 155592 236648 155644 236700
rect 213828 236648 213880 236700
rect 220176 236648 220228 236700
rect 257344 236648 257396 236700
rect 258264 236648 258316 236700
rect 258908 236648 258960 236700
rect 265440 236648 265492 236700
rect 287980 236648 288032 236700
rect 334992 236648 335044 236700
rect 209504 236580 209556 236632
rect 227812 236580 227864 236632
rect 227996 236580 228048 236632
rect 229100 236580 229152 236632
rect 231216 236580 231268 236632
rect 237472 236580 237524 236632
rect 237748 236580 237800 236632
rect 242072 236580 242124 236632
rect 242256 236580 242308 236632
rect 244004 236580 244056 236632
rect 244648 236580 244700 236632
rect 247960 236580 248012 236632
rect 248328 236580 248380 236632
rect 248972 236580 249024 236632
rect 249708 236580 249760 236632
rect 252836 236580 252888 236632
rect 265532 236580 265584 236632
rect 213828 236512 213880 236564
rect 223948 236444 224000 236496
rect 224316 236444 224368 236496
rect 224684 236512 224736 236564
rect 224868 236512 224920 236564
rect 230756 236512 230808 236564
rect 230940 236512 230992 236564
rect 241888 236512 241940 236564
rect 242440 236512 242492 236564
rect 253480 236512 253532 236564
rect 262772 236512 262824 236564
rect 226064 236444 226116 236496
rect 258448 236444 258500 236496
rect 269856 236512 269908 236564
rect 223764 236376 223816 236428
rect 226340 236376 226392 236428
rect 238208 236376 238260 236428
rect 247868 236376 247920 236428
rect 327724 236376 327776 236428
rect 265900 236308 265952 236360
rect 266820 236308 266872 236360
rect 245108 236240 245160 236292
rect 245568 236240 245620 236292
rect 261024 236240 261076 236292
rect 261852 236240 261904 236292
rect 214472 236172 214524 236224
rect 215024 236172 215076 236224
rect 226432 236104 226484 236156
rect 227628 236104 227680 236156
rect 261484 236104 261536 236156
rect 276204 236104 276256 236156
rect 261208 236036 261260 236088
rect 267280 236036 267332 236088
rect 207756 235968 207808 236020
rect 208032 235968 208084 236020
rect 217692 235968 217744 236020
rect 244648 235968 244700 236020
rect 255320 235968 255372 236020
rect 255688 235968 255740 236020
rect 285588 235968 285640 236020
rect 286876 235968 286928 236020
rect 289360 235968 289412 236020
rect 289728 235968 289780 236020
rect 210884 235900 210936 235952
rect 217324 235900 217376 235952
rect 219164 235900 219216 235952
rect 221832 235900 221884 235952
rect 222016 235900 222068 235952
rect 233424 235900 233476 235952
rect 233700 235900 233752 235952
rect 233884 235900 233936 235952
rect 237472 235900 237524 235952
rect 253112 235900 253164 235952
rect 253664 235900 253716 235952
rect 274548 235900 274600 235952
rect 330024 235900 330076 235952
rect 223764 235832 223816 235884
rect 259828 235832 259880 235884
rect 268292 235832 268344 235884
rect 285680 235832 285732 235884
rect 286968 235832 287020 235884
rect 287704 235832 287756 235884
rect 240232 235764 240284 235816
rect 276020 235764 276072 235816
rect 223856 235696 223908 235748
rect 224500 235696 224552 235748
rect 226156 235696 226208 235748
rect 226524 235696 226576 235748
rect 244924 235696 244976 235748
rect 291108 235696 291160 235748
rect 236000 235628 236052 235680
rect 279976 235628 280028 235680
rect 221004 235560 221056 235612
rect 233056 235560 233108 235612
rect 244740 235560 244792 235612
rect 285680 235560 285732 235612
rect 222016 235492 222068 235544
rect 230480 235492 230532 235544
rect 232872 235492 232924 235544
rect 234620 235492 234672 235544
rect 242808 235492 242860 235544
rect 283564 235492 283616 235544
rect 216036 235424 216088 235476
rect 236552 235424 236604 235476
rect 243820 235424 243872 235476
rect 248604 235424 248656 235476
rect 269488 235424 269540 235476
rect 269580 235424 269632 235476
rect 270132 235424 270184 235476
rect 282736 235424 282788 235476
rect 211068 235356 211120 235408
rect 221004 235356 221056 235408
rect 239220 235356 239272 235408
rect 239772 235356 239824 235408
rect 243176 235356 243228 235408
rect 262864 235356 262916 235408
rect 268292 235356 268344 235408
rect 270408 235356 270460 235408
rect 280896 235356 280948 235408
rect 218888 235288 218940 235340
rect 244740 235288 244792 235340
rect 253480 235288 253532 235340
rect 253848 235288 253900 235340
rect 262036 235288 262088 235340
rect 277400 235288 277452 235340
rect 219256 235220 219308 235272
rect 255596 235220 255648 235272
rect 263140 235220 263192 235272
rect 282552 235220 282604 235272
rect 331404 235220 331456 235272
rect 239312 235152 239364 235204
rect 240048 235152 240100 235204
rect 243084 235152 243136 235204
rect 243544 235152 243596 235204
rect 252008 235152 252060 235204
rect 265072 235152 265124 235204
rect 267280 235152 267332 235204
rect 269764 235152 269816 235204
rect 278596 235152 278648 235204
rect 227076 235084 227128 235136
rect 239404 235084 239456 235136
rect 254768 235084 254820 235136
rect 269028 235084 269080 235136
rect 216312 235016 216364 235068
rect 227444 235016 227496 235068
rect 240784 235016 240836 235068
rect 300492 235016 300544 235068
rect 216220 234948 216272 235000
rect 210608 234880 210660 234932
rect 217232 234880 217284 234932
rect 235264 234948 235316 235000
rect 294972 234948 295024 235000
rect 254032 234880 254084 234932
rect 255228 234880 255280 234932
rect 245568 234812 245620 234864
rect 245844 234812 245896 234864
rect 213552 234744 213604 234796
rect 246488 234744 246540 234796
rect 246856 234744 246908 234796
rect 210792 234676 210844 234728
rect 217232 234676 217284 234728
rect 247316 234676 247368 234728
rect 247776 234676 247828 234728
rect 256792 234676 256844 234728
rect 257896 234676 257948 234728
rect 258448 234608 258500 234660
rect 291108 234608 291160 234660
rect 291844 234608 291896 234660
rect 214748 234540 214800 234592
rect 215208 234540 215260 234592
rect 240600 234540 240652 234592
rect 244648 234540 244700 234592
rect 249156 234540 249208 234592
rect 257896 234540 257948 234592
rect 260104 234540 260156 234592
rect 267648 234540 267700 234592
rect 272708 234540 272760 234592
rect 273168 234540 273220 234592
rect 286508 234540 286560 234592
rect 243452 234472 243504 234524
rect 303068 234472 303120 234524
rect 208492 234404 208544 234456
rect 209320 234404 209372 234456
rect 239036 234404 239088 234456
rect 245752 234404 245804 234456
rect 300400 234404 300452 234456
rect 202328 234336 202380 234388
rect 202604 234336 202656 234388
rect 228180 234336 228232 234388
rect 237564 234336 237616 234388
rect 282828 234336 282880 234388
rect 188896 234064 188948 234116
rect 214748 234064 214800 234116
rect 184848 233996 184900 234048
rect 211620 233996 211672 234048
rect 244280 234268 244332 234320
rect 250536 234268 250588 234320
rect 258724 234268 258776 234320
rect 259276 234268 259328 234320
rect 306012 234268 306064 234320
rect 235264 234200 235316 234252
rect 235632 234200 235684 234252
rect 276480 234200 276532 234252
rect 235356 234132 235408 234184
rect 275560 234132 275612 234184
rect 239128 234064 239180 234116
rect 239680 234064 239732 234116
rect 279332 234064 279384 234116
rect 241244 233996 241296 234048
rect 242348 233996 242400 234048
rect 280804 233996 280856 234048
rect 172336 233928 172388 233980
rect 202604 233928 202656 233980
rect 235172 233928 235224 233980
rect 235816 233928 235868 233980
rect 156972 233860 157024 233912
rect 208400 233860 208452 233912
rect 211896 233860 211948 233912
rect 212448 233860 212500 233912
rect 216404 233860 216456 233912
rect 250904 233928 250956 233980
rect 258724 233928 258776 233980
rect 284208 233928 284260 233980
rect 241704 233860 241756 233912
rect 242716 233860 242768 233912
rect 243728 233860 243780 233912
rect 278780 233860 278832 233912
rect 280068 233860 280120 233912
rect 246396 233792 246448 233844
rect 257896 233792 257948 233844
rect 284024 233792 284076 233844
rect 232872 233724 232924 233776
rect 233148 233724 233200 233776
rect 239956 233724 240008 233776
rect 218704 233656 218756 233708
rect 251088 233656 251140 233708
rect 272892 233724 272944 233776
rect 263784 233656 263836 233708
rect 264704 233656 264756 233708
rect 267648 233656 267700 233708
rect 270132 233656 270184 233708
rect 278504 233656 278556 233708
rect 253572 233452 253624 233504
rect 253848 233452 253900 233504
rect 242992 233384 243044 233436
rect 243636 233384 243688 233436
rect 239588 233316 239640 233368
rect 298928 233588 298980 233640
rect 226524 233248 226576 233300
rect 227352 233248 227404 233300
rect 245384 233248 245436 233300
rect 245752 233248 245804 233300
rect 205640 233180 205692 233232
rect 206560 233180 206612 233232
rect 229008 233180 229060 233232
rect 246120 233180 246172 233232
rect 246672 233180 246724 233232
rect 253480 233180 253532 233232
rect 253848 233180 253900 233232
rect 254032 233180 254084 233232
rect 269672 233180 269724 233232
rect 270316 233180 270368 233232
rect 270592 233180 270644 233232
rect 276388 233180 276440 233232
rect 579620 233180 579672 233232
rect 251088 233112 251140 233164
rect 309968 233112 310020 233164
rect 236736 233044 236788 233096
rect 237012 233044 237064 233096
rect 295984 233044 296036 233096
rect 246212 232976 246264 233028
rect 305736 232976 305788 233028
rect 249800 232908 249852 232960
rect 253204 232908 253256 232960
rect 253848 232908 253900 232960
rect 296352 232908 296404 232960
rect 236736 232840 236788 232892
rect 277676 232840 277728 232892
rect 250168 232772 250220 232824
rect 251088 232772 251140 232824
rect 253204 232772 253256 232824
rect 286416 232772 286468 232824
rect 191748 232704 191800 232756
rect 216404 232704 216456 232756
rect 240784 232704 240836 232756
rect 194416 232636 194468 232688
rect 221924 232636 221976 232688
rect 244188 232636 244240 232688
rect 273720 232636 273772 232688
rect 276020 232704 276072 232756
rect 277032 232704 277084 232756
rect 279608 232704 279660 232756
rect 281540 232704 281592 232756
rect 293408 232704 293460 232756
rect 276848 232636 276900 232688
rect 283564 232636 283616 232688
rect 329932 232636 329984 232688
rect 152832 232568 152884 232620
rect 205640 232568 205692 232620
rect 228548 232568 228600 232620
rect 231860 232568 231912 232620
rect 237288 232568 237340 232620
rect 238944 232568 238996 232620
rect 252284 232568 252336 232620
rect 279700 232568 279752 232620
rect 334072 232568 334124 232620
rect 161480 232500 161532 232552
rect 191656 232500 191708 232552
rect 193128 232500 193180 232552
rect 252468 232500 252520 232552
rect 254032 232500 254084 232552
rect 262772 232500 262824 232552
rect 276020 232500 276072 232552
rect 280252 232500 280304 232552
rect 337016 232500 337068 232552
rect 248052 232432 248104 232484
rect 270040 232432 270092 232484
rect 270684 232432 270736 232484
rect 270960 232432 271012 232484
rect 265072 232296 265124 232348
rect 283564 232364 283616 232416
rect 236920 232228 236972 232280
rect 237104 232228 237156 232280
rect 279516 232228 279568 232280
rect 270592 232160 270644 232212
rect 271604 232160 271656 232212
rect 273628 232160 273680 232212
rect 274272 232160 274324 232212
rect 270040 232092 270092 232144
rect 275284 232092 275336 232144
rect 233700 232024 233752 232076
rect 234252 232024 234304 232076
rect 241060 231956 241112 232008
rect 241336 231956 241388 232008
rect 256884 231956 256936 232008
rect 261576 231956 261628 232008
rect 195888 231820 195940 231872
rect 252560 231820 252612 231872
rect 255596 231820 255648 231872
rect 256608 231820 256660 231872
rect 256884 231820 256936 231872
rect 258080 231820 258132 231872
rect 199016 231752 199068 231804
rect 200028 231752 200080 231804
rect 228732 231752 228784 231804
rect 233424 231752 233476 231804
rect 234068 231752 234120 231804
rect 262864 231752 262916 231804
rect 274916 231752 274968 231804
rect 275744 231752 275796 231804
rect 276112 231752 276164 231804
rect 276940 231752 276992 231804
rect 293224 231684 293276 231736
rect 250996 231616 251048 231668
rect 301780 231616 301832 231668
rect 199844 231548 199896 231600
rect 259368 231548 259420 231600
rect 247408 231480 247460 231532
rect 296076 231480 296128 231532
rect 232044 231412 232096 231464
rect 232412 231412 232464 231464
rect 244096 231412 244148 231464
rect 275468 231412 275520 231464
rect 248972 231344 249024 231396
rect 280252 231344 280304 231396
rect 253572 231276 253624 231328
rect 283748 231276 283800 231328
rect 152740 231208 152792 231260
rect 199016 231208 199068 231260
rect 248144 231208 248196 231260
rect 276112 231208 276164 231260
rect 289728 231208 289780 231260
rect 332784 231208 332836 231260
rect 256424 231140 256476 231192
rect 290648 231140 290700 231192
rect 336924 231140 336976 231192
rect 196992 231072 197044 231124
rect 256976 231072 257028 231124
rect 261576 231072 261628 231124
rect 338304 231072 338356 231124
rect 260288 231004 260340 231056
rect 281540 231004 281592 231056
rect 269028 230936 269080 230988
rect 289176 230936 289228 230988
rect 289728 230936 289780 230988
rect 239404 230868 239456 230920
rect 298652 230868 298704 230920
rect 252928 230800 252980 230852
rect 312912 230800 312964 230852
rect 247408 230732 247460 230784
rect 248144 230732 248196 230784
rect 255504 230732 255556 230784
rect 256516 230732 256568 230784
rect 199936 230664 199988 230716
rect 259460 230664 259512 230716
rect 197176 230596 197228 230648
rect 255136 230596 255188 230648
rect 199752 230528 199804 230580
rect 259276 230596 259328 230648
rect 198648 230460 198700 230512
rect 257712 230460 257764 230512
rect 214748 230392 214800 230444
rect 216128 230392 216180 230444
rect 232780 230392 232832 230444
rect 233516 230392 233568 230444
rect 244280 230392 244332 230444
rect 245108 230392 245160 230444
rect 249800 230392 249852 230444
rect 250444 230392 250496 230444
rect 271420 230460 271472 230512
rect 271144 230392 271196 230444
rect 273444 230392 273496 230444
rect 274456 230392 274508 230444
rect 275468 230392 275520 230444
rect 244188 230256 244240 230308
rect 244280 230256 244332 230308
rect 239404 230188 239456 230240
rect 240048 230188 240100 230240
rect 301596 230324 301648 230376
rect 245200 230256 245252 230308
rect 303620 230256 303672 230308
rect 304448 230188 304500 230240
rect 221832 230120 221884 230172
rect 243728 230120 243780 230172
rect 246948 230120 247000 230172
rect 249340 230120 249392 230172
rect 298836 230120 298888 230172
rect 233976 230052 234028 230104
rect 240416 230052 240468 230104
rect 288348 230052 288400 230104
rect 215208 229984 215260 230036
rect 240508 229984 240560 230036
rect 280988 229984 281040 230036
rect 212448 229916 212500 229968
rect 239956 229916 240008 229968
rect 242624 229916 242676 229968
rect 282276 229916 282328 229968
rect 212264 229848 212316 229900
rect 239128 229848 239180 229900
rect 244832 229848 244884 229900
rect 245200 229848 245252 229900
rect 246212 229848 246264 229900
rect 246580 229848 246632 229900
rect 269304 229848 269356 229900
rect 269396 229848 269448 229900
rect 276756 229848 276808 229900
rect 223580 229780 223632 229832
rect 224868 229780 224920 229832
rect 233516 229780 233568 229832
rect 278320 229780 278372 229832
rect 218704 229712 218756 229764
rect 234896 229712 234948 229764
rect 223764 229644 223816 229696
rect 224040 229644 224092 229696
rect 228732 229644 228784 229696
rect 244648 229712 244700 229764
rect 245476 229712 245528 229764
rect 246028 229712 246080 229764
rect 246580 229712 246632 229764
rect 248420 229712 248472 229764
rect 249524 229712 249576 229764
rect 251272 229712 251324 229764
rect 252376 229712 252428 229764
rect 252560 229712 252612 229764
rect 253756 229712 253808 229764
rect 254032 229712 254084 229764
rect 254952 229712 255004 229764
rect 255504 229712 255556 229764
rect 256332 229712 256384 229764
rect 265532 229712 265584 229764
rect 285036 229712 285088 229764
rect 335452 229712 335504 229764
rect 249800 229644 249852 229696
rect 254308 229644 254360 229696
rect 254584 229644 254636 229696
rect 269304 229644 269356 229696
rect 272984 229644 273036 229696
rect 227168 229576 227220 229628
rect 241520 229576 241572 229628
rect 241612 229576 241664 229628
rect 242164 229576 242216 229628
rect 245476 229576 245528 229628
rect 249340 229576 249392 229628
rect 253572 229576 253624 229628
rect 253756 229576 253808 229628
rect 259828 229576 259880 229628
rect 260840 229576 260892 229628
rect 223764 229508 223816 229560
rect 224224 229508 224276 229560
rect 239588 229508 239640 229560
rect 256148 229508 256200 229560
rect 222108 229440 222160 229492
rect 302884 229440 302936 229492
rect 201224 229372 201276 229424
rect 271972 229372 272024 229424
rect 241520 229304 241572 229356
rect 248328 229304 248380 229356
rect 223304 229100 223356 229152
rect 244188 229100 244240 229152
rect 208216 229032 208268 229084
rect 226616 229032 226668 229084
rect 237288 229032 237340 229084
rect 298744 229032 298796 229084
rect 161572 228964 161624 229016
rect 207848 228964 207900 229016
rect 156696 228896 156748 228948
rect 208124 228896 208176 228948
rect 226064 228964 226116 229016
rect 263784 228964 263836 229016
rect 325148 228964 325200 229016
rect 210884 228896 210936 228948
rect 237472 228896 237524 228948
rect 262312 228896 262364 228948
rect 323676 228896 323728 228948
rect 156788 228828 156840 228880
rect 208216 228828 208268 228880
rect 211068 228828 211120 228880
rect 237288 228828 237340 228880
rect 264428 228828 264480 228880
rect 264796 228828 264848 228880
rect 325056 228828 325108 228880
rect 156880 228760 156932 228812
rect 210976 228760 211028 228812
rect 235540 228760 235592 228812
rect 294420 228760 294472 228812
rect 159640 228692 159692 228744
rect 214932 228692 214984 228744
rect 217784 228692 217836 228744
rect 240784 228692 240836 228744
rect 264520 228692 264572 228744
rect 323768 228692 323820 228744
rect 202328 228624 202380 228676
rect 270500 228624 270552 228676
rect 200212 228556 200264 228608
rect 270776 228556 270828 228608
rect 197912 228488 197964 228540
rect 272156 228488 272208 228540
rect 159732 228420 159784 228472
rect 234804 228420 234856 228472
rect 236552 228420 236604 228472
rect 237656 228420 237708 228472
rect 297456 228420 297508 228472
rect 162032 228352 162084 228404
rect 239680 228352 239732 228404
rect 260012 228352 260064 228404
rect 319444 228352 319496 228404
rect 235172 228284 235224 228336
rect 291936 228284 291988 228336
rect 236460 228216 236512 228268
rect 288164 228216 288216 228268
rect 245016 228148 245068 228200
rect 269304 228148 269356 228200
rect 227720 227808 227772 227860
rect 228640 227808 228692 227860
rect 263784 227808 263836 227860
rect 264244 227808 264296 227860
rect 235172 227740 235224 227792
rect 235632 227740 235684 227792
rect 261760 227672 261812 227724
rect 271328 227672 271380 227724
rect 238116 227604 238168 227656
rect 260012 227604 260064 227656
rect 231124 227536 231176 227588
rect 244464 227536 244516 227588
rect 252100 227536 252152 227588
rect 313004 227536 313056 227588
rect 239680 227468 239732 227520
rect 259920 227468 259972 227520
rect 260564 227468 260616 227520
rect 321100 227468 321152 227520
rect 234160 227400 234212 227452
rect 282644 227400 282696 227452
rect 228456 227332 228508 227384
rect 248972 227332 249024 227384
rect 256700 227332 256752 227384
rect 304356 227332 304408 227384
rect 238576 227264 238628 227316
rect 262956 227264 263008 227316
rect 223212 227196 223264 227248
rect 249340 227196 249392 227248
rect 258264 227196 258316 227248
rect 292580 227196 292632 227248
rect 161664 227128 161716 227180
rect 207756 227128 207808 227180
rect 223120 227128 223172 227180
rect 237380 227128 237432 227180
rect 238484 227128 238536 227180
rect 265164 227128 265216 227180
rect 291752 227128 291804 227180
rect 292212 227128 292264 227180
rect 328552 227128 328604 227180
rect 161020 227060 161072 227112
rect 236920 227060 236972 227112
rect 263508 227060 263560 227112
rect 291936 227060 291988 227112
rect 335360 227060 335412 227112
rect 160928 226992 160980 227044
rect 236552 226992 236604 227044
rect 257620 226992 257672 227044
rect 291752 226992 291804 227044
rect 292580 226992 292632 227044
rect 293224 226992 293276 227044
rect 338120 226992 338172 227044
rect 224408 226924 224460 226976
rect 224592 226924 224644 226976
rect 239772 226924 239824 226976
rect 259644 226924 259696 226976
rect 237012 226856 237064 226908
rect 259736 226856 259788 226908
rect 240876 226788 240928 226840
rect 260932 226856 260984 226908
rect 338212 226788 338264 226840
rect 248696 226720 248748 226772
rect 249616 226720 249668 226772
rect 262404 226720 262456 226772
rect 339592 226720 339644 226772
rect 270776 226312 270828 226364
rect 271328 226312 271380 226364
rect 241888 226244 241940 226296
rect 327356 226244 327408 226296
rect 239036 226176 239088 226228
rect 239220 226176 239272 226228
rect 300216 226176 300268 226228
rect 246488 226108 246540 226160
rect 246764 226108 246816 226160
rect 251824 226108 251876 226160
rect 311348 226108 311400 226160
rect 246856 226040 246908 226092
rect 305644 226040 305696 226092
rect 247776 225972 247828 226024
rect 307024 225972 307076 226024
rect 243084 225904 243136 225956
rect 301504 225904 301556 225956
rect 246120 225836 246172 225888
rect 246856 225836 246908 225888
rect 259276 225836 259328 225888
rect 314108 225836 314160 225888
rect 222016 225768 222068 225820
rect 239036 225768 239088 225820
rect 245568 225768 245620 225820
rect 299572 225768 299624 225820
rect 300584 225768 300636 225820
rect 163504 225700 163556 225752
rect 232044 225700 232096 225752
rect 244188 225700 244240 225752
rect 296720 225700 296772 225752
rect 297732 225700 297784 225752
rect 154212 225632 154264 225684
rect 229928 225632 229980 225684
rect 246488 225632 246540 225684
rect 305920 225632 305972 225684
rect 160836 225564 160888 225616
rect 236460 225564 236512 225616
rect 260932 225564 260984 225616
rect 327448 225564 327500 225616
rect 241796 225496 241848 225548
rect 292396 225496 292448 225548
rect 241888 225428 241940 225480
rect 242532 225428 242584 225480
rect 243084 225428 243136 225480
rect 243544 225428 243596 225480
rect 242624 225360 242676 225412
rect 289268 225428 289320 225480
rect 267096 225360 267148 225412
rect 267372 225360 267424 225412
rect 241704 224952 241756 225004
rect 242624 224952 242676 225004
rect 260196 224884 260248 224936
rect 262404 224884 262456 224936
rect 263048 224884 263100 224936
rect 273444 224884 273496 224936
rect 273904 224884 273956 224936
rect 310060 224816 310112 224868
rect 248696 224748 248748 224800
rect 249432 224748 249484 224800
rect 252008 224748 252060 224800
rect 252376 224748 252428 224800
rect 311532 224748 311584 224800
rect 232504 224680 232556 224732
rect 292028 224680 292080 224732
rect 232688 224612 232740 224664
rect 238300 224612 238352 224664
rect 297364 224612 297416 224664
rect 238392 224544 238444 224596
rect 296168 224544 296220 224596
rect 240048 224476 240100 224528
rect 294696 224476 294748 224528
rect 240784 224408 240836 224460
rect 241428 224408 241480 224460
rect 288072 224408 288124 224460
rect 240968 224340 241020 224392
rect 282368 224340 282420 224392
rect 233700 224272 233752 224324
rect 273996 224272 274048 224324
rect 226248 224204 226300 224256
rect 239312 224204 239364 224256
rect 240048 224204 240100 224256
rect 241060 224204 241112 224256
rect 241520 224204 241572 224256
rect 283656 224204 283708 224256
rect 241612 224136 241664 224188
rect 251272 224136 251324 224188
rect 286324 224136 286376 224188
rect 243728 224068 243780 224120
rect 244004 224068 244056 224120
rect 277124 224068 277176 224120
rect 206928 224000 206980 224052
rect 229836 224000 229888 224052
rect 237932 224000 237984 224052
rect 300860 224000 300912 224052
rect 265532 223932 265584 223984
rect 265808 223932 265860 223984
rect 206836 223796 206888 223848
rect 227352 223592 227404 223644
rect 233700 223592 233752 223644
rect 258632 223592 258684 223644
rect 264152 223592 264204 223644
rect 258816 223524 258868 223576
rect 259184 223524 259236 223576
rect 319812 223524 319864 223576
rect 259368 223456 259420 223508
rect 262956 223456 263008 223508
rect 264152 223456 264204 223508
rect 319720 223456 319772 223508
rect 256884 223388 256936 223440
rect 257344 223388 257396 223440
rect 318248 223388 318300 223440
rect 256792 223320 256844 223372
rect 257436 223320 257488 223372
rect 318156 223320 318208 223372
rect 257712 223252 257764 223304
rect 254216 223184 254268 223236
rect 254860 223184 254912 223236
rect 262956 223252 263008 223304
rect 316684 223252 316736 223304
rect 255596 223116 255648 223168
rect 256148 223116 256200 223168
rect 259368 223116 259420 223168
rect 316868 223184 316920 223236
rect 314292 223116 314344 223168
rect 254308 223048 254360 223100
rect 314200 223048 314252 223100
rect 289084 222980 289136 223032
rect 158628 222912 158680 222964
rect 205640 222912 205692 222964
rect 229376 222912 229428 222964
rect 230020 222912 230072 222964
rect 232780 222912 232832 222964
rect 276664 222912 276716 222964
rect 162308 222844 162360 222896
rect 237104 222844 237156 222896
rect 247500 222844 247552 222896
rect 247776 222844 247828 222896
rect 306472 222980 306524 223032
rect 307116 222980 307168 223032
rect 253112 222776 253164 222828
rect 271972 222776 272024 222828
rect 272524 222776 272576 222828
rect 262312 222708 262364 222760
rect 262956 222708 263008 222760
rect 242992 222096 243044 222148
rect 243636 222096 243688 222148
rect 248604 222096 248656 222148
rect 249340 222096 249392 222148
rect 252744 222096 252796 222148
rect 253204 222096 253256 222148
rect 254124 222096 254176 222148
rect 254676 222096 254728 222148
rect 254952 222096 255004 222148
rect 328460 222096 328512 222148
rect 252652 222028 252704 222080
rect 253480 222028 253532 222080
rect 252192 221960 252244 222012
rect 312820 222028 312872 222080
rect 254768 221960 254820 222012
rect 315304 221960 315356 222012
rect 232596 221892 232648 221944
rect 253296 221892 253348 221944
rect 254952 221892 255004 221944
rect 255504 221892 255556 221944
rect 255964 221892 256016 221944
rect 316776 221892 316828 221944
rect 253940 221824 253992 221876
rect 254676 221824 254728 221876
rect 314384 221824 314436 221876
rect 253480 221756 253532 221808
rect 312636 221756 312688 221808
rect 253204 221688 253256 221740
rect 312728 221688 312780 221740
rect 243636 221620 243688 221672
rect 287888 221620 287940 221672
rect 230756 221552 230808 221604
rect 231492 221552 231544 221604
rect 271880 221552 271932 221604
rect 228640 221484 228692 221536
rect 262220 221484 262272 221536
rect 162216 221416 162268 221468
rect 236736 221416 236788 221468
rect 249340 221416 249392 221468
rect 339500 221416 339552 221468
rect 254032 221348 254084 221400
rect 254768 221348 254820 221400
rect 223948 220736 224000 220788
rect 224316 220736 224368 220788
rect 227444 220736 227496 220788
rect 288256 220736 288308 220788
rect 223856 220668 223908 220720
rect 224500 220668 224552 220720
rect 224316 220600 224368 220652
rect 284484 220668 284536 220720
rect 224500 220464 224552 220516
rect 284300 220600 284352 220652
rect 226432 220396 226484 220448
rect 227444 220396 227496 220448
rect 286600 220532 286652 220584
rect 226524 220260 226576 220312
rect 227260 220260 227312 220312
rect 229284 220260 229336 220312
rect 283840 220464 283892 220516
rect 225880 220192 225932 220244
rect 275008 220396 275060 220448
rect 248512 220328 248564 220380
rect 249156 220328 249208 220380
rect 158076 220056 158128 220108
rect 229284 220056 229336 220108
rect 249156 220056 249208 220108
rect 309784 220056 309836 220108
rect 229192 219376 229244 219428
rect 229928 219376 229980 219428
rect 228916 219308 228968 219360
rect 289452 219376 289504 219428
rect 230572 219308 230624 219360
rect 231768 219308 231820 219360
rect 290464 219308 290516 219360
rect 246396 219240 246448 219292
rect 249984 219240 250036 219292
rect 309876 219240 309928 219292
rect 256516 219172 256568 219224
rect 314016 219172 314068 219224
rect 246764 219104 246816 219156
rect 289544 219104 289596 219156
rect 229928 219036 229980 219088
rect 273352 219036 273404 219088
rect 243912 218968 243964 219020
rect 282184 218968 282236 219020
rect 152648 218764 152700 218816
rect 228272 218764 228324 218816
rect 228916 218764 228968 218816
rect 160744 218696 160796 218748
rect 237564 218696 237616 218748
rect 249524 218696 249576 218748
rect 335360 218696 335412 218748
rect 336004 218696 336056 218748
rect 249248 218016 249300 218068
rect 249524 218016 249576 218068
rect 204168 217948 204220 218000
rect 225512 217948 225564 218000
rect 180156 217404 180208 217456
rect 212908 217404 212960 217456
rect 303620 217404 303672 217456
rect 304264 217404 304316 217456
rect 165344 217336 165396 217388
rect 204168 217336 204220 217388
rect 166816 217268 166868 217320
rect 226708 217268 226760 217320
rect 246580 217268 246632 217320
rect 303620 217268 303672 217320
rect 205640 216588 205692 216640
rect 206928 216588 206980 216640
rect 224684 216588 224736 216640
rect 188620 216044 188672 216096
rect 213000 216044 213052 216096
rect 155408 215976 155460 216028
rect 205640 215976 205692 216028
rect 161756 215908 161808 215960
rect 223488 215908 223540 215960
rect 247132 215908 247184 215960
rect 247868 215908 247920 215960
rect 317420 215908 317472 215960
rect 205640 215228 205692 215280
rect 206836 215228 206888 215280
rect 227536 215228 227588 215280
rect 173900 214684 173952 214736
rect 174728 214684 174780 214736
rect 176108 214684 176160 214736
rect 210516 214684 210568 214736
rect 159364 214616 159416 214668
rect 205640 214616 205692 214668
rect 3424 214548 3476 214600
rect 200764 214548 200816 214600
rect 252560 214548 252612 214600
rect 253572 214548 253624 214600
rect 313924 214548 313976 214600
rect 167000 214480 167052 214532
rect 167736 214480 167788 214532
rect 168380 214480 168432 214532
rect 168840 214480 168892 214532
rect 169760 214480 169812 214532
rect 170312 214480 170364 214532
rect 171140 214480 171192 214532
rect 172152 214480 172204 214532
rect 172520 214480 172572 214532
rect 173256 214480 173308 214532
rect 173992 214480 174044 214532
rect 174360 214480 174412 214532
rect 186412 214480 186464 214532
rect 186872 214480 186924 214532
rect 187792 214480 187844 214532
rect 188988 214480 189040 214532
rect 189080 214480 189132 214532
rect 189816 214480 189868 214532
rect 190460 214480 190512 214532
rect 190920 214480 190972 214532
rect 191932 214480 191984 214532
rect 193036 214480 193088 214532
rect 193312 214480 193364 214532
rect 193496 214480 193548 214532
rect 194600 214480 194652 214532
rect 195336 214480 195388 214532
rect 186320 214412 186372 214464
rect 187240 214412 187292 214464
rect 189172 214412 189224 214464
rect 189448 214412 189500 214464
rect 190552 214412 190604 214464
rect 190736 214412 190788 214464
rect 193220 214412 193272 214464
rect 194508 214412 194560 214464
rect 194692 214412 194744 214464
rect 194968 214412 195020 214464
rect 186412 214344 186464 214396
rect 186688 214344 186740 214396
rect 201408 213868 201460 213920
rect 223580 213868 223632 213920
rect 182364 213392 182416 213444
rect 210700 213392 210752 213444
rect 181996 213324 182048 213376
rect 216496 213324 216548 213376
rect 157984 213256 158036 213308
rect 201408 213256 201460 213308
rect 242532 213256 242584 213308
rect 252560 213256 252612 213308
rect 184756 213188 184808 213240
rect 244372 213188 244424 213240
rect 250628 213188 250680 213240
rect 311164 213188 311216 213240
rect 175740 212440 175792 212492
rect 180064 212440 180116 212492
rect 199384 212440 199436 212492
rect 220360 212440 220412 212492
rect 173900 212372 173952 212424
rect 178684 212372 178736 212424
rect 181260 212372 181312 212424
rect 184204 212372 184256 212424
rect 184388 212372 184440 212424
rect 176660 212304 176712 212356
rect 176936 212304 176988 212356
rect 183560 212304 183612 212356
rect 184296 212304 184348 212356
rect 184940 212304 184992 212356
rect 185400 212304 185452 212356
rect 205548 212372 205600 212424
rect 197084 212304 197136 212356
rect 164240 212236 164292 212288
rect 164792 212236 164844 212288
rect 165712 212236 165764 212288
rect 166908 212236 166960 212288
rect 176844 212236 176896 212288
rect 177672 212236 177724 212288
rect 178040 212236 178092 212288
rect 178776 212236 178828 212288
rect 183652 212236 183704 212288
rect 183928 212236 183980 212288
rect 185124 212236 185176 212288
rect 185768 212236 185820 212288
rect 185860 212236 185912 212288
rect 188344 212236 188396 212288
rect 195980 212236 196032 212288
rect 196440 212236 196492 212288
rect 197360 212236 197412 212288
rect 198556 212236 198608 212288
rect 198924 212236 198976 212288
rect 200028 212236 200080 212288
rect 221648 212236 221700 212288
rect 173532 212168 173584 212220
rect 173808 212168 173860 212220
rect 188804 212168 188856 212220
rect 194140 212168 194192 212220
rect 221556 212168 221608 212220
rect 175372 212100 175424 212152
rect 216588 212100 216640 212152
rect 159272 212032 159324 212084
rect 201224 212032 201276 212084
rect 202696 212032 202748 212084
rect 203340 212032 203392 212084
rect 204076 212032 204128 212084
rect 204812 212032 204864 212084
rect 180524 211964 180576 212016
rect 221740 211964 221792 212016
rect 165712 211896 165764 211948
rect 165896 211896 165948 211948
rect 172060 211896 172112 211948
rect 213736 211896 213788 211948
rect 155224 211828 155276 211880
rect 204076 211828 204128 211880
rect 28264 211760 28316 211812
rect 202696 211760 202748 211812
rect 203708 211760 203760 211812
rect 272064 211760 272116 211812
rect 167644 211692 167696 211744
rect 168288 211692 168340 211744
rect 178592 211692 178644 211744
rect 185860 211692 185912 211744
rect 195980 211692 196032 211744
rect 196164 211692 196216 211744
rect 168748 211352 168800 211404
rect 169668 211352 169720 211404
rect 187332 211352 187384 211404
rect 187792 211352 187844 211404
rect 202144 211352 202196 211404
rect 169760 211284 169812 211336
rect 173532 211284 173584 211336
rect 178684 211284 178736 211336
rect 203708 211284 203760 211336
rect 162584 211216 162636 211268
rect 166540 211216 166592 211268
rect 168288 211216 168340 211268
rect 196256 211216 196308 211268
rect 157892 211148 157944 211200
rect 202328 211148 202380 211200
rect 197360 211080 197412 211132
rect 197544 211080 197596 211132
rect 179604 210876 179656 210928
rect 179788 210876 179840 210928
rect 200212 210808 200264 210860
rect 201132 210808 201184 210860
rect 184940 210740 184992 210792
rect 185216 210740 185268 210792
rect 3516 210536 3568 210588
rect 178684 210536 178736 210588
rect 183100 210536 183152 210588
rect 213184 210536 213236 210588
rect 3424 210468 3476 210520
rect 184388 210468 184440 210520
rect 3608 210400 3660 210452
rect 187792 210400 187844 210452
rect 205272 210400 205324 210452
rect 218796 210400 218848 210452
rect 198372 209992 198424 210044
rect 204352 209992 204404 210044
rect 205364 209992 205416 210044
rect 160560 209924 160612 209976
rect 200212 209924 200264 209976
rect 156604 209856 156656 209908
rect 153844 209788 153896 209840
rect 198372 209788 198424 209840
rect 199568 209856 199620 209908
rect 199936 209856 199988 209908
rect 204260 209788 204312 209840
rect 159456 209380 159508 209432
rect 163596 209380 163648 209432
rect 160652 209176 160704 209228
rect 201684 209380 201736 209432
rect 146944 209108 146996 209160
rect 203156 209516 203208 209568
rect 203892 209516 203944 209568
rect 120816 209040 120868 209092
rect 202880 209448 202932 209500
rect 204996 209380 205048 209432
rect 11704 208360 11756 208412
rect 209320 207680 209372 207732
rect 264520 207680 264572 207732
rect 209412 207612 209464 207664
rect 265808 207612 265860 207664
rect 209596 206320 209648 206372
rect 260288 206320 260340 206372
rect 209504 206252 209556 206304
rect 264428 206252 264480 206304
rect 209688 204960 209740 205012
rect 261668 204960 261720 205012
rect 249800 204892 249852 204944
rect 250444 204892 250496 204944
rect 327264 204824 327316 204876
rect 327816 204824 327868 204876
rect 247960 203600 248012 203652
rect 332600 203600 332652 203652
rect 229008 203532 229060 203584
rect 342260 203532 342312 203584
rect 3332 202784 3384 202836
rect 159272 202784 159324 202836
rect 208952 202104 209004 202156
rect 266728 202104 266780 202156
rect 210516 200744 210568 200796
rect 224592 200744 224644 200796
rect 210700 199384 210752 199436
rect 225144 199384 225196 199436
rect 577504 193128 577556 193180
rect 579620 193128 579672 193180
rect 3148 188980 3200 189032
rect 160560 188980 160612 189032
rect 257528 187688 257580 187740
rect 257804 187688 257856 187740
rect 449900 187688 449952 187740
rect 257620 186328 257672 186380
rect 257988 186328 258040 186380
rect 447140 186328 447192 186380
rect 242624 184152 242676 184204
rect 260840 184152 260892 184204
rect 256240 183540 256292 183592
rect 256516 183540 256568 183592
rect 425060 183540 425112 183592
rect 210332 180072 210384 180124
rect 222292 180072 222344 180124
rect 209228 175924 209280 175976
rect 267188 175924 267240 175976
rect 248236 175244 248288 175296
rect 325700 175244 325752 175296
rect 260288 175176 260340 175228
rect 260748 175176 260800 175228
rect 260288 173884 260340 173936
rect 478880 173884 478932 173936
rect 246764 171096 246816 171148
rect 305000 171096 305052 171148
rect 245016 168376 245068 168428
rect 245292 168376 245344 168428
rect 298100 168376 298152 168428
rect 283656 167016 283708 167068
rect 284116 167016 284168 167068
rect 340880 167016 340932 167068
rect 3332 164160 3384 164212
rect 160652 164160 160704 164212
rect 157800 162256 157852 162308
rect 158076 162256 158128 162308
rect 161664 161508 161716 161560
rect 162400 161508 162452 161560
rect 158720 161100 158772 161152
rect 159640 161100 159692 161152
rect 208400 161372 208452 161424
rect 155868 160624 155920 160676
rect 162124 160624 162176 160676
rect 155500 160420 155552 160472
rect 157064 160216 157116 160268
rect 161848 160148 161900 160200
rect 159916 160012 159968 160064
rect 162124 159944 162176 159996
rect 161756 159876 161808 159928
rect 150440 159808 150492 159860
rect 159548 159808 159600 159860
rect 159916 159808 159968 159860
rect 162676 159876 162728 159928
rect 162952 159876 163004 159928
rect 163320 159876 163372 159928
rect 163136 159808 163188 159860
rect 164148 159808 164200 159860
rect 164424 159808 164476 159860
rect 132500 159740 132552 159792
rect 135260 159672 135312 159724
rect 164700 159740 164752 159792
rect 165344 159740 165396 159792
rect 165528 159876 165580 159928
rect 166172 159808 166224 159860
rect 167736 159876 167788 159928
rect 229560 161236 229612 161288
rect 207940 161168 207992 161220
rect 208308 161168 208360 161220
rect 207480 161100 207532 161152
rect 256148 161100 256200 161152
rect 207940 161032 207992 161084
rect 254860 161032 254912 161084
rect 209228 160964 209280 161016
rect 246304 160964 246356 161016
rect 208400 160896 208452 160948
rect 224500 160896 224552 160948
rect 169760 159876 169812 159928
rect 165620 159740 165672 159792
rect 167552 159740 167604 159792
rect 139400 159604 139452 159656
rect 158444 159604 158496 159656
rect 125600 159536 125652 159588
rect 160008 159604 160060 159656
rect 163044 159604 163096 159656
rect 163688 159604 163740 159656
rect 167460 159672 167512 159724
rect 167736 159672 167788 159724
rect 172704 159808 172756 159860
rect 170956 159740 171008 159792
rect 170680 159672 170732 159724
rect 171232 159672 171284 159724
rect 171784 159672 171836 159724
rect 172888 159740 172940 159792
rect 96620 159468 96672 159520
rect 156880 159468 156932 159520
rect 78680 159400 78732 159452
rect 152648 159400 152700 159452
rect 152924 159400 152976 159452
rect 164424 159536 164476 159588
rect 174084 159808 174136 159860
rect 174820 159808 174872 159860
rect 176384 159876 176436 159928
rect 177672 159876 177724 159928
rect 173900 159740 173952 159792
rect 168288 159536 168340 159588
rect 170680 159536 170732 159588
rect 161296 159468 161348 159520
rect 173256 159604 173308 159656
rect 173992 159604 174044 159656
rect 174268 159604 174320 159656
rect 171692 159536 171744 159588
rect 178960 159740 179012 159792
rect 227444 160760 227496 160812
rect 230112 160692 230164 160744
rect 186504 159876 186556 159928
rect 209228 160216 209280 160268
rect 192024 159876 192076 159928
rect 193772 159876 193824 159928
rect 199660 159876 199712 159928
rect 200672 159876 200724 159928
rect 207940 160080 207992 160132
rect 209596 160148 209648 160200
rect 208952 159944 209004 159996
rect 206468 159876 206520 159928
rect 206744 159876 206796 159928
rect 208768 159876 208820 159928
rect 205916 159808 205968 159860
rect 207664 159808 207716 159860
rect 197912 159740 197964 159792
rect 198556 159740 198608 159792
rect 199384 159740 199436 159792
rect 203524 159740 203576 159792
rect 203800 159740 203852 159792
rect 209044 159740 209096 159792
rect 207756 159672 207808 159724
rect 158536 159400 158588 159452
rect 165528 159400 165580 159452
rect 166908 159400 166960 159452
rect 167184 159400 167236 159452
rect 169576 159400 169628 159452
rect 175096 159468 175148 159520
rect 185400 159604 185452 159656
rect 208584 159604 208636 159656
rect 182548 159536 182600 159588
rect 242164 159536 242216 159588
rect 178960 159468 179012 159520
rect 3700 159332 3752 159384
rect 157892 159332 157944 159384
rect 159916 159332 159968 159384
rect 173256 159400 173308 159452
rect 154396 159196 154448 159248
rect 164240 159264 164292 159316
rect 165344 159264 165396 159316
rect 172612 159332 172664 159384
rect 173164 159332 173216 159384
rect 181720 159332 181772 159384
rect 190184 159468 190236 159520
rect 211804 159468 211856 159520
rect 195428 159400 195480 159452
rect 219256 159400 219308 159452
rect 210240 159332 210292 159384
rect 161204 159196 161256 159248
rect 161572 159128 161624 159180
rect 162584 159128 162636 159180
rect 164424 159196 164476 159248
rect 167368 159264 167420 159316
rect 167736 159264 167788 159316
rect 166540 159196 166592 159248
rect 201316 159264 201368 159316
rect 208860 159264 208912 159316
rect 153016 159060 153068 159112
rect 161848 159060 161900 159112
rect 152740 158992 152792 159044
rect 168932 159060 168984 159112
rect 171048 159128 171100 159180
rect 176200 159060 176252 159112
rect 176844 159060 176896 159112
rect 178960 159060 179012 159112
rect 152924 158924 152976 158976
rect 168564 158992 168616 159044
rect 170772 158992 170824 159044
rect 163136 158924 163188 158976
rect 163412 158924 163464 158976
rect 164332 158924 164384 158976
rect 165252 158924 165304 158976
rect 167184 158924 167236 158976
rect 169944 158924 169996 158976
rect 171508 158924 171560 158976
rect 172060 158924 172112 158976
rect 175096 158924 175148 158976
rect 161388 158856 161440 158908
rect 178224 158856 178276 158908
rect 161940 158788 161992 158840
rect 176016 158788 176068 158840
rect 164148 158720 164200 158772
rect 164424 158720 164476 158772
rect 164700 158720 164752 158772
rect 166816 158720 166868 158772
rect 154304 158652 154356 158704
rect 163780 158584 163832 158636
rect 163044 158516 163096 158568
rect 164332 158652 164384 158704
rect 164608 158584 164660 158636
rect 165528 158584 165580 158636
rect 172152 158720 172204 158772
rect 169208 158584 169260 158636
rect 169760 158584 169812 158636
rect 164332 158516 164384 158568
rect 172796 158652 172848 158704
rect 173440 158652 173492 158704
rect 176568 158584 176620 158636
rect 176844 158584 176896 158636
rect 162308 158448 162360 158500
rect 168288 158448 168340 158500
rect 172980 158516 173032 158568
rect 151176 158380 151228 158432
rect 151636 158380 151688 158432
rect 165620 158380 165672 158432
rect 167368 158380 167420 158432
rect 170588 158380 170640 158432
rect 153936 158312 153988 158364
rect 164332 158312 164384 158364
rect 165896 158312 165948 158364
rect 166356 158312 166408 158364
rect 176844 158448 176896 158500
rect 177120 158584 177172 158636
rect 190828 159128 190880 159180
rect 191288 159128 191340 159180
rect 195520 159128 195572 159180
rect 200672 159128 200724 159180
rect 203800 159196 203852 159248
rect 204536 159196 204588 159248
rect 201316 159128 201368 159180
rect 202328 159128 202380 159180
rect 203432 159128 203484 159180
rect 205088 159128 205140 159180
rect 205548 159128 205600 159180
rect 206744 159128 206796 159180
rect 207480 159128 207532 159180
rect 207756 159128 207808 159180
rect 209228 159128 209280 159180
rect 264244 159128 264296 159180
rect 181720 159060 181772 159112
rect 232872 159060 232924 159112
rect 181904 158992 181956 159044
rect 232504 158992 232556 159044
rect 229928 158924 229980 158976
rect 184204 158856 184256 158908
rect 243636 158856 243688 158908
rect 182364 158720 182416 158772
rect 183284 158720 183336 158772
rect 183652 158720 183704 158772
rect 184204 158720 184256 158772
rect 189356 158788 189408 158840
rect 189632 158788 189684 158840
rect 196164 158788 196216 158840
rect 197176 158788 197228 158840
rect 198556 158788 198608 158840
rect 199660 158788 199712 158840
rect 200672 158788 200724 158840
rect 256240 158788 256292 158840
rect 231492 158720 231544 158772
rect 182272 158652 182324 158704
rect 183468 158652 183520 158704
rect 184388 158652 184440 158704
rect 186320 158652 186372 158704
rect 188252 158652 188304 158704
rect 189356 158652 189408 158704
rect 189908 158652 189960 158704
rect 194416 158652 194468 158704
rect 195152 158652 195204 158704
rect 196624 158652 196676 158704
rect 200028 158652 200080 158704
rect 202328 158652 202380 158704
rect 202880 158652 202932 158704
rect 203340 158652 203392 158704
rect 184756 158584 184808 158636
rect 186872 158584 186924 158636
rect 188528 158584 188580 158636
rect 194324 158584 194376 158636
rect 203524 158584 203576 158636
rect 187148 158516 187200 158568
rect 189908 158516 189960 158568
rect 190184 158516 190236 158568
rect 201316 158516 201368 158568
rect 177120 158448 177172 158500
rect 177396 158448 177448 158500
rect 182732 158448 182784 158500
rect 188252 158448 188304 158500
rect 188344 158448 188396 158500
rect 191196 158448 191248 158500
rect 196532 158448 196584 158500
rect 206744 158652 206796 158704
rect 207204 158652 207256 158704
rect 251824 158652 251876 158704
rect 203800 158584 203852 158636
rect 204168 158584 204220 158636
rect 204812 158584 204864 158636
rect 209504 158584 209556 158636
rect 204260 158516 204312 158568
rect 209320 158516 209372 158568
rect 203708 158448 203760 158500
rect 247684 158448 247736 158500
rect 172612 158380 172664 158432
rect 148324 158244 148376 158296
rect 160560 158244 160612 158296
rect 162216 158244 162268 158296
rect 171692 158312 171744 158364
rect 172060 158312 172112 158364
rect 174636 158312 174688 158364
rect 175556 158312 175608 158364
rect 166724 158244 166776 158296
rect 172336 158244 172388 158296
rect 124864 158108 124916 158160
rect 163964 158108 164016 158160
rect 60740 158040 60792 158092
rect 166908 158176 166960 158228
rect 168288 158176 168340 158228
rect 172428 158176 172480 158228
rect 171232 158108 171284 158160
rect 171508 158108 171560 158160
rect 169760 158040 169812 158092
rect 170128 158040 170180 158092
rect 172612 158040 172664 158092
rect 186320 158244 186372 158296
rect 192024 158244 192076 158296
rect 177396 158176 177448 158228
rect 177672 158176 177724 158228
rect 184112 158176 184164 158228
rect 198004 158176 198056 158228
rect 181352 158108 181404 158160
rect 190276 158108 190328 158160
rect 191012 158108 191064 158160
rect 180524 158040 180576 158092
rect 191104 158040 191156 158092
rect 46204 157972 46256 158024
rect 161480 157972 161532 158024
rect 162768 157972 162820 158024
rect 163504 157972 163556 158024
rect 174268 157972 174320 158024
rect 180248 157972 180300 158024
rect 190184 157972 190236 158024
rect 156696 157904 156748 157956
rect 165160 157904 165212 157956
rect 168932 157904 168984 157956
rect 169300 157904 169352 157956
rect 169484 157904 169536 157956
rect 176108 157904 176160 157956
rect 178960 157904 179012 157956
rect 184112 157904 184164 157956
rect 184756 157904 184808 157956
rect 186504 157904 186556 157956
rect 160836 157836 160888 157888
rect 164240 157836 164292 157888
rect 165344 157836 165396 157888
rect 177120 157836 177172 157888
rect 193496 158108 193548 158160
rect 192668 158040 192720 158092
rect 196348 158040 196400 158092
rect 192116 157972 192168 158024
rect 194140 157972 194192 158024
rect 191564 157904 191616 157956
rect 195612 157836 195664 157888
rect 162032 157768 162084 157820
rect 179052 157768 179104 157820
rect 185216 157768 185268 157820
rect 190184 157768 190236 157820
rect 190276 157768 190328 157820
rect 195428 157768 195480 157820
rect 161020 157700 161072 157752
rect 176844 157700 176896 157752
rect 177672 157700 177724 157752
rect 188252 157700 188304 157752
rect 195336 157700 195388 157752
rect 197360 157836 197412 157888
rect 200212 157836 200264 157888
rect 201776 158380 201828 158432
rect 209688 158380 209740 158432
rect 200948 158312 201000 158364
rect 210700 158312 210752 158364
rect 207480 158244 207532 158296
rect 252008 158244 252060 158296
rect 207572 158176 207624 158228
rect 252100 158176 252152 158228
rect 207020 158108 207072 158160
rect 253204 158108 253256 158160
rect 207848 158040 207900 158092
rect 207940 158040 207992 158092
rect 208308 158040 208360 158092
rect 208400 158040 208452 158092
rect 272248 158040 272300 158092
rect 200672 157972 200724 158024
rect 201224 157972 201276 158024
rect 209688 157972 209740 158024
rect 283656 157972 283708 158024
rect 307116 157972 307168 158024
rect 324412 157972 324464 158024
rect 205180 157836 205232 157888
rect 207112 157904 207164 157956
rect 249340 157904 249392 157956
rect 208032 157836 208084 157888
rect 199292 157768 199344 157820
rect 200120 157768 200172 157820
rect 204168 157700 204220 157752
rect 160744 157632 160796 157684
rect 165344 157632 165396 157684
rect 160928 157564 160980 157616
rect 177488 157632 177540 157684
rect 195704 157632 195756 157684
rect 199476 157632 199528 157684
rect 200212 157632 200264 157684
rect 208124 157768 208176 157820
rect 163688 157496 163740 157548
rect 170220 157564 170272 157616
rect 176568 157564 176620 157616
rect 182732 157564 182784 157616
rect 191104 157564 191156 157616
rect 198188 157564 198240 157616
rect 198280 157564 198332 157616
rect 258908 157700 258960 157752
rect 166356 157496 166408 157548
rect 200948 157496 201000 157548
rect 163504 157428 163556 157480
rect 166724 157428 166776 157480
rect 171784 157428 171836 157480
rect 157984 157360 158036 157412
rect 162860 157360 162912 157412
rect 164148 157360 164200 157412
rect 164240 157360 164292 157412
rect 169484 157360 169536 157412
rect 185768 157428 185820 157480
rect 187240 157428 187292 157480
rect 189632 157428 189684 157480
rect 192668 157428 192720 157480
rect 195980 157428 196032 157480
rect 255412 157632 255464 157684
rect 207296 157428 207348 157480
rect 250444 157428 250496 157480
rect 207940 157360 207992 157412
rect 204168 157292 204220 157344
rect 207204 157292 207256 157344
rect 154488 157224 154540 157276
rect 164976 157224 165028 157276
rect 208584 157224 208636 157276
rect 270776 157224 270828 157276
rect 271788 157224 271840 157276
rect 162124 157156 162176 157208
rect 162860 157156 162912 157208
rect 172980 157156 173032 157208
rect 233516 157156 233568 157208
rect 162216 157088 162268 157140
rect 171600 157088 171652 157140
rect 191104 157088 191156 157140
rect 246580 157088 246632 157140
rect 174360 157020 174412 157072
rect 234160 157020 234212 157072
rect 123484 156952 123536 157004
rect 167644 156952 167696 157004
rect 175740 156952 175792 157004
rect 235448 156952 235500 157004
rect 106280 156884 106332 156936
rect 170680 156884 170732 156936
rect 181076 156884 181128 156936
rect 240140 156884 240192 156936
rect 240968 156884 241020 156936
rect 99380 156816 99432 156868
rect 162124 156816 162176 156868
rect 189356 156816 189408 156868
rect 247960 156816 248012 156868
rect 85580 156748 85632 156800
rect 169024 156748 169076 156800
rect 179604 156748 179656 156800
rect 200856 156748 200908 156800
rect 81440 156680 81492 156732
rect 168748 156680 168800 156732
rect 178500 156680 178552 156732
rect 207756 156680 207808 156732
rect 271788 156680 271840 156732
rect 289084 156680 289136 156732
rect 74540 156612 74592 156664
rect 168196 156612 168248 156664
rect 171140 156612 171192 156664
rect 171508 156612 171560 156664
rect 178776 156612 178828 156664
rect 209504 156612 209556 156664
rect 213644 156612 213696 156664
rect 162124 156544 162176 156596
rect 169760 156544 169812 156596
rect 186044 156544 186096 156596
rect 191104 156544 191156 156596
rect 192944 156476 192996 156528
rect 207020 156544 207072 156596
rect 151728 156408 151780 156460
rect 163504 156408 163556 156460
rect 161388 156340 161440 156392
rect 174912 156340 174964 156392
rect 172888 156272 172940 156324
rect 220544 156476 220596 156528
rect 288532 156612 288584 156664
rect 430580 156612 430632 156664
rect 164240 156204 164292 156256
rect 164976 156204 165028 156256
rect 195796 156204 195848 156256
rect 200856 156272 200908 156324
rect 211804 156272 211856 156324
rect 200120 156136 200172 156188
rect 200948 156136 201000 156188
rect 167184 156068 167236 156120
rect 168104 156068 168156 156120
rect 160744 155932 160796 155984
rect 166356 155932 166408 155984
rect 168656 155932 168708 155984
rect 169116 155932 169168 155984
rect 169944 155932 169996 155984
rect 170312 155932 170364 155984
rect 171232 155932 171284 155984
rect 171876 155932 171928 155984
rect 177120 155932 177172 155984
rect 181444 155932 181496 155984
rect 211804 155932 211856 155984
rect 212264 155932 212316 155984
rect 289360 155932 289412 155984
rect 518900 155932 518952 155984
rect 149704 155864 149756 155916
rect 150348 155864 150400 155916
rect 165068 155864 165120 155916
rect 169300 155864 169352 155916
rect 169668 155864 169720 155916
rect 175464 155864 175516 155916
rect 176384 155864 176436 155916
rect 155776 155728 155828 155780
rect 166632 155728 166684 155780
rect 161848 155660 161900 155712
rect 163228 155660 163280 155712
rect 168472 155660 168524 155712
rect 169208 155660 169260 155712
rect 171140 155660 171192 155712
rect 175740 155660 175792 155712
rect 187516 155864 187568 155916
rect 210608 155864 210660 155916
rect 203064 155796 203116 155848
rect 282276 155796 282328 155848
rect 282552 155796 282604 155848
rect 178040 155728 178092 155780
rect 201500 155728 201552 155780
rect 207204 155728 207256 155780
rect 207756 155728 207808 155780
rect 215944 155728 215996 155780
rect 235264 155660 235316 155712
rect 164792 155592 164844 155644
rect 175188 155592 175240 155644
rect 219072 155592 219124 155644
rect 173348 155524 173400 155576
rect 173532 155524 173584 155576
rect 215760 155524 215812 155576
rect 176292 155456 176344 155508
rect 178040 155456 178092 155508
rect 180156 155456 180208 155508
rect 220636 155456 220688 155508
rect 225604 155456 225656 155508
rect 252560 155456 252612 155508
rect 253204 155456 253256 155508
rect 153200 155388 153252 155440
rect 174360 155388 174412 155440
rect 202604 155388 202656 155440
rect 237012 155388 237064 155440
rect 144920 155320 144972 155372
rect 173716 155320 173768 155372
rect 179328 155320 179380 155372
rect 210332 155320 210384 155372
rect 25504 155252 25556 155304
rect 164332 155252 164384 155304
rect 198004 155252 198056 155304
rect 221832 155252 221884 155304
rect 6920 155184 6972 155236
rect 155868 155184 155920 155236
rect 155960 155184 156012 155236
rect 174544 155184 174596 155236
rect 178040 155184 178092 155236
rect 216312 155184 216364 155236
rect 282276 155184 282328 155236
rect 522304 155184 522356 155236
rect 190736 155116 190788 155168
rect 202144 155116 202196 155168
rect 203616 155116 203668 155168
rect 204076 155116 204128 155168
rect 183744 155048 183796 155100
rect 271144 155048 271196 155100
rect 179880 154980 179932 155032
rect 212448 154980 212500 155032
rect 182456 154912 182508 154964
rect 252560 154912 252612 154964
rect 188804 154844 188856 154896
rect 207112 154844 207164 154896
rect 167552 154776 167604 154828
rect 168288 154776 168340 154828
rect 177672 154776 177724 154828
rect 180064 154776 180116 154828
rect 212448 154572 212500 154624
rect 213184 154572 213236 154624
rect 275652 154572 275704 154624
rect 494060 154572 494112 154624
rect 192392 154504 192444 154556
rect 207572 154504 207624 154556
rect 178316 154368 178368 154420
rect 200856 154436 200908 154488
rect 205824 154436 205876 154488
rect 282276 154436 282328 154488
rect 197452 154368 197504 154420
rect 197912 154368 197964 154420
rect 202052 154368 202104 154420
rect 277400 154368 277452 154420
rect 175832 154300 175884 154352
rect 176568 154300 176620 154352
rect 235632 154300 235684 154352
rect 173440 154232 173492 154284
rect 173716 154232 173768 154284
rect 228548 154232 228600 154284
rect 182916 154164 182968 154216
rect 233148 154164 233200 154216
rect 182180 154096 182232 154148
rect 183192 154096 183244 154148
rect 187976 154096 188028 154148
rect 238208 154096 238260 154148
rect 175004 154028 175056 154080
rect 217324 154028 217376 154080
rect 138020 153960 138072 154012
rect 172520 153960 172572 154012
rect 185492 153960 185544 154012
rect 223304 153960 223356 154012
rect 92480 153892 92532 153944
rect 169576 153892 169628 153944
rect 180616 153892 180668 153944
rect 214564 153892 214616 153944
rect 57980 153824 58032 153876
rect 156788 153824 156840 153876
rect 178592 153824 178644 153876
rect 208400 153824 208452 153876
rect 209596 153824 209648 153876
rect 269120 154096 269172 154148
rect 270132 154096 270184 154148
rect 250444 153824 250496 153876
rect 282276 153824 282328 153876
rect 557540 153824 557592 153876
rect 189080 153756 189132 153808
rect 202880 153756 202932 153808
rect 180708 153688 180760 153740
rect 220728 153688 220780 153740
rect 228364 153688 228416 153740
rect 183836 153620 183888 153672
rect 276296 153620 276348 153672
rect 195612 153552 195664 153604
rect 207296 153552 207348 153604
rect 184940 153416 184992 153468
rect 185860 153416 185912 153468
rect 197636 153348 197688 153400
rect 198004 153348 198056 153400
rect 296628 153280 296680 153332
rect 507860 153280 507912 153332
rect 205732 153212 205784 153264
rect 206008 153212 206060 153264
rect 206192 153212 206244 153264
rect 206652 153212 206704 153264
rect 172612 153144 172664 153196
rect 176568 153144 176620 153196
rect 202236 153144 202288 153196
rect 202604 153144 202656 153196
rect 205640 153144 205692 153196
rect 206376 153144 206428 153196
rect 175464 153076 175516 153128
rect 176476 153076 176528 153128
rect 189264 153076 189316 153128
rect 189632 153076 189684 153128
rect 205272 153076 205324 153128
rect 270132 153212 270184 153264
rect 483020 153212 483072 153264
rect 217324 153144 217376 153196
rect 217784 153144 217836 153196
rect 280436 153144 280488 153196
rect 579896 153144 579948 153196
rect 287980 153076 288032 153128
rect 288348 153076 288400 153128
rect 188896 153008 188948 153060
rect 209688 153008 209740 153060
rect 209780 153008 209832 153060
rect 218980 153008 219032 153060
rect 175280 152940 175332 152992
rect 176016 152940 176068 152992
rect 187700 152940 187752 152992
rect 247776 152940 247828 152992
rect 183284 152872 183336 152924
rect 241336 152872 241388 152924
rect 246304 152872 246356 152924
rect 176752 152804 176804 152856
rect 179328 152804 179380 152856
rect 181812 152804 181864 152856
rect 235356 152804 235408 152856
rect 195980 152736 196032 152788
rect 196992 152736 197044 152788
rect 197176 152736 197228 152788
rect 239588 152736 239640 152788
rect 174636 152668 174688 152720
rect 133880 152600 133932 152652
rect 173716 152600 173768 152652
rect 186320 152600 186372 152652
rect 187332 152600 187384 152652
rect 190552 152600 190604 152652
rect 215116 152668 215168 152720
rect 104900 152532 104952 152584
rect 170864 152532 170916 152584
rect 46940 152464 46992 152516
rect 155592 152464 155644 152516
rect 165804 152464 165856 152516
rect 166448 152464 166500 152516
rect 163228 152396 163280 152448
rect 163780 152396 163832 152448
rect 176660 152464 176712 152516
rect 177028 152464 177080 152516
rect 177304 152464 177356 152516
rect 177948 152464 178000 152516
rect 179512 152532 179564 152584
rect 180432 152532 180484 152584
rect 180984 152532 181036 152584
rect 176936 152396 176988 152448
rect 177764 152396 177816 152448
rect 173256 152328 173308 152380
rect 173808 152328 173860 152380
rect 180892 152464 180944 152516
rect 181996 152464 182048 152516
rect 182180 152464 182232 152516
rect 182732 152464 182784 152516
rect 183744 152464 183796 152516
rect 184572 152464 184624 152516
rect 186504 152532 186556 152584
rect 186964 152532 187016 152584
rect 187700 152532 187752 152584
rect 188712 152532 188764 152584
rect 189080 152532 189132 152584
rect 190368 152532 190420 152584
rect 194600 152532 194652 152584
rect 194876 152532 194928 152584
rect 207848 152600 207900 152652
rect 307116 152600 307168 152652
rect 228732 152532 228784 152584
rect 217324 152464 217376 152516
rect 181168 152396 181220 152448
rect 181904 152396 181956 152448
rect 183652 152396 183704 152448
rect 184848 152396 184900 152448
rect 184940 152396 184992 152448
rect 186228 152396 186280 152448
rect 186596 152396 186648 152448
rect 187056 152396 187108 152448
rect 187792 152396 187844 152448
rect 188436 152396 188488 152448
rect 189172 152396 189224 152448
rect 189816 152396 189868 152448
rect 190644 152396 190696 152448
rect 190920 152396 190972 152448
rect 191932 152396 191984 152448
rect 192852 152396 192904 152448
rect 196164 152396 196216 152448
rect 196440 152396 196492 152448
rect 197452 152396 197504 152448
rect 197820 152396 197872 152448
rect 198740 152396 198792 152448
rect 199384 152396 199436 152448
rect 200120 152396 200172 152448
rect 200580 152396 200632 152448
rect 201684 152396 201736 152448
rect 202512 152396 202564 152448
rect 202604 152396 202656 152448
rect 284392 152396 284444 152448
rect 512000 152532 512052 152584
rect 288348 152464 288400 152516
rect 550640 152464 550692 152516
rect 234068 152328 234120 152380
rect 179512 152260 179564 152312
rect 179972 152260 180024 152312
rect 180156 152260 180208 152312
rect 165620 152192 165672 152244
rect 166540 152192 166592 152244
rect 178684 152192 178736 152244
rect 179420 152124 179472 152176
rect 179696 152124 179748 152176
rect 186504 152124 186556 152176
rect 187608 152124 187660 152176
rect 192208 152124 192260 152176
rect 193128 152124 193180 152176
rect 193496 152124 193548 152176
rect 194048 152124 194100 152176
rect 177764 152056 177816 152108
rect 180156 152056 180208 152108
rect 193220 152056 193272 152108
rect 193864 152056 193916 152108
rect 197636 152192 197688 152244
rect 198648 152192 198700 152244
rect 201776 152192 201828 152244
rect 202788 152192 202840 152244
rect 205916 152260 205968 152312
rect 206192 152260 206244 152312
rect 209872 152260 209924 152312
rect 210884 152260 210936 152312
rect 211988 152192 212040 152244
rect 209872 152056 209924 152108
rect 193312 151988 193364 152040
rect 194232 151988 194284 152040
rect 205640 151988 205692 152040
rect 206928 151988 206980 152040
rect 194692 151784 194744 151836
rect 195060 151784 195112 151836
rect 159732 151716 159784 151768
rect 161480 151716 161532 151768
rect 181260 151716 181312 151768
rect 214380 151716 214432 151768
rect 215208 151716 215260 151768
rect 186688 151648 186740 151700
rect 213552 151648 213604 151700
rect 182640 151580 182692 151632
rect 242716 151580 242768 151632
rect 185676 151512 185728 151564
rect 245384 151512 245436 151564
rect 181628 151444 181680 151496
rect 240784 151444 240836 151496
rect 183560 151376 183612 151428
rect 243544 151376 243596 151428
rect 189908 151308 189960 151360
rect 247868 151308 247920 151360
rect 188528 151240 188580 151292
rect 246488 151240 246540 151292
rect 180800 151172 180852 151224
rect 236000 151172 236052 151224
rect 151084 151104 151136 151156
rect 174084 151104 174136 151156
rect 195428 151104 195480 151156
rect 241520 151104 241572 151156
rect 245384 151104 245436 151156
rect 295984 151104 296036 151156
rect 142160 151036 142212 151088
rect 172704 151036 172756 151088
rect 198188 151036 198240 151088
rect 233240 151036 233292 151088
rect 279700 151036 279752 151088
rect 381636 151036 381688 151088
rect 201224 150968 201276 151020
rect 229100 150968 229152 151020
rect 229836 150968 229888 151020
rect 183192 150900 183244 150952
rect 251272 150900 251324 150952
rect 192300 150832 192352 150884
rect 279700 150832 279752 150884
rect 236000 150492 236052 150544
rect 236920 150492 236972 150544
rect 214380 150424 214432 150476
rect 215944 150424 215996 150476
rect 233240 150424 233292 150476
rect 233976 150424 234028 150476
rect 241520 150424 241572 150476
rect 242164 150424 242216 150476
rect 242716 150424 242768 150476
rect 243636 150424 243688 150476
rect 251272 150424 251324 150476
rect 251824 150424 251876 150476
rect 197360 150356 197412 150408
rect 292212 150356 292264 150408
rect 201500 150288 201552 150340
rect 214656 150288 214708 150340
rect 184020 150220 184072 150272
rect 274456 150220 274508 150272
rect 188068 150152 188120 150204
rect 275192 150152 275244 150204
rect 195336 150084 195388 150136
rect 260840 150084 260892 150136
rect 274640 150084 274692 150136
rect 274916 150084 274968 150136
rect 190184 150016 190236 150068
rect 244924 150016 244976 150068
rect 181536 149948 181588 150000
rect 219440 149948 219492 150000
rect 220728 149948 220780 150000
rect 200856 149880 200908 149932
rect 238392 149880 238444 149932
rect 178868 149812 178920 149864
rect 211068 149812 211120 149864
rect 191840 149744 191892 149796
rect 223212 149744 223264 149796
rect 275192 149744 275244 149796
rect 327080 149744 327132 149796
rect 71780 149676 71832 149728
rect 156880 149676 156932 149728
rect 176568 149676 176620 149728
rect 182088 149676 182140 149728
rect 217508 149676 217560 149728
rect 220728 149676 220780 149728
rect 232504 149676 232556 149728
rect 292212 149676 292264 149728
rect 451280 149676 451332 149728
rect 187240 149608 187292 149660
rect 216220 149608 216272 149660
rect 185860 149540 185912 149592
rect 218888 149540 218940 149592
rect 183008 149472 183060 149524
rect 274640 149472 274692 149524
rect 151820 149064 151872 149116
rect 174176 149064 174228 149116
rect 206008 149064 206060 149116
rect 206560 149064 206612 149116
rect 274456 149064 274508 149116
rect 275100 149064 275152 149116
rect 202880 148996 202932 149048
rect 228824 148996 228876 149048
rect 201408 148928 201460 148980
rect 270040 148928 270092 148980
rect 270316 148928 270368 148980
rect 202328 148860 202380 148912
rect 269120 148860 269172 148912
rect 184388 148792 184440 148844
rect 244096 148792 244148 148844
rect 187976 148724 188028 148776
rect 248052 148724 248104 148776
rect 184664 148656 184716 148708
rect 243728 148656 243780 148708
rect 278044 148656 278096 148708
rect 185584 148588 185636 148640
rect 245016 148588 245068 148640
rect 151912 148520 151964 148572
rect 173900 148520 173952 148572
rect 191196 148520 191248 148572
rect 249248 148520 249300 148572
rect 133144 148452 133196 148504
rect 171968 148452 172020 148504
rect 191288 148452 191340 148504
rect 191564 148452 191616 148504
rect 194140 148452 194192 148504
rect 251916 148452 251968 148504
rect 82820 148384 82872 148436
rect 152832 148384 152884 148436
rect 192668 148384 192720 148436
rect 249156 148384 249208 148436
rect 281540 148384 281592 148436
rect 345020 148384 345072 148436
rect 15844 148316 15896 148368
rect 163412 148316 163464 148368
rect 191380 148316 191432 148368
rect 249432 148316 249484 148368
rect 270316 148316 270368 148368
rect 500960 148316 501012 148368
rect 174176 148248 174228 148300
rect 227352 148248 227404 148300
rect 194416 148180 194468 148232
rect 227168 148180 227220 148232
rect 189632 148112 189684 148164
rect 281540 148112 281592 148164
rect 200856 148044 200908 148096
rect 201408 148044 201460 148096
rect 173900 147636 173952 147688
rect 175372 147636 175424 147688
rect 176844 147568 176896 147620
rect 182824 147568 182876 147620
rect 201960 147568 202012 147620
rect 296628 147568 296680 147620
rect 187884 147500 187936 147552
rect 276112 147500 276164 147552
rect 276388 147500 276440 147552
rect 206100 147432 206152 147484
rect 284300 147432 284352 147484
rect 182364 147364 182416 147416
rect 243452 147364 243504 147416
rect 249432 147364 249484 147416
rect 249708 147364 249760 147416
rect 273260 147364 273312 147416
rect 193496 147296 193548 147348
rect 254676 147296 254728 147348
rect 143540 147024 143592 147076
rect 173624 147228 173676 147280
rect 233332 147228 233384 147280
rect 193956 147160 194008 147212
rect 253756 147160 253808 147212
rect 193588 147092 193640 147144
rect 253480 147092 253532 147144
rect 194876 147024 194928 147076
rect 254584 147024 254636 147076
rect 68284 146956 68336 147008
rect 151268 146956 151320 147008
rect 164884 146956 164936 147008
rect 165252 146956 165304 147008
rect 165896 146956 165948 147008
rect 166264 146956 166316 147008
rect 276388 147024 276440 147076
rect 316684 147024 316736 147076
rect 14464 146888 14516 146940
rect 161664 146888 161716 146940
rect 405740 146956 405792 147008
rect 225420 146888 225472 146940
rect 243452 146888 243504 146940
rect 253296 146888 253348 146940
rect 284300 146888 284352 146940
rect 285128 146888 285180 146940
rect 561680 146888 561732 146940
rect 181812 146820 181864 146872
rect 239404 146820 239456 146872
rect 203708 146752 203760 146804
rect 253572 146752 253624 146804
rect 202236 146684 202288 146736
rect 250628 146684 250680 146736
rect 196256 146616 196308 146668
rect 255964 146616 256016 146668
rect 154212 146208 154264 146260
rect 154488 146208 154540 146260
rect 169300 146208 169352 146260
rect 175556 146208 175608 146260
rect 176108 146208 176160 146260
rect 201684 146208 201736 146260
rect 293960 146208 294012 146260
rect 294604 146208 294656 146260
rect 201776 146140 201828 146192
rect 289360 146140 289412 146192
rect 190736 146072 190788 146124
rect 270316 146072 270368 146124
rect 183744 146004 183796 146056
rect 245476 146004 245528 146056
rect 189448 145936 189500 145988
rect 250904 145936 250956 145988
rect 185308 145868 185360 145920
rect 246672 145868 246724 145920
rect 176108 145800 176160 145852
rect 236092 145800 236144 145852
rect 282184 145800 282236 145852
rect 198004 145732 198056 145784
rect 257344 145732 257396 145784
rect 118700 145664 118752 145716
rect 172060 145664 172112 145716
rect 198832 145664 198884 145716
rect 258172 145664 258224 145716
rect 270316 145664 270368 145716
rect 359464 145664 359516 145716
rect 95884 145596 95936 145648
rect 154488 145596 154540 145648
rect 88984 145528 89036 145580
rect 168656 145528 168708 145580
rect 226984 145596 227036 145648
rect 250904 145596 250956 145648
rect 356060 145596 356112 145648
rect 200856 145528 200908 145580
rect 258724 145528 258776 145580
rect 293960 145528 294012 145580
rect 514024 145528 514076 145580
rect 179696 145460 179748 145512
rect 218060 145460 218112 145512
rect 179328 145392 179380 145444
rect 213276 145392 213328 145444
rect 175464 144848 175516 144900
rect 176568 144848 176620 144900
rect 202880 144848 202932 144900
rect 204076 144848 204128 144900
rect 218060 144848 218112 144900
rect 227076 144848 227128 144900
rect 185216 144780 185268 144832
rect 278228 144780 278280 144832
rect 284944 144780 284996 144832
rect 189356 144712 189408 144764
rect 280252 144712 280304 144764
rect 281448 144712 281500 144764
rect 203892 144644 203944 144696
rect 268936 144644 268988 144696
rect 201132 144576 201184 144628
rect 259828 144576 259880 144628
rect 201224 144508 201276 144560
rect 260104 144508 260156 144560
rect 176200 144440 176252 144492
rect 221464 144440 221516 144492
rect 222016 144440 222068 144492
rect 222200 144440 222252 144492
rect 179604 144372 179656 144424
rect 176568 144304 176620 144356
rect 216036 144304 216088 144356
rect 281448 144304 281500 144356
rect 319444 144304 319496 144356
rect 93860 144236 93912 144288
rect 169116 144236 169168 144288
rect 200304 144236 200356 144288
rect 201224 144236 201276 144288
rect 204076 144236 204128 144288
rect 228640 144236 228692 144288
rect 290924 144236 290976 144288
rect 436744 144236 436796 144288
rect 13084 144168 13136 144220
rect 161572 144168 161624 144220
rect 202696 144168 202748 144220
rect 262404 144168 262456 144220
rect 268936 144168 268988 144220
rect 532700 144168 532752 144220
rect 196164 144100 196216 144152
rect 290648 144100 290700 144152
rect 290924 144100 290976 144152
rect 174636 144032 174688 144084
rect 176200 144032 176252 144084
rect 185124 143488 185176 143540
rect 186228 143488 186280 143540
rect 186688 143488 186740 143540
rect 269212 143488 269264 143540
rect 269304 143488 269356 143540
rect 269764 143488 269816 143540
rect 185032 143420 185084 143472
rect 203616 143352 203668 143404
rect 283104 143352 283156 143404
rect 283564 143352 283616 143404
rect 164516 143284 164568 143336
rect 224316 143284 224368 143336
rect 187792 143216 187844 143268
rect 243820 143216 243872 143268
rect 169760 143148 169812 143200
rect 170128 143148 170180 143200
rect 222936 143148 222988 143200
rect 186228 143080 186280 143132
rect 231124 143080 231176 143132
rect 143632 143012 143684 143064
rect 173348 143012 173400 143064
rect 182272 143012 182324 143064
rect 107660 142944 107712 142996
rect 169760 142944 169812 142996
rect 49700 142876 49752 142928
rect 165712 142876 165764 142928
rect 222108 142876 222160 142928
rect 264244 142876 264296 142928
rect 269212 142876 269264 142928
rect 273444 142876 273496 142928
rect 309876 142876 309928 142928
rect 33140 142808 33192 142860
rect 164240 142808 164292 142860
rect 197084 142808 197136 142860
rect 255320 142808 255372 142860
rect 283104 142808 283156 142860
rect 376024 142808 376076 142860
rect 187700 142060 187752 142112
rect 283012 142060 283064 142112
rect 194784 141992 194836 142044
rect 289176 141992 289228 142044
rect 204352 141924 204404 141976
rect 278136 141924 278188 141976
rect 121460 141516 121512 141568
rect 171232 141856 171284 141908
rect 234620 141856 234672 141908
rect 183652 141788 183704 141840
rect 245200 141788 245252 141840
rect 189264 141720 189316 141772
rect 190368 141720 190420 141772
rect 249064 141720 249116 141772
rect 205824 141652 205876 141704
rect 265348 141652 265400 141704
rect 179144 141584 179196 141636
rect 223120 141584 223172 141636
rect 178224 141516 178276 141568
rect 179052 141516 179104 141568
rect 218704 141516 218756 141568
rect 243820 141516 243872 141568
rect 323584 141516 323636 141568
rect 44180 141448 44232 141500
rect 166264 141448 166316 141500
rect 177580 141448 177632 141500
rect 179236 141448 179288 141500
rect 233884 141448 233936 141500
rect 245200 141448 245252 141500
rect 267004 141448 267056 141500
rect 289176 141448 289228 141500
rect 415400 141448 415452 141500
rect 31024 141380 31076 141432
rect 164516 141380 164568 141432
rect 206928 141380 206980 141432
rect 267924 141380 267976 141432
rect 278136 141380 278188 141432
rect 547144 141380 547196 141432
rect 205916 140836 205968 140888
rect 206928 140836 206980 140888
rect 205824 140768 205876 140820
rect 206468 140768 206520 140820
rect 190644 140700 190696 140752
rect 285036 140700 285088 140752
rect 197636 140632 197688 140684
rect 272616 140632 272668 140684
rect 167276 140564 167328 140616
rect 229468 140564 229520 140616
rect 184940 140496 184992 140548
rect 246856 140496 246908 140548
rect 167368 140428 167420 140480
rect 227260 140428 227312 140480
rect 169944 140360 169996 140412
rect 170404 140360 170456 140412
rect 225696 140360 225748 140412
rect 169760 140292 169812 140344
rect 170036 140292 170088 140344
rect 222844 140292 222896 140344
rect 115204 140156 115256 140208
rect 171876 140156 171928 140208
rect 302884 140156 302936 140208
rect 40040 140088 40092 140140
rect 165160 140088 165212 140140
rect 285036 140088 285088 140140
rect 363604 140088 363656 140140
rect 17224 140020 17276 140072
rect 163504 140020 163556 140072
rect 272616 140020 272668 140072
rect 465080 140020 465132 140072
rect 167276 139408 167328 139460
rect 167644 139408 167696 139460
rect 186596 139340 186648 139392
rect 274824 139340 274876 139392
rect 275376 139340 275428 139392
rect 193404 139272 193456 139324
rect 271972 139272 272024 139324
rect 205088 139204 205140 139256
rect 269028 139204 269080 139256
rect 168104 139136 168156 139188
rect 227996 139136 228048 139188
rect 179512 139068 179564 139120
rect 226248 139068 226300 139120
rect 115940 138796 115992 138848
rect 171324 138796 171376 138848
rect 275376 138796 275428 138848
rect 314016 138796 314068 138848
rect 62120 138728 62172 138780
rect 167368 138728 167420 138780
rect 271972 138728 272024 138780
rect 399484 138728 399536 138780
rect 52460 138660 52512 138712
rect 165804 138660 165856 138712
rect 269028 138660 269080 138712
rect 554780 138660 554832 138712
rect 167736 137980 167788 138032
rect 168104 137980 168156 138032
rect 194692 137912 194744 137964
rect 285772 137912 285824 137964
rect 205732 137844 205784 137896
rect 272248 137844 272300 137896
rect 146300 137300 146352 137352
rect 173256 137300 173308 137352
rect 283012 137300 283064 137352
rect 338120 137300 338172 137352
rect 26240 137232 26292 137284
rect 164424 137232 164476 137284
rect 180432 137232 180484 137284
rect 220084 137232 220136 137284
rect 285772 137232 285824 137284
rect 419540 137232 419592 137284
rect 272248 136620 272300 136672
rect 564440 136620 564492 136672
rect 196992 136552 197044 136604
rect 261576 136552 261628 136604
rect 262128 136552 262180 136604
rect 205640 136484 205692 136536
rect 270868 136484 270920 136536
rect 271788 136484 271840 136536
rect 189172 136416 189224 136468
rect 249616 136416 249668 136468
rect 219440 136348 219492 136400
rect 220084 136348 220136 136400
rect 238024 136348 238076 136400
rect 249616 136008 249668 136060
rect 351920 136008 351972 136060
rect 262128 135940 262180 135992
rect 440240 135940 440292 135992
rect 4804 135872 4856 135924
rect 161756 135872 161808 135924
rect 180524 135872 180576 135924
rect 223580 135872 223632 135924
rect 271788 135872 271840 135924
rect 571984 135872 572036 135924
rect 191564 135192 191616 135244
rect 250996 135192 251048 135244
rect 91100 134580 91152 134632
rect 168380 134580 168432 134632
rect 181904 134580 181956 134632
rect 241520 134580 241572 134632
rect 250996 134580 251048 134632
rect 369860 134580 369912 134632
rect 8300 134512 8352 134564
rect 162860 134512 162912 134564
rect 208124 134512 208176 134564
rect 575480 134512 575532 134564
rect 191472 133832 191524 133884
rect 285680 133832 285732 133884
rect 197452 133764 197504 133816
rect 291936 133764 291988 133816
rect 186320 133696 186372 133748
rect 246028 133696 246080 133748
rect 246028 133288 246080 133340
rect 246948 133288 247000 133340
rect 320180 133288 320232 133340
rect 98000 133220 98052 133272
rect 169760 133220 169812 133272
rect 285680 133220 285732 133272
rect 376760 133220 376812 133272
rect 48320 133152 48372 133204
rect 166172 133152 166224 133204
rect 166264 133152 166316 133204
rect 174728 133152 174780 133204
rect 291936 133152 291988 133204
rect 455420 133152 455472 133204
rect 192024 132404 192076 132456
rect 287796 132404 287848 132456
rect 198924 132336 198976 132388
rect 293224 132336 293276 132388
rect 186504 132268 186556 132320
rect 247040 132268 247092 132320
rect 247040 131860 247092 131912
rect 248328 131860 248380 131912
rect 301504 131860 301556 131912
rect 287796 131792 287848 131844
rect 387800 131792 387852 131844
rect 110512 131724 110564 131776
rect 170864 131724 170916 131776
rect 177764 131724 177816 131776
rect 186320 131724 186372 131776
rect 293224 131724 293276 131776
rect 468484 131724 468536 131776
rect 193312 131044 193364 131096
rect 255228 131044 255280 131096
rect 169024 130364 169076 130416
rect 176108 130364 176160 130416
rect 255228 130364 255280 130416
rect 408500 130364 408552 130416
rect 195704 129684 195756 129736
rect 268200 129684 268252 129736
rect 269028 129684 269080 129736
rect 199660 129616 199712 129668
rect 270408 129616 270460 129668
rect 117320 129072 117372 129124
rect 171784 129072 171836 129124
rect 269028 129072 269080 129124
rect 422944 129072 422996 129124
rect 66260 129004 66312 129056
rect 168288 129004 168340 129056
rect 181996 129004 182048 129056
rect 237380 129004 237432 129056
rect 270408 129004 270460 129056
rect 480260 129004 480312 129056
rect 200120 128256 200172 128308
rect 274088 128256 274140 128308
rect 274548 128256 274600 128308
rect 195980 128188 196032 128240
rect 256056 128188 256108 128240
rect 122104 127644 122156 127696
rect 172428 127644 172480 127696
rect 256056 127644 256108 127696
rect 256608 127644 256660 127696
rect 444380 127644 444432 127696
rect 69020 127576 69072 127628
rect 167736 127576 167788 127628
rect 274088 127576 274140 127628
rect 490012 127576 490064 127628
rect 186412 126896 186464 126948
rect 280804 126896 280856 126948
rect 281448 126896 281500 126948
rect 198556 126828 198608 126880
rect 288440 126828 288492 126880
rect 289728 126828 289780 126880
rect 191932 126760 191984 126812
rect 253480 126760 253532 126812
rect 253848 126760 253900 126812
rect 281448 126352 281500 126404
rect 307852 126352 307904 126404
rect 253480 126284 253532 126336
rect 390560 126284 390612 126336
rect 289728 126216 289780 126268
rect 458180 126216 458232 126268
rect 176568 125536 176620 125588
rect 180156 125536 180208 125588
rect 198740 125536 198792 125588
rect 274732 125536 274784 125588
rect 275376 125536 275428 125588
rect 189080 125468 189132 125520
rect 251088 125468 251140 125520
rect 102140 124924 102192 124976
rect 170404 124924 170456 124976
rect 251088 124924 251140 124976
rect 337384 124924 337436 124976
rect 56600 124856 56652 124908
rect 166080 124856 166132 124908
rect 275376 124856 275428 124908
rect 476120 124856 476172 124908
rect 192944 124108 192996 124160
rect 252468 124108 252520 124160
rect 201592 124040 201644 124092
rect 261484 124040 261536 124092
rect 262128 124040 262180 124092
rect 252468 123496 252520 123548
rect 394700 123496 394752 123548
rect 86960 123428 87012 123480
rect 169484 123428 169536 123480
rect 262128 123428 262180 123480
rect 503720 123428 503772 123480
rect 194508 122068 194560 122120
rect 412640 122068 412692 122120
rect 60832 120708 60884 120760
rect 167092 120708 167144 120760
rect 22744 119348 22796 119400
rect 163228 119348 163280 119400
rect 184572 119348 184624 119400
rect 273260 119348 273312 119400
rect 162860 117988 162912 118040
rect 173992 117988 174044 118040
rect 24124 117920 24176 117972
rect 163044 117920 163096 117972
rect 193220 117240 193272 117292
rect 253388 117240 253440 117292
rect 39304 116560 39356 116612
rect 164700 116560 164752 116612
rect 253388 116560 253440 116612
rect 404360 116560 404412 116612
rect 43444 115200 43496 115252
rect 166816 115200 166868 115252
rect 279424 113092 279476 113144
rect 580172 113092 580224 113144
rect 9680 112412 9732 112464
rect 163412 112412 163464 112464
rect 3148 111732 3200 111784
rect 120816 111732 120868 111784
rect 131120 111052 131172 111104
rect 173072 111052 173124 111104
rect 183468 111052 183520 111104
rect 262220 111052 262272 111104
rect 52552 109692 52604 109744
rect 165620 109692 165672 109744
rect 201132 109692 201184 109744
rect 489184 109692 489236 109744
rect 70400 108264 70452 108316
rect 167460 108264 167512 108316
rect 177304 108264 177356 108316
rect 184296 108264 184348 108316
rect 201224 108264 201276 108316
rect 492680 108264 492732 108316
rect 79324 106904 79376 106956
rect 169208 106904 169260 106956
rect 179052 105612 179104 105664
rect 201592 105612 201644 105664
rect 13820 105544 13872 105596
rect 163136 105544 163188 105596
rect 190368 105544 190420 105596
rect 347780 105544 347832 105596
rect 95240 104116 95292 104168
rect 169852 104116 169904 104168
rect 31760 102756 31812 102808
rect 164608 102756 164660 102808
rect 202696 101396 202748 101448
rect 517520 101396 517572 101448
rect 341524 100648 341576 100700
rect 580172 100648 580224 100700
rect 19340 99968 19392 100020
rect 157892 99968 157944 100020
rect 111800 98608 111852 98660
rect 171508 98608 171560 98660
rect 27620 97248 27672 97300
rect 153936 97248 153988 97300
rect 35900 94460 35952 94512
rect 156696 94460 156748 94512
rect 203984 94460 204036 94512
rect 535460 94460 535512 94512
rect 11060 93100 11112 93152
rect 148324 93100 148376 93152
rect 205548 91740 205600 91792
rect 553400 91740 553452 91792
rect 206560 90312 206612 90364
rect 556252 90312 556304 90364
rect 206468 88952 206520 89004
rect 560300 88952 560352 89004
rect 206652 87592 206704 87644
rect 564532 87592 564584 87644
rect 179144 86232 179196 86284
rect 205640 86232 205692 86284
rect 206744 86232 206796 86284
rect 567200 86232 567252 86284
rect 3516 85484 3568 85536
rect 28264 85484 28316 85536
rect 206836 84804 206888 84856
rect 569224 84804 569276 84856
rect 208216 83444 208268 83496
rect 574100 83444 574152 83496
rect 208308 80656 208360 80708
rect 578240 80656 578292 80708
rect 42800 77936 42852 77988
rect 151176 77936 151228 77988
rect 198648 73788 198700 73840
rect 454040 73788 454092 73840
rect 3516 71680 3568 71732
rect 146944 71680 146996 71732
rect 176660 68280 176712 68332
rect 187700 68280 187752 68332
rect 3056 59304 3108 59356
rect 155224 59304 155276 59356
rect 177948 58624 178000 58676
rect 191104 58624 191156 58676
rect 3516 45500 3568 45552
rect 156604 45500 156656 45552
rect 204168 37884 204220 37936
rect 525800 37884 525852 37936
rect 206928 36524 206980 36576
rect 568580 36524 568632 36576
rect 201316 35164 201368 35216
rect 499580 35164 499632 35216
rect 204076 33736 204128 33788
rect 524420 33736 524472 33788
rect 2872 33056 2924 33108
rect 11704 33056 11756 33108
rect 176016 28908 176068 28960
rect 176660 28908 176712 28960
rect 334624 20612 334676 20664
rect 580080 20612 580132 20664
rect 205456 18572 205508 18624
rect 539692 18572 539744 18624
rect 38660 17212 38712 17264
rect 165436 17212 165488 17264
rect 197176 17212 197228 17264
rect 433340 17212 433392 17264
rect 202788 15852 202840 15904
rect 505376 15852 505428 15904
rect 88892 14424 88944 14476
rect 168932 14424 168984 14476
rect 25320 13064 25372 13116
rect 164884 13064 164936 13116
rect 143540 11772 143592 11824
rect 144736 11772 144788 11824
rect 15752 11704 15804 11756
rect 163780 11704 163832 11756
rect 20168 10276 20220 10328
rect 124864 10276 124916 10328
rect 190460 10276 190512 10328
rect 376024 10276 376076 10328
rect 195888 9052 195940 9104
rect 422576 9052 422628 9104
rect 197084 8984 197136 9036
rect 433248 8984 433300 9036
rect 103336 8916 103388 8968
rect 170772 8916 170824 8968
rect 196072 8916 196124 8968
rect 443828 8916 443880 8968
rect 73804 7556 73856 7608
rect 167644 7556 167696 7608
rect 204260 7556 204312 7608
rect 546684 7556 546736 7608
rect 3424 6808 3476 6860
rect 153844 6808 153896 6860
rect 193128 6264 193180 6316
rect 383568 6264 383620 6316
rect 193036 6196 193088 6248
rect 387156 6196 387208 6248
rect 199844 6128 199896 6180
rect 475752 6128 475804 6180
rect 176292 5516 176344 5568
rect 177856 5516 177908 5568
rect 5264 4768 5316 4820
rect 46204 4768 46256 4820
rect 64328 4768 64380 4820
rect 167920 4768 167972 4820
rect 209688 4088 209740 4140
rect 210976 4088 211028 4140
rect 232504 4088 232556 4140
rect 246396 4088 246448 4140
rect 250444 4088 250496 4140
rect 264152 4088 264204 4140
rect 267004 4088 267056 4140
rect 13544 4020 13596 4072
rect 17224 4020 17276 4072
rect 235264 4020 235316 4072
rect 211804 3952 211856 4004
rect 221556 3952 221608 4004
rect 242808 4020 242860 4072
rect 249984 3952 250036 4004
rect 180156 3884 180208 3936
rect 181444 3884 181496 3936
rect 184296 3884 184348 3936
rect 194416 3884 194468 3936
rect 213184 3884 213236 3936
rect 225144 3884 225196 3936
rect 228364 3884 228416 3936
rect 235816 3884 235868 3936
rect 243636 3884 243688 3936
rect 253112 3884 253164 3936
rect 253296 3952 253348 4004
rect 267648 4020 267700 4072
rect 265348 3952 265400 4004
rect 274640 3952 274692 4004
rect 302884 4088 302936 4140
rect 306748 4088 306800 4140
rect 307024 4088 307076 4140
rect 322112 4088 322164 4140
rect 323584 4088 323636 4140
rect 327540 4088 327592 4140
rect 284944 4020 284996 4072
rect 303160 4020 303212 4072
rect 315304 4020 315356 4072
rect 316224 4020 316276 4072
rect 319444 4020 319496 4072
rect 288992 3952 289044 4004
rect 311164 3952 311216 4004
rect 320824 3952 320876 4004
rect 321100 4020 321152 4072
rect 331588 4088 331640 4140
rect 363604 4088 363656 4140
rect 367008 4088 367060 4140
rect 429844 4088 429896 4140
rect 432052 4088 432104 4140
rect 489184 4088 489236 4140
rect 489920 4088 489972 4140
rect 547144 4088 547196 4140
rect 547880 4088 547932 4140
rect 327816 4020 327868 4072
rect 329288 4020 329340 4072
rect 337384 4020 337436 4072
rect 359924 4020 359976 4072
rect 349160 3952 349212 4004
rect 268844 3884 268896 3936
rect 269764 3884 269816 3936
rect 292580 3884 292632 3936
rect 309784 3884 309836 3936
rect 346952 3884 347004 3936
rect 381636 3884 381688 3936
rect 384764 3884 384816 3936
rect 180064 3816 180116 3868
rect 189724 3816 189776 3868
rect 214564 3816 214616 3868
rect 232228 3816 232280 3868
rect 243544 3816 243596 3868
rect 272432 3816 272484 3868
rect 301504 3816 301556 3868
rect 324320 3816 324372 3868
rect 327724 3816 327776 3868
rect 329196 3816 329248 3868
rect 329288 3816 329340 3868
rect 368204 3816 368256 3868
rect 384304 3816 384356 3868
rect 398840 3816 398892 3868
rect 186964 3748 187016 3800
rect 203892 3748 203944 3800
rect 217324 3748 217376 3800
rect 239312 3748 239364 3800
rect 243728 3748 243780 3800
rect 286600 3748 286652 3800
rect 313924 3748 313976 3800
rect 403624 3748 403676 3800
rect 123484 3680 123536 3732
rect 133144 3680 133196 3732
rect 135260 3680 135312 3732
rect 136456 3680 136508 3732
rect 186044 3680 186096 3732
rect 291384 3680 291436 3732
rect 305644 3680 305696 3732
rect 311440 3680 311492 3732
rect 314016 3680 314068 3732
rect 317328 3680 317380 3732
rect 320824 3680 320876 3732
rect 364616 3680 364668 3732
rect 381544 3680 381596 3732
rect 520740 3748 520792 3800
rect 12348 3612 12400 3664
rect 15844 3612 15896 3664
rect 37188 3612 37240 3664
rect 68284 3612 68336 3664
rect 2872 3544 2924 3596
rect 13084 3544 13136 3596
rect 60740 3544 60792 3596
rect 61660 3544 61712 3596
rect 67916 3544 67968 3596
rect 69112 3544 69164 3596
rect 71044 3544 71096 3596
rect 77392 3612 77444 3664
rect 80704 3612 80756 3664
rect 86868 3612 86920 3664
rect 88984 3612 89036 3664
rect 109316 3612 109368 3664
rect 112444 3612 112496 3664
rect 118792 3612 118844 3664
rect 120724 3612 120776 3664
rect 121092 3612 121144 3664
rect 122104 3612 122156 3664
rect 124680 3612 124732 3664
rect 123392 3544 123444 3596
rect 126980 3544 127032 3596
rect 128176 3544 128228 3596
rect 129372 3612 129424 3664
rect 160192 3612 160244 3664
rect 170772 3612 170824 3664
rect 174636 3612 174688 3664
rect 179236 3612 179288 3664
rect 200304 3612 200356 3664
rect 215944 3612 215996 3664
rect 242900 3612 242952 3664
rect 251824 3612 251876 3664
rect 254676 3612 254728 3664
rect 254768 3612 254820 3664
rect 374000 3612 374052 3664
rect 387064 3612 387116 3664
rect 573916 3612 573968 3664
rect 162124 3544 162176 3596
rect 169576 3544 169628 3596
rect 174544 3544 174596 3596
rect 179328 3544 179380 3596
rect 184940 3544 184992 3596
rect 186228 3544 186280 3596
rect 294880 3544 294932 3596
rect 295984 3544 296036 3596
rect 299480 3544 299532 3596
rect 299572 3544 299624 3596
rect 300768 3544 300820 3596
rect 305736 3544 305788 3596
rect 307668 3544 307720 3596
rect 307852 3544 307904 3596
rect 309048 3544 309100 3596
rect 316684 3544 316736 3596
rect 321100 3544 321152 3596
rect 321468 3544 321520 3596
rect 510068 3544 510120 3596
rect 1676 3476 1728 3528
rect 14464 3476 14516 3528
rect 17040 3476 17092 3528
rect 18604 3476 18656 3528
rect 23020 3476 23072 3528
rect 24124 3476 24176 3528
rect 38384 3476 38436 3528
rect 39304 3476 39356 3528
rect 41880 3476 41932 3528
rect 43444 3476 43496 3528
rect 46664 3476 46716 3528
rect 6460 3408 6512 3460
rect 157984 3408 158036 3460
rect 160100 3476 160152 3528
rect 161296 3476 161348 3528
rect 168380 3476 168432 3528
rect 176384 3476 176436 3528
rect 182088 3476 182140 3528
rect 183744 3476 183796 3528
rect 160744 3408 160796 3460
rect 166080 3408 166132 3460
rect 173164 3408 173216 3460
rect 181536 3408 181588 3460
rect 191104 3476 191156 3528
rect 192024 3476 192076 3528
rect 193864 3476 193916 3528
rect 195612 3476 195664 3528
rect 196624 3476 196676 3528
rect 199108 3476 199160 3528
rect 199936 3476 199988 3528
rect 468300 3476 468352 3528
rect 468484 3476 468536 3528
rect 469864 3476 469916 3528
rect 472624 3476 472676 3528
rect 473452 3476 473504 3528
rect 498200 3476 498252 3528
rect 499028 3476 499080 3528
rect 520924 3476 520976 3528
rect 521844 3476 521896 3528
rect 522304 3476 522356 3528
rect 523040 3476 523092 3528
rect 564440 3476 564492 3528
rect 565268 3476 565320 3528
rect 193220 3408 193272 3460
rect 200028 3408 200080 3460
rect 472256 3408 472308 3460
rect 78588 3340 78640 3392
rect 79324 3340 79376 3392
rect 110420 3340 110472 3392
rect 111616 3340 111668 3392
rect 114008 3340 114060 3392
rect 115204 3340 115256 3392
rect 118700 3340 118752 3392
rect 119896 3340 119948 3392
rect 126980 3340 127032 3392
rect 129004 3340 129056 3392
rect 149520 3340 149572 3392
rect 151084 3340 151136 3392
rect 182824 3340 182876 3392
rect 196808 3340 196860 3392
rect 239404 3340 239456 3392
rect 253480 3340 253532 3392
rect 253572 3340 253624 3392
rect 258264 3340 258316 3392
rect 264244 3340 264296 3392
rect 271236 3340 271288 3392
rect 275284 3340 275336 3392
rect 278320 3340 278372 3392
rect 307668 3340 307720 3392
rect 315028 3340 315080 3392
rect 324412 3340 324464 3392
rect 325608 3340 325660 3392
rect 327540 3340 327592 3392
rect 335084 3340 335136 3392
rect 340972 3340 341024 3392
rect 342168 3340 342220 3392
rect 349252 3340 349304 3392
rect 350448 3340 350500 3392
rect 359464 3340 359516 3392
rect 363512 3340 363564 3392
rect 374092 3340 374144 3392
rect 375288 3340 375340 3392
rect 376116 3340 376168 3392
rect 381176 3340 381228 3392
rect 390560 3340 390612 3392
rect 391848 3340 391900 3392
rect 398932 3340 398984 3392
rect 400128 3340 400180 3392
rect 407212 3340 407264 3392
rect 408408 3340 408460 3392
rect 423772 3340 423824 3392
rect 424968 3340 425020 3392
rect 570604 3340 570656 3392
rect 577412 3340 577464 3392
rect 4068 3272 4120 3324
rect 4804 3272 4856 3324
rect 24216 3272 24268 3324
rect 25504 3272 25556 3324
rect 93952 3272 94004 3324
rect 95884 3272 95936 3324
rect 162492 3272 162544 3324
rect 166264 3272 166316 3324
rect 246304 3272 246356 3324
rect 257068 3272 257120 3324
rect 265624 3272 265676 3324
rect 266544 3272 266596 3324
rect 271144 3272 271196 3324
rect 274824 3272 274876 3324
rect 571984 3272 572036 3324
rect 572720 3272 572772 3324
rect 27712 3204 27764 3256
rect 31024 3204 31076 3256
rect 31300 3204 31352 3256
rect 36544 3204 36596 3256
rect 115204 3204 115256 3256
rect 117964 3204 118016 3256
rect 160100 3204 160152 3256
rect 161480 3204 161532 3256
rect 241244 3204 241296 3256
rect 251180 3204 251232 3256
rect 253112 3204 253164 3256
rect 249708 3136 249760 3188
rect 254768 3136 254820 3188
rect 309876 3204 309928 3256
rect 313832 3204 313884 3256
rect 260656 3136 260708 3188
rect 543004 3136 543056 3188
rect 545488 3136 545540 3188
rect 552756 3136 552808 3188
rect 556160 3136 556212 3188
rect 569224 3136 569276 3188
rect 571524 3136 571576 3188
rect 189816 3068 189868 3120
rect 190828 3068 190880 3120
rect 210424 3068 210476 3120
rect 218060 3068 218112 3120
rect 287704 3068 287756 3120
rect 290188 3068 290240 3120
rect 307116 3068 307168 3120
rect 310244 3068 310296 3120
rect 471244 3068 471296 3120
rect 474556 3068 474608 3120
rect 167184 3000 167236 3052
rect 169024 3000 169076 3052
rect 184204 3000 184256 3052
rect 186136 3000 186188 3052
rect 225604 3000 225656 3052
rect 228732 3000 228784 3052
rect 278044 3000 278096 3052
rect 281908 3000 281960 3052
rect 282184 3000 282236 3052
rect 285404 3000 285456 3052
rect 289084 3000 289136 3052
rect 296076 3000 296128 3052
rect 399484 3000 399536 3052
rect 402520 3000 402572 3052
rect 422944 3000 422996 3052
rect 423772 3000 423824 3052
rect 436744 3000 436796 3052
rect 437940 3000 437992 3052
rect 514024 3000 514076 3052
rect 515956 3000 516008 3052
rect 201408 2932 201460 2984
rect 205088 2932 205140 2984
rect 240784 2932 240836 2984
rect 247592 2932 247644 2984
rect 18236 2864 18288 2916
rect 22744 2864 22796 2916
rect 242164 2864 242216 2916
rect 244096 2864 244148 2916
rect 247684 2864 247736 2916
rect 248788 2864 248840 2916
rect 291844 2864 291896 2916
rect 293684 2864 293736 2916
rect 318156 2864 318208 2916
rect 319720 2864 319772 2916
rect 448520 2456 448572 2508
rect 449808 2456 449860 2508
rect 415400 2048 415452 2100
rect 416688 2048 416740 2100
rect 440240 2048 440292 2100
rect 441528 2048 441580 2100
<< metal2 >>
rect 8086 703520 8198 704960
rect 23492 703582 24164 703610
rect 8128 700330 8156 703520
rect 8116 700324 8168 700330
rect 8116 700266 8168 700272
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 3422 671256 3478 671265
rect 3422 671191 3478 671200
rect 3436 671090 3464 671191
rect 3424 671084 3476 671090
rect 3424 671026 3476 671032
rect 7564 671084 7616 671090
rect 7564 671026 7616 671032
rect 2778 658200 2834 658209
rect 2778 658135 2834 658144
rect 2792 657014 2820 658135
rect 2780 657008 2832 657014
rect 2780 656950 2832 656956
rect 4804 657008 4856 657014
rect 4804 656950 4856 656956
rect 3424 632120 3476 632126
rect 3422 632088 3424 632097
rect 3476 632088 3478 632097
rect 3422 632023 3478 632032
rect 3422 619168 3478 619177
rect 3422 619103 3478 619112
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3238 566944 3294 566953
rect 3238 566879 3294 566888
rect 3252 565894 3280 566879
rect 3240 565888 3292 565894
rect 3240 565830 3292 565836
rect 3330 553888 3386 553897
rect 3330 553823 3386 553832
rect 3344 553450 3372 553823
rect 3332 553444 3384 553450
rect 3332 553386 3384 553392
rect 2962 527912 3018 527921
rect 2962 527847 3018 527856
rect 2976 527202 3004 527847
rect 2964 527196 3016 527202
rect 2964 527138 3016 527144
rect 3054 501800 3110 501809
rect 3054 501735 3110 501744
rect 3068 501022 3096 501735
rect 3056 501016 3108 501022
rect 3056 500958 3108 500964
rect 3054 475688 3110 475697
rect 3054 475623 3110 475632
rect 3068 474774 3096 475623
rect 3056 474768 3108 474774
rect 3056 474710 3108 474716
rect 3054 449576 3110 449585
rect 3054 449511 3110 449520
rect 3068 448662 3096 449511
rect 3056 448656 3108 448662
rect 3056 448598 3108 448604
rect 3436 420238 3464 619103
rect 3514 606112 3570 606121
rect 3514 606047 3570 606056
rect 3528 605878 3556 606047
rect 3516 605872 3568 605878
rect 3516 605814 3568 605820
rect 3514 514856 3570 514865
rect 3514 514791 3516 514800
rect 3568 514791 3570 514800
rect 3516 514762 3568 514768
rect 3514 462632 3570 462641
rect 3514 462567 3516 462576
rect 3568 462567 3570 462576
rect 3516 462538 3568 462544
rect 3514 423600 3570 423609
rect 3514 423535 3570 423544
rect 3528 422346 3556 423535
rect 3516 422340 3568 422346
rect 3516 422282 3568 422288
rect 3424 420232 3476 420238
rect 3424 420174 3476 420180
rect 4816 414730 4844 656950
rect 7576 419490 7604 671026
rect 10324 553444 10376 553450
rect 10324 553386 10376 553392
rect 8944 462596 8996 462602
rect 8944 462538 8996 462544
rect 8956 421598 8984 462538
rect 8944 421592 8996 421598
rect 8944 421534 8996 421540
rect 7564 419484 7616 419490
rect 7564 419426 7616 419432
rect 10336 418130 10364 553386
rect 13084 514820 13136 514826
rect 13084 514762 13136 514768
rect 10324 418124 10376 418130
rect 10324 418066 10376 418072
rect 4804 414724 4856 414730
rect 4804 414666 4856 414672
rect 3422 410544 3478 410553
rect 3422 410479 3478 410488
rect 3436 407114 3464 410479
rect 3424 407108 3476 407114
rect 3424 407050 3476 407056
rect 13096 403646 13124 514762
rect 23492 407794 23520 703582
rect 24136 703474 24164 703582
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 24320 703474 24348 703520
rect 24136 703446 24348 703474
rect 40052 467158 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 104912 703582 105308 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 40040 467152 40092 467158
rect 40040 467094 40092 467100
rect 71792 411942 71820 702986
rect 89180 702434 89208 703520
rect 88352 702406 89208 702434
rect 88352 449206 88380 702406
rect 104912 465730 104940 703582
rect 105280 703474 105308 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 136652 703582 137692 703610
rect 105464 703474 105492 703520
rect 105280 703446 105492 703474
rect 104900 465724 104952 465730
rect 104900 465666 104952 465672
rect 136652 450566 136680 703582
rect 137664 703474 137692 703582
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 234632 703582 235028 703610
rect 137848 703474 137876 703520
rect 137664 703446 137876 703474
rect 154132 702434 154160 703520
rect 170324 702434 170352 703520
rect 202800 703050 202828 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 153212 702406 154160 702434
rect 169772 702406 170352 702434
rect 142804 605872 142856 605878
rect 142804 605814 142856 605820
rect 136640 450560 136692 450566
rect 136640 450502 136692 450508
rect 88340 449200 88392 449206
rect 88340 449142 88392 449148
rect 142816 416090 142844 605814
rect 142804 416084 142856 416090
rect 142804 416026 142856 416032
rect 71780 411936 71832 411942
rect 71780 411878 71832 411884
rect 23480 407788 23532 407794
rect 23480 407730 23532 407736
rect 13084 403640 13136 403646
rect 13084 403582 13136 403588
rect 3424 397520 3476 397526
rect 3422 397488 3424 397497
rect 3476 397488 3478 397497
rect 3422 397423 3478 397432
rect 153212 373998 153240 702406
rect 169772 464370 169800 702406
rect 195244 565888 195296 565894
rect 195244 565830 195296 565836
rect 169760 464364 169812 464370
rect 169760 464306 169812 464312
rect 195256 405006 195284 565830
rect 195244 405000 195296 405006
rect 195244 404942 195296 404948
rect 153200 373992 153252 373998
rect 153200 373934 153252 373940
rect 3422 371376 3478 371385
rect 3422 371311 3478 371320
rect 3436 371278 3464 371311
rect 3424 371272 3476 371278
rect 3424 371214 3476 371220
rect 201512 367810 201540 702986
rect 218992 699718 219020 703520
rect 218980 699712 219032 699718
rect 218980 699654 219032 699660
rect 220084 699712 220136 699718
rect 220084 699654 220136 699660
rect 219256 374672 219308 374678
rect 219256 374614 219308 374620
rect 201500 367804 201552 367810
rect 201500 367746 201552 367752
rect 3146 358456 3202 358465
rect 3146 358391 3202 358400
rect 3160 357474 3188 358391
rect 3148 357468 3200 357474
rect 3148 357410 3200 357416
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3344 345098 3372 345335
rect 3332 345092 3384 345098
rect 3332 345034 3384 345040
rect 218704 321768 218756 321774
rect 218704 321710 218756 321716
rect 206744 321700 206796 321706
rect 206744 321642 206796 321648
rect 201408 321632 201460 321638
rect 201408 321574 201460 321580
rect 202786 321600 202842 321609
rect 3422 319288 3478 319297
rect 3422 319223 3478 319232
rect 3436 318850 3464 319223
rect 3424 318844 3476 318850
rect 3424 318786 3476 318792
rect 197360 318844 197412 318850
rect 197360 318786 197412 318792
rect 4066 306232 4122 306241
rect 4122 306190 4200 306218
rect 4066 306167 4122 306176
rect 4172 299470 4200 306190
rect 193220 300144 193272 300150
rect 193220 300086 193272 300092
rect 4160 299464 4212 299470
rect 4160 299406 4212 299412
rect 178684 297288 178736 297294
rect 178684 297230 178736 297236
rect 176660 297084 176712 297090
rect 176660 297026 176712 297032
rect 173900 296948 173952 296954
rect 173900 296890 173952 296896
rect 169760 296064 169812 296070
rect 169760 296006 169812 296012
rect 167000 294840 167052 294846
rect 167000 294782 167052 294788
rect 164240 294636 164292 294642
rect 164240 294578 164292 294584
rect 157800 293276 157852 293282
rect 157800 293218 157852 293224
rect 3422 293176 3478 293185
rect 3422 293111 3478 293120
rect 3436 292602 3464 293111
rect 3424 292596 3476 292602
rect 3424 292538 3476 292544
rect 3054 267200 3110 267209
rect 3054 267135 3110 267144
rect 3068 266422 3096 267135
rect 3056 266416 3108 266422
rect 3056 266358 3108 266364
rect 14464 266416 14516 266422
rect 14464 266358 14516 266364
rect 3422 254144 3478 254153
rect 3422 254079 3478 254088
rect 3436 253978 3464 254079
rect 3424 253972 3476 253978
rect 3424 253914 3476 253920
rect 3330 241088 3386 241097
rect 3330 241023 3386 241032
rect 3344 239426 3372 241023
rect 14476 240786 14504 266358
rect 154396 242208 154448 242214
rect 154396 242150 154448 242156
rect 153014 241904 153070 241913
rect 153014 241839 153070 241848
rect 151726 241768 151782 241777
rect 151726 241703 151782 241712
rect 151634 241632 151690 241641
rect 151634 241567 151690 241576
rect 14464 240780 14516 240786
rect 14464 240722 14516 240728
rect 3332 239420 3384 239426
rect 3332 239362 3384 239368
rect 151544 238808 151596 238814
rect 151544 238750 151596 238756
rect 150346 229800 150402 229809
rect 150346 229735 150402 229744
rect 3422 214976 3478 214985
rect 3422 214911 3478 214920
rect 3436 214606 3464 214911
rect 3424 214600 3476 214606
rect 3424 214542 3476 214548
rect 28264 211812 28316 211818
rect 28264 211754 28316 211760
rect 3516 210588 3568 210594
rect 3516 210530 3568 210536
rect 3424 210520 3476 210526
rect 3424 210462 3476 210468
rect 3332 202836 3384 202842
rect 3332 202778 3384 202784
rect 3344 201929 3372 202778
rect 3330 201920 3386 201929
rect 3330 201855 3386 201864
rect 3148 189032 3200 189038
rect 3148 188974 3200 188980
rect 3160 188873 3188 188974
rect 3146 188864 3202 188873
rect 3146 188799 3202 188808
rect 3332 164212 3384 164218
rect 3332 164154 3384 164160
rect 3344 162897 3372 164154
rect 3330 162888 3386 162897
rect 3330 162823 3386 162832
rect 3148 111784 3200 111790
rect 3148 111726 3200 111732
rect 3160 110673 3188 111726
rect 3146 110664 3202 110673
rect 3146 110599 3202 110608
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 2872 33108 2924 33114
rect 2872 33050 2924 33056
rect 2884 32473 2912 33050
rect 2870 32464 2926 32473
rect 2870 32399 2926 32408
rect 3436 19417 3464 210462
rect 3528 97617 3556 210530
rect 3608 210452 3660 210458
rect 3608 210394 3660 210400
rect 3620 136785 3648 210394
rect 11704 208412 11756 208418
rect 11704 208354 11756 208360
rect 3700 159384 3752 159390
rect 3700 159326 3752 159332
rect 3712 149841 3740 159326
rect 6920 155236 6972 155242
rect 6920 155178 6972 155184
rect 3698 149832 3754 149841
rect 3698 149767 3754 149776
rect 3606 136776 3662 136785
rect 3606 136711 3662 136720
rect 4804 135924 4856 135930
rect 4804 135866 4856 135872
rect 3514 97608 3570 97617
rect 3514 97543 3570 97552
rect 3516 85536 3568 85542
rect 3516 85478 3568 85484
rect 3528 84697 3556 85478
rect 3514 84688 3570 84697
rect 3514 84623 3570 84632
rect 3516 71732 3568 71738
rect 3516 71674 3568 71680
rect 3528 71641 3556 71674
rect 3514 71632 3570 71641
rect 3514 71567 3570 71576
rect 3516 45552 3568 45558
rect 3514 45520 3516 45529
rect 3568 45520 3570 45529
rect 3514 45455 3570 45464
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 2872 3596 2924 3602
rect 2872 3538 2924 3544
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 1688 480 1716 3470
rect 2884 480 2912 3538
rect 4816 3330 4844 135866
rect 6932 16574 6960 155178
rect 8300 134564 8352 134570
rect 8300 134506 8352 134512
rect 8312 16574 8340 134506
rect 9680 112464 9732 112470
rect 9680 112406 9732 112412
rect 6932 16546 7696 16574
rect 8312 16546 8800 16574
rect 5264 4820 5316 4826
rect 5264 4762 5316 4768
rect 4068 3324 4120 3330
rect 4068 3266 4120 3272
rect 4804 3324 4856 3330
rect 4804 3266 4856 3272
rect 4080 480 4108 3266
rect 5276 480 5304 4762
rect 6460 3460 6512 3466
rect 6460 3402 6512 3408
rect 6472 480 6500 3402
rect 7668 480 7696 16546
rect 8772 480 8800 16546
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 112406
rect 11060 93152 11112 93158
rect 11060 93094 11112 93100
rect 11072 16574 11100 93094
rect 11716 33114 11744 208354
rect 25504 155304 25556 155310
rect 25504 155246 25556 155252
rect 15844 148368 15896 148374
rect 15844 148310 15896 148316
rect 14464 146940 14516 146946
rect 14464 146882 14516 146888
rect 13084 144220 13136 144226
rect 13084 144162 13136 144168
rect 11704 33108 11756 33114
rect 11704 33050 11756 33056
rect 11072 16546 11192 16574
rect 11164 480 11192 16546
rect 12348 3664 12400 3670
rect 12348 3606 12400 3612
rect 12360 480 12388 3606
rect 13096 3602 13124 144162
rect 13820 105596 13872 105602
rect 13820 105538 13872 105544
rect 13832 16574 13860 105538
rect 13832 16546 14320 16574
rect 13544 4072 13596 4078
rect 13544 4014 13596 4020
rect 13084 3596 13136 3602
rect 13084 3538 13136 3544
rect 13556 480 13584 4014
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 14476 3534 14504 146882
rect 15752 11756 15804 11762
rect 15752 11698 15804 11704
rect 14464 3528 14516 3534
rect 14464 3470 14516 3476
rect 15764 3482 15792 11698
rect 15856 3670 15884 148310
rect 18602 145616 18658 145625
rect 18602 145551 18658 145560
rect 17224 140072 17276 140078
rect 17224 140014 17276 140020
rect 17236 4078 17264 140014
rect 17224 4072 17276 4078
rect 17224 4014 17276 4020
rect 15844 3664 15896 3670
rect 15844 3606 15896 3612
rect 18616 3534 18644 145551
rect 20718 122088 20774 122097
rect 20718 122023 20774 122032
rect 19340 100020 19392 100026
rect 19340 99962 19392 99968
rect 19352 16574 19380 99962
rect 20732 16574 20760 122023
rect 22744 119400 22796 119406
rect 22744 119342 22796 119348
rect 19352 16546 19472 16574
rect 20732 16546 21864 16574
rect 17040 3528 17092 3534
rect 15764 3454 15976 3482
rect 17040 3470 17092 3476
rect 18604 3528 18656 3534
rect 18604 3470 18656 3476
rect 15948 480 15976 3454
rect 17052 480 17080 3470
rect 18236 2916 18288 2922
rect 18236 2858 18288 2864
rect 18248 480 18276 2858
rect 19444 480 19472 16546
rect 20168 10328 20220 10334
rect 20168 10270 20220 10276
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20180 354 20208 10270
rect 21836 480 21864 16546
rect 22756 2922 22784 119342
rect 24124 117972 24176 117978
rect 24124 117914 24176 117920
rect 24136 3534 24164 117914
rect 25320 13116 25372 13122
rect 25320 13058 25372 13064
rect 23020 3528 23072 3534
rect 23020 3470 23072 3476
rect 24124 3528 24176 3534
rect 24124 3470 24176 3476
rect 22744 2916 22796 2922
rect 22744 2858 22796 2864
rect 23032 480 23060 3470
rect 24216 3324 24268 3330
rect 24216 3266 24268 3272
rect 24228 480 24256 3266
rect 25332 480 25360 13058
rect 25516 3330 25544 155246
rect 26240 137284 26292 137290
rect 26240 137226 26292 137232
rect 25504 3324 25556 3330
rect 25504 3266 25556 3272
rect 20598 354 20710 480
rect 20180 326 20710 354
rect 20598 -960 20710 326
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 137226
rect 27620 97300 27672 97306
rect 27620 97242 27672 97248
rect 27632 16574 27660 97242
rect 28276 85542 28304 211754
rect 146944 209160 146996 209166
rect 146944 209102 146996 209108
rect 120816 209092 120868 209098
rect 120816 209034 120868 209040
rect 96620 159520 96672 159526
rect 96620 159462 96672 159468
rect 78680 159452 78732 159458
rect 78680 159394 78732 159400
rect 60740 158092 60792 158098
rect 60740 158034 60792 158040
rect 46204 158024 46256 158030
rect 46204 157966 46256 157972
rect 28998 153776 29054 153785
rect 28998 153711 29054 153720
rect 28264 85536 28316 85542
rect 28264 85478 28316 85484
rect 29012 16574 29040 153711
rect 34518 151056 34574 151065
rect 34518 150991 34574 151000
rect 33140 142860 33192 142866
rect 33140 142802 33192 142808
rect 31024 141432 31076 141438
rect 31024 141374 31076 141380
rect 27632 16546 28488 16574
rect 29012 16546 30144 16574
rect 27712 3256 27764 3262
rect 27712 3198 27764 3204
rect 27724 480 27752 3198
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28460 354 28488 16546
rect 30116 480 30144 16546
rect 31036 3262 31064 141374
rect 31760 102808 31812 102814
rect 31760 102750 31812 102756
rect 31772 16574 31800 102750
rect 33152 16574 33180 142802
rect 31772 16546 31984 16574
rect 33152 16546 33640 16574
rect 31024 3256 31076 3262
rect 31024 3198 31076 3204
rect 31300 3256 31352 3262
rect 31300 3198 31352 3204
rect 31312 480 31340 3198
rect 28878 354 28990 480
rect 28460 326 28990 354
rect 28878 -960 28990 326
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 31956 354 31984 16546
rect 33612 480 33640 16546
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34532 354 34560 150991
rect 44180 141500 44232 141506
rect 44180 141442 44232 141448
rect 40040 140140 40092 140146
rect 40040 140082 40092 140088
rect 36542 130384 36598 130393
rect 36542 130319 36598 130328
rect 35900 94512 35952 94518
rect 35900 94454 35952 94460
rect 35912 16574 35940 94454
rect 35912 16546 36032 16574
rect 36004 480 36032 16546
rect 36556 3262 36584 130319
rect 39304 116612 39356 116618
rect 39304 116554 39356 116560
rect 38660 17264 38712 17270
rect 38660 17206 38712 17212
rect 38672 16574 38700 17206
rect 38672 16546 39160 16574
rect 37188 3664 37240 3670
rect 37188 3606 37240 3612
rect 36544 3256 36596 3262
rect 36544 3198 36596 3204
rect 37200 480 37228 3606
rect 38384 3528 38436 3534
rect 38384 3470 38436 3476
rect 38396 480 38424 3470
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39132 354 39160 16546
rect 39316 3534 39344 116554
rect 40052 16574 40080 140082
rect 43444 115252 43496 115258
rect 43444 115194 43496 115200
rect 42800 77988 42852 77994
rect 42800 77930 42852 77936
rect 40052 16546 40264 16574
rect 39304 3528 39356 3534
rect 39304 3470 39356 3476
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 40236 354 40264 16546
rect 41880 3528 41932 3534
rect 41880 3470 41932 3476
rect 41892 480 41920 3470
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 39550 -960 39662 326
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 42812 354 42840 77930
rect 43456 3534 43484 115194
rect 44192 6914 44220 141442
rect 44270 113792 44326 113801
rect 44270 113727 44326 113736
rect 44284 16574 44312 113727
rect 44284 16546 45048 16574
rect 44192 6886 44312 6914
rect 43444 3528 43496 3534
rect 43444 3470 43496 3476
rect 44284 480 44312 6886
rect 43046 354 43158 480
rect 42812 326 43158 354
rect 43046 -960 43158 326
rect 44242 -960 44354 480
rect 45020 354 45048 16546
rect 46216 4826 46244 157966
rect 57980 153876 58032 153882
rect 57980 153818 58032 153824
rect 46940 152516 46992 152522
rect 46940 152458 46992 152464
rect 46952 16574 46980 152458
rect 51078 151192 51134 151201
rect 51078 151127 51134 151136
rect 49700 142928 49752 142934
rect 49700 142870 49752 142876
rect 48320 133204 48372 133210
rect 48320 133146 48372 133152
rect 48332 16574 48360 133146
rect 49712 16574 49740 142870
rect 46952 16546 47440 16574
rect 48332 16546 48544 16574
rect 49712 16546 50200 16574
rect 46204 4820 46256 4826
rect 46204 4762 46256 4768
rect 46664 3528 46716 3534
rect 46664 3470 46716 3476
rect 46676 480 46704 3470
rect 45438 354 45550 480
rect 45020 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 48516 354 48544 16546
rect 50172 480 50200 16546
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 47830 -960 47942 326
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51092 354 51120 151127
rect 53838 149696 53894 149705
rect 53838 149631 53894 149640
rect 52460 138712 52512 138718
rect 52460 138654 52512 138660
rect 52472 6914 52500 138654
rect 52552 109744 52604 109750
rect 52552 109686 52604 109692
rect 52564 16574 52592 109686
rect 53852 16574 53880 149631
rect 55218 131744 55274 131753
rect 55218 131679 55274 131688
rect 55232 16574 55260 131679
rect 56600 124908 56652 124914
rect 56600 124850 56652 124856
rect 56612 16574 56640 124850
rect 57992 16574 58020 153818
rect 59358 137320 59414 137329
rect 59358 137255 59414 137264
rect 52564 16546 53328 16574
rect 53852 16546 54984 16574
rect 55232 16546 56088 16574
rect 56612 16546 56824 16574
rect 57992 16546 58480 16574
rect 52472 6886 52592 6914
rect 52564 480 52592 6886
rect 51326 354 51438 480
rect 51092 326 51438 354
rect 51326 -960 51438 326
rect 52522 -960 52634 480
rect 53300 354 53328 16546
rect 54956 480 54984 16546
rect 56060 480 56088 16546
rect 53718 354 53830 480
rect 53300 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 16546
rect 58452 480 58480 16546
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59372 354 59400 137255
rect 60752 3602 60780 158034
rect 74540 156664 74592 156670
rect 74540 156606 74592 156612
rect 71042 153912 71098 153921
rect 71042 153847 71098 153856
rect 64878 151328 64934 151337
rect 64878 151263 64934 151272
rect 62120 138780 62172 138786
rect 62120 138722 62172 138728
rect 60832 120760 60884 120766
rect 60832 120702 60884 120708
rect 60740 3596 60792 3602
rect 60740 3538 60792 3544
rect 60844 480 60872 120702
rect 62132 16574 62160 138722
rect 64892 16574 64920 151263
rect 68284 147008 68336 147014
rect 68284 146950 68336 146956
rect 66260 129056 66312 129062
rect 66260 128998 66312 129004
rect 66272 16574 66300 128998
rect 62132 16546 63264 16574
rect 64892 16546 65104 16574
rect 66272 16546 66760 16574
rect 61660 3596 61712 3602
rect 61660 3538 61712 3544
rect 59606 354 59718 480
rect 59372 326 59718 354
rect 59606 -960 59718 326
rect 60802 -960 60914 480
rect 61672 354 61700 3538
rect 63236 480 63264 16546
rect 64328 4820 64380 4826
rect 64328 4762 64380 4768
rect 64340 480 64368 4762
rect 61998 354 62110 480
rect 61672 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65076 354 65104 16546
rect 66732 480 66760 16546
rect 68296 3670 68324 146950
rect 69020 127628 69072 127634
rect 69020 127570 69072 127576
rect 69032 16574 69060 127570
rect 70400 108316 70452 108322
rect 70400 108258 70452 108264
rect 70412 16574 70440 108258
rect 69032 16546 69888 16574
rect 70412 16546 70992 16574
rect 68284 3664 68336 3670
rect 68284 3606 68336 3612
rect 67916 3596 67968 3602
rect 67916 3538 67968 3544
rect 69112 3596 69164 3602
rect 69112 3538 69164 3544
rect 67928 480 67956 3538
rect 69124 480 69152 3538
rect 65494 354 65606 480
rect 65076 326 65606 354
rect 65494 -960 65606 326
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 69860 354 69888 16546
rect 70964 3482 70992 16546
rect 71056 3602 71084 153847
rect 71780 149728 71832 149734
rect 71780 149670 71832 149676
rect 71792 16574 71820 149670
rect 74552 16574 74580 156606
rect 75918 148336 75974 148345
rect 75918 148271 75974 148280
rect 71792 16546 72648 16574
rect 74552 16546 75040 16574
rect 71044 3596 71096 3602
rect 71044 3538 71096 3544
rect 70964 3454 71544 3482
rect 71516 480 71544 3454
rect 72620 480 72648 16546
rect 73804 7608 73856 7614
rect 73804 7550 73856 7556
rect 73816 480 73844 7550
rect 75012 480 75040 16546
rect 70278 354 70390 480
rect 69860 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 75932 354 75960 148271
rect 78692 16574 78720 159394
rect 85580 156800 85632 156806
rect 85580 156742 85632 156748
rect 81440 156732 81492 156738
rect 81440 156674 81492 156680
rect 80702 135960 80758 135969
rect 80702 135895 80758 135904
rect 80058 126304 80114 126313
rect 80058 126239 80114 126248
rect 79324 106956 79376 106962
rect 79324 106898 79376 106904
rect 78692 16546 79272 16574
rect 77392 3664 77444 3670
rect 77392 3606 77444 3612
rect 77404 480 77432 3606
rect 78588 3392 78640 3398
rect 78588 3334 78640 3340
rect 78600 480 78628 3334
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79244 354 79272 16546
rect 79336 3398 79364 106898
rect 80072 16574 80100 126239
rect 80072 16546 80652 16574
rect 80624 3482 80652 16546
rect 80716 3670 80744 135895
rect 81452 16574 81480 156674
rect 82820 148436 82872 148442
rect 82820 148378 82872 148384
rect 82832 16574 82860 148378
rect 84198 130520 84254 130529
rect 84198 130455 84254 130464
rect 81452 16546 81664 16574
rect 82832 16546 83320 16574
rect 80704 3664 80756 3670
rect 80704 3606 80756 3612
rect 80624 3454 80928 3482
rect 79324 3392 79376 3398
rect 79324 3334 79376 3340
rect 80900 480 80928 3454
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 83292 480 83320 16546
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84212 354 84240 130455
rect 85592 16574 85620 156742
rect 92480 153944 92532 153950
rect 92480 153886 92532 153892
rect 89718 152416 89774 152425
rect 89718 152351 89774 152360
rect 88984 145580 89036 145586
rect 88984 145522 89036 145528
rect 86960 123480 87012 123486
rect 86960 123422 87012 123428
rect 86972 16574 87000 123422
rect 85592 16546 85712 16574
rect 86972 16546 87552 16574
rect 85684 480 85712 16546
rect 86868 3664 86920 3670
rect 86868 3606 86920 3612
rect 86880 480 86908 3606
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87524 354 87552 16546
rect 88892 14476 88944 14482
rect 88892 14418 88944 14424
rect 88904 3482 88932 14418
rect 88996 3670 89024 145522
rect 89732 16574 89760 152351
rect 91100 134632 91152 134638
rect 91100 134574 91152 134580
rect 91112 16574 91140 134574
rect 89732 16546 89944 16574
rect 91112 16546 91600 16574
rect 88984 3664 89036 3670
rect 88984 3606 89036 3612
rect 88904 3454 89208 3482
rect 89180 480 89208 3454
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91572 480 91600 16546
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 153886
rect 95884 145648 95936 145654
rect 95884 145590 95936 145596
rect 93860 144288 93912 144294
rect 93860 144230 93912 144236
rect 93872 16574 93900 144230
rect 95240 104168 95292 104174
rect 95240 104110 95292 104116
rect 95252 16574 95280 104110
rect 93872 16546 94728 16574
rect 95252 16546 95832 16574
rect 93952 3324 94004 3330
rect 93952 3266 94004 3272
rect 93964 480 93992 3266
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 94700 354 94728 16546
rect 95118 354 95230 480
rect 94700 326 95230 354
rect 95804 354 95832 16546
rect 95896 3330 95924 145590
rect 96632 16574 96660 159462
rect 106280 156936 106332 156942
rect 106280 156878 106332 156884
rect 99380 156868 99432 156874
rect 99380 156810 99432 156816
rect 98000 133272 98052 133278
rect 98000 133214 98052 133220
rect 98012 16574 98040 133214
rect 99392 16574 99420 156810
rect 100758 155272 100814 155281
rect 100758 155207 100814 155216
rect 96632 16546 97488 16574
rect 98012 16546 98224 16574
rect 99392 16546 99880 16574
rect 95884 3324 95936 3330
rect 95884 3266 95936 3272
rect 97460 480 97488 16546
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 95118 -960 95230 326
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98196 354 98224 16546
rect 99852 480 99880 16546
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 100772 354 100800 155207
rect 104900 152584 104952 152590
rect 104900 152526 104952 152532
rect 103518 146976 103574 146985
rect 103518 146911 103574 146920
rect 102140 124976 102192 124982
rect 102140 124918 102192 124924
rect 102152 16574 102180 124918
rect 103532 16574 103560 146911
rect 104912 16574 104940 152526
rect 106292 16574 106320 156878
rect 110418 149832 110474 149841
rect 110418 149767 110474 149776
rect 107660 142996 107712 143002
rect 107660 142938 107712 142944
rect 107672 16574 107700 142938
rect 102152 16546 102272 16574
rect 103532 16546 104112 16574
rect 104912 16546 105768 16574
rect 106292 16546 106504 16574
rect 107672 16546 108160 16574
rect 102244 480 102272 16546
rect 103336 8968 103388 8974
rect 103336 8910 103388 8916
rect 103348 480 103376 8910
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 16546
rect 105740 480 105768 16546
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 108132 480 108160 16546
rect 109316 3664 109368 3670
rect 109316 3606 109368 3612
rect 109328 480 109356 3606
rect 110432 3398 110460 149767
rect 120722 147112 120778 147121
rect 120722 147047 120778 147056
rect 118700 145716 118752 145722
rect 118700 145658 118752 145664
rect 117962 144120 118018 144129
rect 117962 144055 118018 144064
rect 115204 140208 115256 140214
rect 115204 140150 115256 140156
rect 110512 131776 110564 131782
rect 110512 131718 110564 131724
rect 110420 3392 110472 3398
rect 110420 3334 110472 3340
rect 110524 480 110552 131718
rect 112442 122224 112498 122233
rect 112442 122159 112498 122168
rect 111800 98660 111852 98666
rect 111800 98602 111852 98608
rect 111812 16574 111840 98602
rect 111812 16546 112392 16574
rect 111616 3392 111668 3398
rect 111616 3334 111668 3340
rect 111628 480 111656 3334
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 16546
rect 112456 3670 112484 122159
rect 112444 3664 112496 3670
rect 112444 3606 112496 3612
rect 115216 3398 115244 140150
rect 115940 138848 115992 138854
rect 115940 138790 115992 138796
rect 115952 16574 115980 138790
rect 117320 129124 117372 129130
rect 117320 129066 117372 129072
rect 115952 16546 116440 16574
rect 114008 3392 114060 3398
rect 114008 3334 114060 3340
rect 115204 3392 115256 3398
rect 115204 3334 115256 3340
rect 114020 480 114048 3334
rect 115204 3256 115256 3262
rect 115204 3198 115256 3204
rect 115216 480 115244 3198
rect 116412 480 116440 16546
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117332 354 117360 129066
rect 117976 3262 118004 144055
rect 118712 3398 118740 145658
rect 120736 3670 120764 147047
rect 120828 111790 120856 209034
rect 132500 159792 132552 159798
rect 132500 159734 132552 159740
rect 125600 159588 125652 159594
rect 125600 159530 125652 159536
rect 124864 158160 124916 158166
rect 124864 158102 124916 158108
rect 123484 157004 123536 157010
rect 123484 156946 123536 156952
rect 121460 141568 121512 141574
rect 121460 141510 121512 141516
rect 120816 111784 120868 111790
rect 120816 111726 120868 111732
rect 121472 16574 121500 141510
rect 122104 127696 122156 127702
rect 122104 127638 122156 127644
rect 121472 16546 122052 16574
rect 118792 3664 118844 3670
rect 118792 3606 118844 3612
rect 120724 3664 120776 3670
rect 120724 3606 120776 3612
rect 121092 3664 121144 3670
rect 121092 3606 121144 3612
rect 118700 3392 118752 3398
rect 118700 3334 118752 3340
rect 117964 3256 118016 3262
rect 117964 3198 118016 3204
rect 118804 480 118832 3606
rect 119896 3392 119948 3398
rect 119896 3334 119948 3340
rect 119908 480 119936 3334
rect 121104 480 121132 3606
rect 122024 3482 122052 16546
rect 122116 3670 122144 127638
rect 123496 6914 123524 156946
rect 124876 10334 124904 158102
rect 124864 10328 124916 10334
rect 124864 10270 124916 10276
rect 123404 6886 123524 6914
rect 122104 3664 122156 3670
rect 122104 3606 122156 3612
rect 123404 3602 123432 6886
rect 123484 3732 123536 3738
rect 123484 3674 123536 3680
rect 123392 3596 123444 3602
rect 123392 3538 123444 3544
rect 122024 3454 122328 3482
rect 122300 480 122328 3454
rect 123496 480 123524 3674
rect 124680 3664 124732 3670
rect 124680 3606 124732 3612
rect 124692 480 124720 3606
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125612 354 125640 159530
rect 126978 154048 127034 154057
rect 126978 153983 127034 153992
rect 126992 3602 127020 153983
rect 129002 136096 129058 136105
rect 129002 136031 129058 136040
rect 126980 3596 127032 3602
rect 126980 3538 127032 3544
rect 128176 3596 128228 3602
rect 128176 3538 128228 3544
rect 126980 3392 127032 3398
rect 126980 3334 127032 3340
rect 126992 480 127020 3334
rect 128188 480 128216 3538
rect 129016 3398 129044 136031
rect 129738 126440 129794 126449
rect 129738 126375 129794 126384
rect 129752 16574 129780 126375
rect 131120 111104 131172 111110
rect 131120 111046 131172 111052
rect 131132 16574 131160 111046
rect 132512 16574 132540 159734
rect 135260 159724 135312 159730
rect 135260 159666 135312 159672
rect 133880 152652 133932 152658
rect 133880 152594 133932 152600
rect 133144 148504 133196 148510
rect 133144 148446 133196 148452
rect 129752 16546 130608 16574
rect 131132 16546 131344 16574
rect 132512 16546 133000 16574
rect 129372 3664 129424 3670
rect 129372 3606 129424 3612
rect 129004 3392 129056 3398
rect 129004 3334 129056 3340
rect 129384 480 129412 3606
rect 130580 480 130608 16546
rect 125846 354 125958 480
rect 125612 326 125958 354
rect 125846 -960 125958 326
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131316 354 131344 16546
rect 132972 480 133000 16546
rect 133156 3738 133184 148446
rect 133144 3732 133196 3738
rect 133144 3674 133196 3680
rect 131734 354 131846 480
rect 131316 326 131846 354
rect 131734 -960 131846 326
rect 132930 -960 133042 480
rect 133892 354 133920 152594
rect 135272 3738 135300 159666
rect 139400 159656 139452 159662
rect 139400 159598 139452 159604
rect 138020 154012 138072 154018
rect 138020 153954 138072 153960
rect 135350 149968 135406 149977
rect 135350 149903 135406 149912
rect 135260 3732 135312 3738
rect 135260 3674 135312 3680
rect 135364 3482 135392 149903
rect 136638 148472 136694 148481
rect 136638 148407 136694 148416
rect 136652 16574 136680 148407
rect 138032 16574 138060 153954
rect 139412 16574 139440 159598
rect 144920 155372 144972 155378
rect 144920 155314 144972 155320
rect 142160 151088 142212 151094
rect 142160 151030 142212 151036
rect 140778 140040 140834 140049
rect 140778 139975 140834 139984
rect 140792 16574 140820 139975
rect 136652 16546 137232 16574
rect 138032 16546 138888 16574
rect 139412 16546 139624 16574
rect 140792 16546 141280 16574
rect 136456 3732 136508 3738
rect 136456 3674 136508 3680
rect 135272 3454 135392 3482
rect 135272 480 135300 3454
rect 136468 480 136496 3674
rect 134126 354 134238 480
rect 133892 326 134238 354
rect 134126 -960 134238 326
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137204 354 137232 16546
rect 138860 480 138888 16546
rect 137622 354 137734 480
rect 137204 326 137734 354
rect 137622 -960 137734 326
rect 138818 -960 138930 480
rect 139596 354 139624 16546
rect 141252 480 141280 16546
rect 140014 354 140126 480
rect 139596 326 140126 354
rect 140014 -960 140126 326
rect 141210 -960 141322 480
rect 142172 354 142200 151030
rect 143540 147076 143592 147082
rect 143540 147018 143592 147024
rect 143552 11830 143580 147018
rect 143632 143064 143684 143070
rect 143632 143006 143684 143012
rect 143540 11824 143592 11830
rect 143540 11766 143592 11772
rect 143644 6914 143672 143006
rect 144932 16574 144960 155314
rect 146300 137352 146352 137358
rect 146300 137294 146352 137300
rect 146312 16574 146340 137294
rect 146956 71738 146984 209102
rect 148324 158296 148376 158302
rect 148324 158238 148376 158244
rect 147678 141400 147734 141409
rect 147678 141335 147734 141344
rect 146944 71732 146996 71738
rect 146944 71674 146996 71680
rect 147692 16574 147720 141335
rect 148336 93158 148364 158238
rect 150360 155922 150388 229735
rect 150440 159860 150492 159866
rect 150440 159802 150492 159808
rect 149704 155916 149756 155922
rect 149704 155858 149756 155864
rect 150348 155916 150400 155922
rect 150348 155858 150400 155864
rect 149716 151065 149744 155858
rect 149702 151056 149758 151065
rect 149702 150991 149758 151000
rect 148324 93152 148376 93158
rect 148324 93094 148376 93100
rect 150452 16574 150480 159802
rect 151556 158953 151584 238750
rect 151266 158944 151322 158953
rect 151266 158879 151322 158888
rect 151542 158944 151598 158953
rect 151542 158879 151598 158888
rect 151176 158432 151228 158438
rect 151176 158374 151228 158380
rect 151084 151156 151136 151162
rect 151084 151098 151136 151104
rect 144932 16546 145512 16574
rect 146312 16546 147168 16574
rect 147692 16546 147904 16574
rect 150452 16546 150664 16574
rect 144736 11824 144788 11830
rect 144736 11766 144788 11772
rect 143552 6886 143672 6914
rect 143552 480 143580 6886
rect 144748 480 144776 11766
rect 142406 354 142518 480
rect 142172 326 142518 354
rect 142406 -960 142518 326
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145484 354 145512 16546
rect 147140 480 147168 16546
rect 145902 354 146014 480
rect 145484 326 146014 354
rect 145902 -960 146014 326
rect 147098 -960 147210 480
rect 147876 354 147904 16546
rect 149520 3392 149572 3398
rect 149520 3334 149572 3340
rect 149532 480 149560 3334
rect 150636 480 150664 16546
rect 151096 3398 151124 151098
rect 151188 77994 151216 158374
rect 151280 147014 151308 158879
rect 151648 158438 151676 241567
rect 151636 158432 151688 158438
rect 151636 158374 151688 158380
rect 151740 156466 151768 241703
rect 152922 240816 152978 240825
rect 152922 240751 152978 240760
rect 152832 232620 152884 232626
rect 152832 232562 152884 232568
rect 152740 231260 152792 231266
rect 152740 231202 152792 231208
rect 152648 218816 152700 218822
rect 152648 218758 152700 218764
rect 152554 159624 152610 159633
rect 152554 159559 152610 159568
rect 151728 156460 151780 156466
rect 151728 156402 151780 156408
rect 152568 152425 152596 159559
rect 152660 159458 152688 218758
rect 152648 159452 152700 159458
rect 152648 159394 152700 159400
rect 152752 159050 152780 231202
rect 152740 159044 152792 159050
rect 152740 158986 152792 158992
rect 152844 156777 152872 232562
rect 152936 159633 152964 240751
rect 152922 159624 152978 159633
rect 152922 159559 152978 159568
rect 152924 159452 152976 159458
rect 152924 159394 152976 159400
rect 152936 158982 152964 159394
rect 153028 159118 153056 241839
rect 153108 240848 153160 240854
rect 153108 240790 153160 240796
rect 153016 159112 153068 159118
rect 153016 159054 153068 159060
rect 152924 158976 152976 158982
rect 152924 158918 152976 158924
rect 152830 156768 152886 156777
rect 152830 156703 152886 156712
rect 152554 152416 152610 152425
rect 152554 152351 152610 152360
rect 151820 149116 151872 149122
rect 151820 149058 151872 149064
rect 151268 147008 151320 147014
rect 151268 146950 151320 146956
rect 151176 77988 151228 77994
rect 151176 77930 151228 77936
rect 151084 3392 151136 3398
rect 151084 3334 151136 3340
rect 151832 480 151860 149058
rect 151912 148572 151964 148578
rect 151912 148514 151964 148520
rect 151924 16574 151952 148514
rect 152844 148442 152872 156703
rect 152832 148436 152884 148442
rect 152832 148378 152884 148384
rect 153120 147529 153148 240790
rect 154304 238944 154356 238950
rect 154304 238886 154356 238892
rect 154212 225684 154264 225690
rect 154212 225626 154264 225632
rect 154118 220144 154174 220153
rect 154118 220079 154174 220088
rect 153844 209840 153896 209846
rect 153844 209782 153896 209788
rect 153200 155440 153252 155446
rect 153200 155382 153252 155388
rect 153106 147520 153162 147529
rect 153106 147455 153162 147464
rect 153212 16574 153240 155382
rect 151924 16546 153056 16574
rect 153212 16546 153792 16574
rect 153028 480 153056 16546
rect 148294 354 148406 480
rect 147876 326 148406 354
rect 148294 -960 148406 326
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 153764 354 153792 16546
rect 153856 6866 153884 209782
rect 153936 158364 153988 158370
rect 153936 158306 153988 158312
rect 153948 97306 153976 158306
rect 154132 147665 154160 220079
rect 154118 147656 154174 147665
rect 154118 147591 154174 147600
rect 154224 146266 154252 225626
rect 154316 158710 154344 238886
rect 154408 159254 154436 242150
rect 154488 241528 154540 241534
rect 154488 241470 154540 241476
rect 154396 159248 154448 159254
rect 154396 159190 154448 159196
rect 154304 158704 154356 158710
rect 154304 158646 154356 158652
rect 154500 157282 154528 241470
rect 157246 240952 157302 240961
rect 157246 240887 157302 240896
rect 157062 240680 157118 240689
rect 157062 240615 157118 240624
rect 155684 240168 155736 240174
rect 155684 240110 155736 240116
rect 155498 239456 155554 239465
rect 155498 239391 155554 239400
rect 155408 216028 155460 216034
rect 155408 215970 155460 215976
rect 155224 211880 155276 211886
rect 155224 211822 155276 211828
rect 154488 157276 154540 157282
rect 154488 157218 154540 157224
rect 154578 153096 154634 153105
rect 154578 153031 154634 153040
rect 154212 146260 154264 146266
rect 154212 146202 154264 146208
rect 154488 146260 154540 146266
rect 154488 146202 154540 146208
rect 154500 145654 154528 146202
rect 154488 145648 154540 145654
rect 154488 145590 154540 145596
rect 153936 97300 153988 97306
rect 153936 97242 153988 97248
rect 154592 16574 154620 153031
rect 155236 59362 155264 211822
rect 155420 161474 155448 215970
rect 155328 161446 155448 161474
rect 155328 160177 155356 161446
rect 155512 160478 155540 239391
rect 155592 236700 155644 236706
rect 155592 236642 155644 236648
rect 155500 160472 155552 160478
rect 155500 160414 155552 160420
rect 155314 160168 155370 160177
rect 155314 160103 155370 160112
rect 155328 153785 155356 160103
rect 155512 153921 155540 160414
rect 155604 157049 155632 236642
rect 155696 159905 155724 240110
rect 155774 239728 155830 239737
rect 155774 239663 155830 239672
rect 156512 239692 156564 239698
rect 155682 159896 155738 159905
rect 155682 159831 155738 159840
rect 155590 157040 155646 157049
rect 155590 156975 155646 156984
rect 155498 153912 155554 153921
rect 155498 153847 155554 153856
rect 155314 153776 155370 153785
rect 155314 153711 155370 153720
rect 155604 152522 155632 156975
rect 155788 155786 155816 239663
rect 156512 239634 156564 239640
rect 155866 239592 155922 239601
rect 155866 239527 155922 239536
rect 155880 160682 155908 239527
rect 155868 160676 155920 160682
rect 155868 160618 155920 160624
rect 155776 155780 155828 155786
rect 155776 155722 155828 155728
rect 155592 152516 155644 152522
rect 155592 152458 155644 152464
rect 155788 149705 155816 155722
rect 155880 155242 155908 160618
rect 156524 156641 156552 239634
rect 156972 233912 157024 233918
rect 156972 233854 157024 233860
rect 156696 228948 156748 228954
rect 156696 228890 156748 228896
rect 156604 209908 156656 209914
rect 156604 209850 156656 209856
rect 156510 156632 156566 156641
rect 156510 156567 156566 156576
rect 155868 155236 155920 155242
rect 155868 155178 155920 155184
rect 155960 155236 156012 155242
rect 155960 155178 156012 155184
rect 155774 149696 155830 149705
rect 155774 149631 155830 149640
rect 155224 59356 155276 59362
rect 155224 59298 155276 59304
rect 155972 16574 156000 155178
rect 156616 45558 156644 209850
rect 156708 160041 156736 228890
rect 156788 228880 156840 228886
rect 156788 228822 156840 228828
rect 156694 160032 156750 160041
rect 156694 159967 156750 159976
rect 156800 158817 156828 228822
rect 156880 228812 156932 228818
rect 156880 228754 156932 228760
rect 156892 159526 156920 228754
rect 156984 160449 157012 233854
rect 156970 160440 157026 160449
rect 156970 160375 157026 160384
rect 156880 159520 156932 159526
rect 156880 159462 156932 159468
rect 156892 159361 156920 159462
rect 156878 159352 156934 159361
rect 156878 159287 156934 159296
rect 156786 158808 156842 158817
rect 156786 158743 156842 158752
rect 156696 157956 156748 157962
rect 156696 157898 156748 157904
rect 156708 94518 156736 157898
rect 156800 153882 156828 158743
rect 156878 156632 156934 156641
rect 156878 156567 156934 156576
rect 156788 153876 156840 153882
rect 156788 153818 156840 153824
rect 156892 149734 156920 156567
rect 156984 151201 157012 160375
rect 157076 160274 157104 240615
rect 157064 160268 157116 160274
rect 157064 160210 157116 160216
rect 157260 157321 157288 240887
rect 157812 211177 157840 293218
rect 160008 241596 160060 241602
rect 160008 241538 160060 241544
rect 158444 239556 158496 239562
rect 158444 239498 158496 239504
rect 158350 235376 158406 235385
rect 158350 235311 158406 235320
rect 158258 228304 158314 228313
rect 158258 228239 158314 228248
rect 158166 221504 158222 221513
rect 158166 221439 158222 221448
rect 158076 220108 158128 220114
rect 158076 220050 158128 220056
rect 157984 213308 158036 213314
rect 157984 213250 158036 213256
rect 157892 211200 157944 211206
rect 157798 211168 157854 211177
rect 157892 211142 157944 211148
rect 157798 211103 157854 211112
rect 157800 162308 157852 162314
rect 157800 162250 157852 162256
rect 157812 157865 157840 162250
rect 157904 159390 157932 211142
rect 157996 162194 158024 213250
rect 158088 162314 158116 220050
rect 158076 162308 158128 162314
rect 158076 162250 158128 162256
rect 157996 162166 158116 162194
rect 157892 159384 157944 159390
rect 157892 159326 157944 159332
rect 157890 158536 157946 158545
rect 157890 158471 157946 158480
rect 157338 157856 157394 157865
rect 157338 157791 157394 157800
rect 157798 157856 157854 157865
rect 157798 157791 157854 157800
rect 157246 157312 157302 157321
rect 157246 157247 157302 157256
rect 157352 155281 157380 157791
rect 157430 157448 157486 157457
rect 157430 157383 157486 157392
rect 157338 155272 157394 155281
rect 157338 155207 157394 155216
rect 157444 154057 157472 157383
rect 157430 154048 157486 154057
rect 157430 153983 157486 153992
rect 157338 153776 157394 153785
rect 157338 153711 157394 153720
rect 156970 151192 157026 151201
rect 156970 151127 157026 151136
rect 156880 149728 156932 149734
rect 156880 149670 156932 149676
rect 156696 94512 156748 94518
rect 156696 94454 156748 94460
rect 156604 45552 156656 45558
rect 156604 45494 156656 45500
rect 157352 16574 157380 153711
rect 157904 100026 157932 158471
rect 157984 157412 158036 157418
rect 157984 157354 158036 157360
rect 157892 100020 157944 100026
rect 157892 99962 157944 99968
rect 154592 16546 155448 16574
rect 155972 16546 156184 16574
rect 157352 16546 157840 16574
rect 153844 6860 153896 6866
rect 153844 6802 153896 6808
rect 155420 480 155448 16546
rect 154182 354 154294 480
rect 153764 326 154294 354
rect 154182 -960 154294 326
rect 155378 -960 155490 480
rect 156156 354 156184 16546
rect 157812 480 157840 16546
rect 157996 3466 158024 157354
rect 158088 157321 158116 162166
rect 158180 157593 158208 221439
rect 158272 160313 158300 228239
rect 158258 160304 158314 160313
rect 158258 160239 158314 160248
rect 158166 157584 158222 157593
rect 158166 157519 158222 157528
rect 158074 157312 158130 157321
rect 158074 157247 158130 157256
rect 158180 153105 158208 157519
rect 158166 153096 158222 153105
rect 158166 153031 158222 153040
rect 158272 148345 158300 160239
rect 158364 157457 158392 235311
rect 158456 159662 158484 239498
rect 158536 239488 158588 239494
rect 158536 239430 158588 239436
rect 158444 159656 158496 159662
rect 158444 159598 158496 159604
rect 158548 159458 158576 239430
rect 159916 236768 159968 236774
rect 159916 236710 159968 236716
rect 159822 231704 159878 231713
rect 159822 231639 159878 231648
rect 159640 228744 159692 228750
rect 159640 228686 159692 228692
rect 159546 225584 159602 225593
rect 159546 225519 159602 225528
rect 158628 222964 158680 222970
rect 158628 222906 158680 222912
rect 158536 159452 158588 159458
rect 158536 159394 158588 159400
rect 158640 158137 158668 222906
rect 159364 214668 159416 214674
rect 159364 214610 159416 214616
rect 159272 212084 159324 212090
rect 159272 212026 159324 212032
rect 159284 202842 159312 212026
rect 159272 202836 159324 202842
rect 159272 202778 159324 202784
rect 158720 161152 158772 161158
rect 158720 161094 158772 161100
rect 158732 159225 158760 161094
rect 159376 160585 159404 214610
rect 159456 209432 159508 209438
rect 159456 209374 159508 209380
rect 159362 160576 159418 160585
rect 159362 160511 159418 160520
rect 158718 159216 158774 159225
rect 158718 159151 158774 159160
rect 158626 158128 158682 158137
rect 158626 158063 158682 158072
rect 158350 157448 158406 157457
rect 158350 157383 158406 157392
rect 158258 148336 158314 148345
rect 158258 148271 158314 148280
rect 158732 16574 158760 159151
rect 159376 151337 159404 160511
rect 159468 158681 159496 209374
rect 159560 159866 159588 225519
rect 159652 161158 159680 228686
rect 159732 228472 159784 228478
rect 159732 228414 159784 228420
rect 159640 161152 159692 161158
rect 159640 161094 159692 161100
rect 159548 159860 159600 159866
rect 159548 159802 159600 159808
rect 159454 158672 159510 158681
rect 159454 158607 159510 158616
rect 159744 158001 159772 228414
rect 159730 157992 159786 158001
rect 159730 157927 159786 157936
rect 159744 151774 159772 157927
rect 159836 156913 159864 231639
rect 159928 160070 159956 236710
rect 159916 160064 159968 160070
rect 159916 160006 159968 160012
rect 159916 159860 159968 159866
rect 159916 159802 159968 159808
rect 159928 159390 159956 159802
rect 160020 159662 160048 241538
rect 161112 238332 161164 238338
rect 161112 238274 161164 238280
rect 161020 227112 161072 227118
rect 161020 227054 161072 227060
rect 160928 227044 160980 227050
rect 160928 226986 160980 226992
rect 160836 225616 160888 225622
rect 160836 225558 160888 225564
rect 160744 218748 160796 218754
rect 160744 218690 160796 218696
rect 160560 209976 160612 209982
rect 160560 209918 160612 209924
rect 160572 189038 160600 209918
rect 160652 209228 160704 209234
rect 160652 209170 160704 209176
rect 160560 189032 160612 189038
rect 160560 188974 160612 188980
rect 160664 164218 160692 209170
rect 160652 164212 160704 164218
rect 160652 164154 160704 164160
rect 160558 159760 160614 159769
rect 160558 159695 160614 159704
rect 160008 159656 160060 159662
rect 160008 159598 160060 159604
rect 159916 159384 159968 159390
rect 159916 159326 159968 159332
rect 160006 158672 160062 158681
rect 160006 158607 160062 158616
rect 160020 157729 160048 158607
rect 160572 158302 160600 159695
rect 160560 158296 160612 158302
rect 160560 158238 160612 158244
rect 160006 157720 160062 157729
rect 160756 157690 160784 218690
rect 160848 157894 160876 225558
rect 160836 157888 160888 157894
rect 160836 157830 160888 157836
rect 160006 157655 160062 157664
rect 160744 157684 160796 157690
rect 159822 156904 159878 156913
rect 159822 156839 159878 156848
rect 160020 154578 160048 157655
rect 160744 157626 160796 157632
rect 160940 157622 160968 226986
rect 161032 157758 161060 227054
rect 161124 161945 161152 238274
rect 161204 238128 161256 238134
rect 161204 238070 161256 238076
rect 161110 161936 161166 161945
rect 161110 161871 161166 161880
rect 161216 159254 161244 238070
rect 161296 238060 161348 238066
rect 161296 238002 161348 238008
rect 161308 159526 161336 238002
rect 161940 237516 161992 237522
rect 161940 237458 161992 237464
rect 161388 237448 161440 237454
rect 161388 237390 161440 237396
rect 161296 159520 161348 159526
rect 161296 159462 161348 159468
rect 161204 159248 161256 159254
rect 161204 159190 161256 159196
rect 161400 158914 161428 237390
rect 161480 232552 161532 232558
rect 161480 232494 161532 232500
rect 161388 158908 161440 158914
rect 161388 158850 161440 158856
rect 161492 158030 161520 232494
rect 161572 229016 161624 229022
rect 161572 228958 161624 228964
rect 161584 159186 161612 228958
rect 161664 227180 161716 227186
rect 161664 227122 161716 227128
rect 161676 161566 161704 227122
rect 161756 215960 161808 215966
rect 161756 215902 161808 215908
rect 161664 161560 161716 161566
rect 161664 161502 161716 161508
rect 161572 159180 161624 159186
rect 161572 159122 161624 159128
rect 161480 158024 161532 158030
rect 161480 157966 161532 157972
rect 161020 157752 161072 157758
rect 161020 157694 161072 157700
rect 160928 157616 160980 157622
rect 160928 157558 160980 157564
rect 161388 156392 161440 156398
rect 161388 156334 161440 156340
rect 160744 155984 160796 155990
rect 160744 155926 160796 155932
rect 160020 154550 160140 154578
rect 159732 151768 159784 151774
rect 159732 151710 159784 151716
rect 159362 151328 159418 151337
rect 159362 151263 159418 151272
rect 160112 147674 160140 154550
rect 160112 147646 160232 147674
rect 160098 144800 160154 144809
rect 160098 144735 160154 144744
rect 158732 16546 158944 16574
rect 157984 3460 158036 3466
rect 157984 3402 158036 3408
rect 158916 480 158944 16546
rect 160112 3534 160140 144735
rect 160204 3670 160232 147646
rect 160192 3664 160244 3670
rect 160192 3606 160244 3612
rect 160100 3528 160152 3534
rect 160100 3470 160152 3476
rect 160756 3466 160784 155926
rect 161400 144809 161428 156334
rect 161480 151768 161532 151774
rect 161480 151710 161532 151716
rect 161386 144800 161442 144809
rect 161386 144735 161442 144744
rect 161296 3528 161348 3534
rect 161296 3470 161348 3476
rect 160744 3460 160796 3466
rect 160744 3402 160796 3408
rect 160100 3256 160152 3262
rect 160100 3198 160152 3204
rect 160112 480 160140 3198
rect 161308 480 161336 3470
rect 161492 3262 161520 151710
rect 161584 144226 161612 159122
rect 161676 146946 161704 161502
rect 161768 159934 161796 215902
rect 161848 160200 161900 160206
rect 161848 160142 161900 160148
rect 161756 159928 161808 159934
rect 161756 159870 161808 159876
rect 161664 146940 161716 146946
rect 161664 146882 161716 146888
rect 161572 144220 161624 144226
rect 161572 144162 161624 144168
rect 161768 135930 161796 159870
rect 161860 159118 161888 160142
rect 161848 159112 161900 159118
rect 161848 159054 161900 159060
rect 161860 155718 161888 159054
rect 161952 158846 161980 237458
rect 162032 228404 162084 228410
rect 162032 228346 162084 228352
rect 161940 158840 161992 158846
rect 161940 158782 161992 158788
rect 162044 157826 162072 228346
rect 163504 225752 163556 225758
rect 163504 225694 163556 225700
rect 162308 222896 162360 222902
rect 162308 222838 162360 222844
rect 162216 221468 162268 221474
rect 162216 221410 162268 221416
rect 162124 160676 162176 160682
rect 162124 160618 162176 160624
rect 162136 160002 162164 160618
rect 162124 159996 162176 160002
rect 162124 159938 162176 159944
rect 162122 159896 162178 159905
rect 162122 159831 162178 159840
rect 162032 157820 162084 157826
rect 162032 157762 162084 157768
rect 162136 157214 162164 159831
rect 162228 158302 162256 221410
rect 162320 158506 162348 222838
rect 163516 215294 163544 225694
rect 163516 215266 163636 215294
rect 162584 211268 162636 211274
rect 162584 211210 162636 211216
rect 162596 211177 162624 211210
rect 162582 211168 162638 211177
rect 162582 211103 162638 211112
rect 163608 209438 163636 215266
rect 164252 212294 164280 294578
rect 165896 294432 165948 294438
rect 165896 294374 165948 294380
rect 165712 294160 165764 294166
rect 165712 294102 165764 294108
rect 164884 293344 164936 293350
rect 164884 293286 164936 293292
rect 164332 293072 164384 293078
rect 164332 293014 164384 293020
rect 164344 229094 164372 293014
rect 164344 229066 164464 229094
rect 164240 212288 164292 212294
rect 164240 212230 164292 212236
rect 164330 211304 164386 211313
rect 164330 211239 164386 211248
rect 164344 209916 164372 211239
rect 164436 209930 164464 229066
rect 164792 212288 164844 212294
rect 164792 212230 164844 212236
rect 164804 209930 164832 212230
rect 164896 211177 164924 293286
rect 165344 217388 165396 217394
rect 165344 217330 165396 217336
rect 164882 211168 164938 211177
rect 164882 211103 164938 211112
rect 164436 209902 164726 209930
rect 164804 209902 165094 209930
rect 165356 209681 165384 217330
rect 165724 212294 165752 294102
rect 165802 275224 165858 275233
rect 165802 275159 165858 275168
rect 165712 212288 165764 212294
rect 165712 212230 165764 212236
rect 165712 211948 165764 211954
rect 165712 211890 165764 211896
rect 165434 211168 165490 211177
rect 165434 211103 165490 211112
rect 165448 209916 165476 211103
rect 165724 209930 165752 211890
rect 165816 210338 165844 275159
rect 165908 211954 165936 294374
rect 166816 217320 166868 217326
rect 166816 217262 166868 217268
rect 165896 211948 165948 211954
rect 165896 211890 165948 211896
rect 166540 211268 166592 211274
rect 166540 211210 166592 211216
rect 165816 210310 165936 210338
rect 165908 209930 165936 210310
rect 165724 209902 165830 209930
rect 165908 209902 166198 209930
rect 166552 209916 166580 211210
rect 166828 209681 166856 217262
rect 167012 214538 167040 294782
rect 168380 294772 168432 294778
rect 168380 294714 168432 294720
rect 168288 290692 168340 290698
rect 168288 290634 168340 290640
rect 167092 244928 167144 244934
rect 167092 244870 167144 244876
rect 167000 214532 167052 214538
rect 167000 214474 167052 214480
rect 166908 212288 166960 212294
rect 166908 212230 166960 212236
rect 166920 209916 166948 212230
rect 167104 209930 167132 244870
rect 167736 214532 167788 214538
rect 167736 214474 167788 214480
rect 167644 211744 167696 211750
rect 167644 211686 167696 211692
rect 167104 209902 167302 209930
rect 167656 209916 167684 211686
rect 167748 209930 167776 214474
rect 168300 211750 168328 290634
rect 168392 214538 168420 294714
rect 169668 286340 169720 286346
rect 169668 286282 169720 286288
rect 168470 278080 168526 278089
rect 168470 278015 168526 278024
rect 168380 214532 168432 214538
rect 168380 214474 168432 214480
rect 168288 211744 168340 211750
rect 168288 211686 168340 211692
rect 168300 211274 168328 211686
rect 168288 211268 168340 211274
rect 168288 211210 168340 211216
rect 168484 209930 168512 278015
rect 168564 247716 168616 247722
rect 168564 247658 168616 247664
rect 168576 229094 168604 247658
rect 168576 229066 169248 229094
rect 168840 214532 168892 214538
rect 168840 214474 168892 214480
rect 168748 211404 168800 211410
rect 168748 211346 168800 211352
rect 167748 209902 168038 209930
rect 168406 209902 168512 209930
rect 168760 209916 168788 211346
rect 168852 209930 168880 214474
rect 169220 209930 169248 229066
rect 169680 211410 169708 286282
rect 169772 214538 169800 296006
rect 171140 295588 171192 295594
rect 171140 295530 171192 295536
rect 169852 294364 169904 294370
rect 169852 294306 169904 294312
rect 169760 214532 169812 214538
rect 169760 214474 169812 214480
rect 169668 211404 169720 211410
rect 169668 211346 169720 211352
rect 169760 211336 169812 211342
rect 169760 211278 169812 211284
rect 169772 209930 169800 211278
rect 169864 210066 169892 294306
rect 169944 290828 169996 290834
rect 169944 290770 169996 290776
rect 169956 229094 169984 290770
rect 169956 229066 170720 229094
rect 170312 214532 170364 214538
rect 170312 214474 170364 214480
rect 169864 210038 169984 210066
rect 169956 209930 169984 210038
rect 170324 209930 170352 214474
rect 170692 209930 170720 229066
rect 171152 214538 171180 295530
rect 172520 295520 172572 295526
rect 172520 295462 172572 295468
rect 171232 294500 171284 294506
rect 171232 294442 171284 294448
rect 171140 214532 171192 214538
rect 171140 214474 171192 214480
rect 171244 209930 171272 294442
rect 171322 287736 171378 287745
rect 171322 287671 171378 287680
rect 171336 229094 171364 287671
rect 172336 233980 172388 233986
rect 172336 233922 172388 233928
rect 171336 229066 171456 229094
rect 171428 209930 171456 229066
rect 172348 219434 172376 233922
rect 171980 219406 172376 219434
rect 168852 209902 169142 209930
rect 169220 209902 169510 209930
rect 169772 209902 169878 209930
rect 169956 209902 170246 209930
rect 170324 209902 170614 209930
rect 170692 209902 170982 209930
rect 171244 209902 171350 209930
rect 171428 209902 171718 209930
rect 165342 209672 165398 209681
rect 165342 209607 165398 209616
rect 166814 209672 166870 209681
rect 166814 209607 166870 209616
rect 171980 209545 172008 219406
rect 172532 214538 172560 295462
rect 172704 293140 172756 293146
rect 172704 293082 172756 293088
rect 172612 292868 172664 292874
rect 172612 292810 172664 292816
rect 172152 214532 172204 214538
rect 172152 214474 172204 214480
rect 172520 214532 172572 214538
rect 172520 214474 172572 214480
rect 172060 211948 172112 211954
rect 172060 211890 172112 211896
rect 172072 209916 172100 211890
rect 172164 209930 172192 214474
rect 172624 209930 172652 292810
rect 172716 229094 172744 293082
rect 173808 290760 173860 290766
rect 173808 290702 173860 290708
rect 172716 229066 172928 229094
rect 172900 209930 172928 229066
rect 173256 214532 173308 214538
rect 173256 214474 173308 214480
rect 173268 209930 173296 214474
rect 173820 212226 173848 290702
rect 173912 214742 173940 296890
rect 173992 295656 174044 295662
rect 173992 295598 174044 295604
rect 173900 214736 173952 214742
rect 173900 214678 173952 214684
rect 174004 214538 174032 295598
rect 175280 292800 175332 292806
rect 175280 292742 175332 292748
rect 174084 289332 174136 289338
rect 174084 289274 174136 289280
rect 173992 214532 174044 214538
rect 173992 214474 174044 214480
rect 173900 212424 173952 212430
rect 173900 212366 173952 212372
rect 173532 212220 173584 212226
rect 173532 212162 173584 212168
rect 173808 212220 173860 212226
rect 173808 212162 173860 212168
rect 173544 211342 173572 212162
rect 173532 211336 173584 211342
rect 173532 211278 173584 211284
rect 172164 209902 172454 209930
rect 172624 209902 172822 209930
rect 172900 209902 173190 209930
rect 173268 209902 173558 209930
rect 173912 209916 173940 212366
rect 174096 209930 174124 289274
rect 175292 229094 175320 292742
rect 175292 229066 176240 229094
rect 174728 214736 174780 214742
rect 174728 214678 174780 214684
rect 176108 214736 176160 214742
rect 176108 214678 176160 214684
rect 174360 214532 174412 214538
rect 174360 214474 174412 214480
rect 174372 209930 174400 214474
rect 174740 209930 174768 214678
rect 175740 212492 175792 212498
rect 175740 212434 175792 212440
rect 175372 212152 175424 212158
rect 175372 212094 175424 212100
rect 174096 209902 174294 209930
rect 174372 209902 174662 209930
rect 174740 209902 175030 209930
rect 175384 209916 175412 212094
rect 175752 209916 175780 212434
rect 176120 209916 176148 214678
rect 176212 209930 176240 229066
rect 176672 212362 176700 297026
rect 176752 295724 176804 295730
rect 176752 295666 176804 295672
rect 176660 212356 176712 212362
rect 176660 212298 176712 212304
rect 176764 212106 176792 295666
rect 176844 294228 176896 294234
rect 176844 294170 176896 294176
rect 176856 212294 176884 294170
rect 176936 292936 176988 292942
rect 176936 292878 176988 292884
rect 176948 229094 176976 292878
rect 178040 289876 178092 289882
rect 178040 289818 178092 289824
rect 176948 229066 177344 229094
rect 176936 212356 176988 212362
rect 176936 212298 176988 212304
rect 176844 212288 176896 212294
rect 176844 212230 176896 212236
rect 176764 212078 176884 212106
rect 176212 209902 176502 209930
rect 176856 209916 176884 212078
rect 176948 209930 176976 212298
rect 177316 209930 177344 229066
rect 178052 212294 178080 289818
rect 178132 279472 178184 279478
rect 178132 279414 178184 279420
rect 177672 212288 177724 212294
rect 177672 212230 177724 212236
rect 178040 212288 178092 212294
rect 178040 212230 178092 212236
rect 177684 209930 177712 212230
rect 178144 209930 178172 279414
rect 178696 212430 178724 297230
rect 187700 297220 187752 297226
rect 187700 297162 187752 297168
rect 183560 296812 183612 296818
rect 183560 296754 183612 296760
rect 182180 294296 182232 294302
rect 182180 294238 182232 294244
rect 179420 293004 179472 293010
rect 179420 292946 179472 292952
rect 179432 215294 179460 292946
rect 180064 289264 180116 289270
rect 180064 289206 180116 289212
rect 179512 280832 179564 280838
rect 179512 280774 179564 280780
rect 179524 229094 179552 280774
rect 179524 229066 179736 229094
rect 179432 215266 179644 215294
rect 178684 212424 178736 212430
rect 178684 212366 178736 212372
rect 178776 212288 178828 212294
rect 178776 212230 178828 212236
rect 178592 211744 178644 211750
rect 178592 211686 178644 211692
rect 178604 209930 178632 211686
rect 178684 211336 178736 211342
rect 178684 211278 178736 211284
rect 178696 210594 178724 211278
rect 178684 210588 178736 210594
rect 178684 210530 178736 210536
rect 178788 209930 178816 212230
rect 179616 210934 179644 215266
rect 179604 210928 179656 210934
rect 179604 210870 179656 210876
rect 179708 210066 179736 229066
rect 180076 212498 180104 289206
rect 180800 283620 180852 283626
rect 180800 283562 180852 283568
rect 180812 229094 180840 283562
rect 180812 229066 181392 229094
rect 180156 217456 180208 217462
rect 180156 217398 180208 217404
rect 180064 212492 180116 212498
rect 180064 212434 180116 212440
rect 179788 210928 179840 210934
rect 179788 210870 179840 210876
rect 179616 210038 179736 210066
rect 179616 209930 179644 210038
rect 176948 209902 177238 209930
rect 177316 209902 177606 209930
rect 177684 209902 177974 209930
rect 178144 209902 178342 209930
rect 178604 209902 178710 209930
rect 178788 209902 179078 209930
rect 179446 209902 179644 209930
rect 179800 209916 179828 210870
rect 180168 209916 180196 217398
rect 181260 212424 181312 212430
rect 181260 212366 181312 212372
rect 180890 212120 180946 212129
rect 180890 212055 180946 212064
rect 180524 212016 180576 212022
rect 180524 211958 180576 211964
rect 180536 209916 180564 211958
rect 180904 209916 180932 212055
rect 181272 209916 181300 212366
rect 181364 209930 181392 229066
rect 182192 215294 182220 294238
rect 182272 290420 182324 290426
rect 182272 290362 182324 290368
rect 182284 229094 182312 290362
rect 182284 229066 183232 229094
rect 182192 215266 182496 215294
rect 182364 213444 182416 213450
rect 182364 213386 182416 213392
rect 181996 213376 182048 213382
rect 181996 213318 182048 213324
rect 181364 209902 181654 209930
rect 182008 209916 182036 213318
rect 182376 209916 182404 213386
rect 182468 209930 182496 215266
rect 183100 210588 183152 210594
rect 183100 210530 183152 210536
rect 182468 209902 182758 209930
rect 183112 209916 183140 210530
rect 183204 209930 183232 229066
rect 183572 212362 183600 296754
rect 184202 289776 184258 289785
rect 184202 289711 184258 289720
rect 183652 289196 183704 289202
rect 183652 289138 183704 289144
rect 183560 212356 183612 212362
rect 183560 212298 183612 212304
rect 183664 212294 183692 289138
rect 183744 282192 183796 282198
rect 183744 282134 183796 282140
rect 183756 229094 183784 282134
rect 183756 229066 183876 229094
rect 183652 212288 183704 212294
rect 183652 212230 183704 212236
rect 183204 209902 183494 209930
rect 183848 209916 183876 229066
rect 184216 212430 184244 289711
rect 186502 289640 186558 289649
rect 186502 289575 186558 289584
rect 186318 289232 186374 289241
rect 186318 289167 186374 289176
rect 184940 289128 184992 289134
rect 184940 289070 184992 289076
rect 185030 289096 185086 289105
rect 184848 234048 184900 234054
rect 184848 233990 184900 233996
rect 184756 213240 184808 213246
rect 184756 213182 184808 213188
rect 184204 212424 184256 212430
rect 184204 212366 184256 212372
rect 184388 212424 184440 212430
rect 184388 212366 184440 212372
rect 184296 212356 184348 212362
rect 184296 212298 184348 212304
rect 183928 212288 183980 212294
rect 183928 212230 183980 212236
rect 183940 209930 183968 212230
rect 184308 209930 184336 212298
rect 184400 210526 184428 212366
rect 184388 210520 184440 210526
rect 184388 210462 184440 210468
rect 183940 209902 184230 209930
rect 184308 209902 184598 209930
rect 184768 209545 184796 213182
rect 184860 209681 184888 233990
rect 184952 212362 184980 289070
rect 185030 289031 185086 289040
rect 184940 212356 184992 212362
rect 184940 212298 184992 212304
rect 184940 210792 184992 210798
rect 184940 210734 184992 210740
rect 184952 209916 184980 210734
rect 185044 209794 185072 289031
rect 185124 284980 185176 284986
rect 185124 284922 185176 284928
rect 185136 212294 185164 284922
rect 185216 239624 185268 239630
rect 185216 239566 185268 239572
rect 185124 212288 185176 212294
rect 185124 212230 185176 212236
rect 185228 210798 185256 239566
rect 186332 214470 186360 289167
rect 186412 273964 186464 273970
rect 186412 273906 186464 273912
rect 186424 214538 186452 273906
rect 186412 214532 186464 214538
rect 186412 214474 186464 214480
rect 186320 214464 186372 214470
rect 186320 214406 186372 214412
rect 186412 214396 186464 214402
rect 186412 214338 186464 214344
rect 185400 212356 185452 212362
rect 185400 212298 185452 212304
rect 185216 210792 185268 210798
rect 185216 210734 185268 210740
rect 185412 209930 185440 212298
rect 185768 212288 185820 212294
rect 185768 212230 185820 212236
rect 185860 212288 185912 212294
rect 185860 212230 185912 212236
rect 185780 209930 185808 212230
rect 185872 211750 185900 212230
rect 185860 211744 185912 211750
rect 185860 211686 185912 211692
rect 185412 209902 185702 209930
rect 185780 209902 186070 209930
rect 186424 209916 186452 214338
rect 186516 209794 186544 289575
rect 186686 289504 186742 289513
rect 186686 289439 186742 289448
rect 186700 214402 186728 289439
rect 186872 214532 186924 214538
rect 186872 214474 186924 214480
rect 186688 214396 186740 214402
rect 186688 214338 186740 214344
rect 186884 209930 186912 214474
rect 187240 214464 187292 214470
rect 187240 214406 187292 214412
rect 187252 209930 187280 214406
rect 187332 211404 187384 211410
rect 187332 211346 187384 211352
rect 187344 210089 187372 211346
rect 187330 210080 187386 210089
rect 187330 210015 187386 210024
rect 187712 209930 187740 297162
rect 189080 296880 189132 296886
rect 189080 296822 189132 296828
rect 188344 293208 188396 293214
rect 188344 293150 188396 293156
rect 187790 289368 187846 289377
rect 187790 289303 187846 289312
rect 187804 214538 187832 289303
rect 187884 242276 187936 242282
rect 187884 242218 187936 242224
rect 187896 229094 187924 242218
rect 187896 229066 188016 229094
rect 187792 214532 187844 214538
rect 187792 214474 187844 214480
rect 187792 211404 187844 211410
rect 187792 211346 187844 211352
rect 187804 210458 187832 211346
rect 187792 210452 187844 210458
rect 187792 210394 187844 210400
rect 187988 209930 188016 229066
rect 188356 212294 188384 293150
rect 188896 234116 188948 234122
rect 188896 234058 188948 234064
rect 188620 216096 188672 216102
rect 188620 216038 188672 216044
rect 188344 212288 188396 212294
rect 188344 212230 188396 212236
rect 186884 209902 187174 209930
rect 187252 209902 187542 209930
rect 187712 209902 187910 209930
rect 187988 209902 188278 209930
rect 188632 209916 188660 216038
rect 188804 212220 188856 212226
rect 188804 212162 188856 212168
rect 185044 209766 185334 209794
rect 186516 209766 186806 209794
rect 188816 209681 188844 212162
rect 184846 209672 184902 209681
rect 184846 209607 184902 209616
rect 188802 209672 188858 209681
rect 188802 209607 188858 209616
rect 188908 209545 188936 234058
rect 189092 214538 189120 296822
rect 190460 295452 190512 295458
rect 190460 295394 190512 295400
rect 189170 290728 189226 290737
rect 189170 290663 189226 290672
rect 188988 214532 189040 214538
rect 188988 214474 189040 214480
rect 189080 214532 189132 214538
rect 189080 214474 189132 214480
rect 189000 209916 189028 214474
rect 189184 214470 189212 290663
rect 189264 272536 189316 272542
rect 189264 272478 189316 272484
rect 189276 229094 189304 272478
rect 189276 229066 189396 229094
rect 189172 214464 189224 214470
rect 189172 214406 189224 214412
rect 189368 209916 189396 229066
rect 190472 214538 190500 295394
rect 192022 290592 192078 290601
rect 192022 290527 192078 290536
rect 191932 290488 191984 290494
rect 191932 290430 191984 290436
rect 190550 290048 190606 290057
rect 190550 289983 190606 289992
rect 189816 214532 189868 214538
rect 189816 214474 189868 214480
rect 190460 214532 190512 214538
rect 190460 214474 190512 214480
rect 189448 214464 189500 214470
rect 189448 214406 189500 214412
rect 189460 209930 189488 214406
rect 189828 209930 189856 214474
rect 190564 214470 190592 289983
rect 191838 289912 191894 289921
rect 191838 289847 191894 289856
rect 190642 276720 190698 276729
rect 190642 276655 190698 276664
rect 190552 214464 190604 214470
rect 190552 214406 190604 214412
rect 189460 209902 189750 209930
rect 189828 209902 190118 209930
rect 190656 209794 190684 276655
rect 190734 243536 190790 243545
rect 190734 243471 190790 243480
rect 190748 229094 190776 243471
rect 191656 238672 191708 238678
rect 191656 238614 191708 238620
rect 191668 232558 191696 238614
rect 191748 232756 191800 232762
rect 191748 232698 191800 232704
rect 191656 232552 191708 232558
rect 191656 232494 191708 232500
rect 190748 229066 191328 229094
rect 190920 214532 190972 214538
rect 190920 214474 190972 214480
rect 190736 214464 190788 214470
rect 190736 214406 190788 214412
rect 190748 209930 190776 214406
rect 190932 209930 190960 214474
rect 191300 209930 191328 229066
rect 190748 209902 190854 209930
rect 190932 209902 191222 209930
rect 191300 209902 191590 209930
rect 190486 209766 190684 209794
rect 191760 209545 191788 232698
rect 191852 209930 191880 289847
rect 191944 214538 191972 290430
rect 191932 214532 191984 214538
rect 191932 214474 191984 214480
rect 192036 209930 192064 290527
rect 192114 286376 192170 286385
rect 192114 286311 192170 286320
rect 192128 229094 192156 286311
rect 192484 238264 192536 238270
rect 192484 238206 192536 238212
rect 192496 232801 192524 238206
rect 192482 232792 192538 232801
rect 192482 232727 192538 232736
rect 193128 232552 193180 232558
rect 193128 232494 193180 232500
rect 192128 229066 192432 229094
rect 192404 209930 192432 229066
rect 193140 219434 193168 232494
rect 192956 219406 193168 219434
rect 191852 209902 191958 209930
rect 192036 209902 192326 209930
rect 192404 209902 192694 209930
rect 192956 209545 192984 219406
rect 193036 214532 193088 214538
rect 193036 214474 193088 214480
rect 193048 209916 193076 214474
rect 193232 214470 193260 300086
rect 194600 299532 194652 299538
rect 194600 299474 194652 299480
rect 193404 298240 193456 298246
rect 193404 298182 193456 298188
rect 193312 298172 193364 298178
rect 193312 298114 193364 298120
rect 193324 214538 193352 298114
rect 193312 214532 193364 214538
rect 193312 214474 193364 214480
rect 193220 214464 193272 214470
rect 193220 214406 193272 214412
rect 193416 209916 193444 298182
rect 193772 238400 193824 238406
rect 193772 238342 193824 238348
rect 193784 233209 193812 238342
rect 193770 233200 193826 233209
rect 193770 233135 193826 233144
rect 194416 232688 194468 232694
rect 194416 232630 194468 232636
rect 193496 214532 193548 214538
rect 193496 214474 193548 214480
rect 193508 209930 193536 214474
rect 194140 212220 194192 212226
rect 194140 212162 194192 212168
rect 193508 209902 193798 209930
rect 194152 209916 194180 212162
rect 194428 209545 194456 232630
rect 194612 214538 194640 299474
rect 195980 297016 196032 297022
rect 195980 296958 196032 296964
rect 194692 290556 194744 290562
rect 194692 290498 194744 290504
rect 194600 214532 194652 214538
rect 194600 214474 194652 214480
rect 194704 214470 194732 290498
rect 194784 271176 194836 271182
rect 194784 271118 194836 271124
rect 194796 229094 194824 271118
rect 195888 231872 195940 231878
rect 195888 231814 195940 231820
rect 194796 229066 194916 229094
rect 194508 214464 194560 214470
rect 194508 214406 194560 214412
rect 194692 214464 194744 214470
rect 194692 214406 194744 214412
rect 194520 209916 194548 214406
rect 194888 209916 194916 229066
rect 195336 214532 195388 214538
rect 195336 214474 195388 214480
rect 194968 214464 195020 214470
rect 194968 214406 195020 214412
rect 194980 209930 195008 214406
rect 195348 209930 195376 214474
rect 194980 209902 195270 209930
rect 195348 209902 195638 209930
rect 195900 209545 195928 231814
rect 195992 212294 196020 296958
rect 196072 290080 196124 290086
rect 196072 290022 196124 290028
rect 195980 212288 196032 212294
rect 195980 212230 196032 212236
rect 195980 211744 196032 211750
rect 195980 211686 196032 211692
rect 195992 209916 196020 211686
rect 196084 209794 196112 290022
rect 196164 269816 196216 269822
rect 196164 269758 196216 269764
rect 196176 211750 196204 269758
rect 197268 236836 197320 236842
rect 197268 236778 197320 236784
rect 196992 231124 197044 231130
rect 196992 231066 197044 231072
rect 197004 219434 197032 231066
rect 197176 230648 197228 230654
rect 197176 230590 197228 230596
rect 196912 219406 197032 219434
rect 196440 212288 196492 212294
rect 196440 212230 196492 212236
rect 196164 211744 196216 211750
rect 196164 211686 196216 211692
rect 196256 211268 196308 211274
rect 196256 211210 196308 211216
rect 196268 210089 196296 211210
rect 196254 210080 196310 210089
rect 196254 210015 196310 210024
rect 196452 209930 196480 212230
rect 196452 209902 196742 209930
rect 196084 209766 196374 209794
rect 196912 209545 196940 219406
rect 197188 215294 197216 230590
rect 197004 215266 197216 215294
rect 197004 209681 197032 215266
rect 197084 212356 197136 212362
rect 197084 212298 197136 212304
rect 197096 209916 197124 212298
rect 196990 209672 197046 209681
rect 196990 209607 197046 209616
rect 197280 209545 197308 236778
rect 197372 212294 197400 318786
rect 201316 317008 201368 317014
rect 201316 316950 201368 316956
rect 200028 311364 200080 311370
rect 200028 311306 200080 311312
rect 197452 301028 197504 301034
rect 197452 300970 197504 300976
rect 197360 212288 197412 212294
rect 197360 212230 197412 212236
rect 197360 211132 197412 211138
rect 197360 211074 197412 211080
rect 197372 209930 197400 211074
rect 197464 210338 197492 300970
rect 198740 293480 198792 293486
rect 198740 293422 198792 293428
rect 198752 292602 198780 293422
rect 198740 292596 198792 292602
rect 198740 292538 198792 292544
rect 197544 290148 197596 290154
rect 197544 290090 197596 290096
rect 197556 211138 197584 290090
rect 198648 230512 198700 230518
rect 198648 230454 198700 230460
rect 197912 228540 197964 228546
rect 197912 228482 197964 228488
rect 197544 211132 197596 211138
rect 197544 211074 197596 211080
rect 197464 210310 197584 210338
rect 197556 209930 197584 210310
rect 197924 209930 197952 228482
rect 198660 219434 198688 230454
rect 198476 219406 198688 219434
rect 198372 210044 198424 210050
rect 198372 209986 198424 209992
rect 197372 209902 197478 209930
rect 197556 209902 197846 209930
rect 197924 209902 198214 209930
rect 198384 209846 198412 209986
rect 198372 209840 198424 209846
rect 198372 209782 198424 209788
rect 198476 209681 198504 219406
rect 198556 212288 198608 212294
rect 198556 212230 198608 212236
rect 198568 209916 198596 212230
rect 198752 209930 198780 292538
rect 199936 253972 199988 253978
rect 199936 253914 199988 253920
rect 198832 246356 198884 246362
rect 198832 246298 198884 246304
rect 198844 210066 198872 246298
rect 199384 240780 199436 240786
rect 199384 240722 199436 240728
rect 198924 239420 198976 239426
rect 198924 239362 198976 239368
rect 198936 212294 198964 239362
rect 199016 231804 199068 231810
rect 199016 231746 199068 231752
rect 199028 231266 199056 231746
rect 199016 231260 199068 231266
rect 199016 231202 199068 231208
rect 199396 212498 199424 240722
rect 199948 240242 199976 253914
rect 199936 240236 199988 240242
rect 199936 240178 199988 240184
rect 200040 231810 200068 311306
rect 200764 290624 200816 290630
rect 200764 290566 200816 290572
rect 200304 240236 200356 240242
rect 200304 240178 200356 240184
rect 200028 231804 200080 231810
rect 200028 231746 200080 231752
rect 199844 231600 199896 231606
rect 199844 231542 199896 231548
rect 199752 230580 199804 230586
rect 199752 230522 199804 230528
rect 199384 212492 199436 212498
rect 199384 212434 199436 212440
rect 198924 212288 198976 212294
rect 198924 212230 198976 212236
rect 198844 210038 199056 210066
rect 199028 209930 199056 210038
rect 198752 209902 198950 209930
rect 199028 209902 199318 209930
rect 198462 209672 198518 209681
rect 198462 209607 198518 209616
rect 171966 209536 172022 209545
rect 171966 209471 172022 209480
rect 184754 209536 184810 209545
rect 184754 209471 184810 209480
rect 188894 209536 188950 209545
rect 188894 209471 188950 209480
rect 191746 209536 191802 209545
rect 191746 209471 191802 209480
rect 192942 209536 192998 209545
rect 192942 209471 192998 209480
rect 194414 209536 194470 209545
rect 194414 209471 194470 209480
rect 195886 209536 195942 209545
rect 195886 209471 195942 209480
rect 196898 209536 196954 209545
rect 196898 209471 196954 209480
rect 197266 209536 197322 209545
rect 199396 209522 199424 212434
rect 199568 209908 199620 209914
rect 199568 209850 199620 209856
rect 199580 209681 199608 209850
rect 199566 209672 199622 209681
rect 199764 209658 199792 230522
rect 199856 209794 199884 231542
rect 199936 230716 199988 230722
rect 199936 230658 199988 230664
rect 199948 209914 199976 230658
rect 200212 228608 200264 228614
rect 200212 228550 200264 228556
rect 200028 212288 200080 212294
rect 200028 212230 200080 212236
rect 200040 209916 200068 212230
rect 200224 210866 200252 228550
rect 200212 210860 200264 210866
rect 200212 210802 200264 210808
rect 200224 209982 200252 210802
rect 200212 209976 200264 209982
rect 200212 209918 200264 209924
rect 200316 209930 200344 240178
rect 200776 214606 200804 290566
rect 201224 229424 201276 229430
rect 201224 229366 201276 229372
rect 200764 214600 200816 214606
rect 200764 214542 200816 214548
rect 199936 209908 199988 209914
rect 200316 209902 200422 209930
rect 200776 209916 200804 214542
rect 201236 212242 201264 229366
rect 201328 226273 201356 316950
rect 201314 226264 201370 226273
rect 201314 226199 201370 226208
rect 201420 213926 201448 321574
rect 202786 321535 202842 321544
rect 202604 311500 202656 311506
rect 202604 311442 202656 311448
rect 202512 307216 202564 307222
rect 202512 307158 202564 307164
rect 202144 300960 202196 300966
rect 202144 300902 202196 300908
rect 201500 290012 201552 290018
rect 201500 289954 201552 289960
rect 201512 229094 201540 289954
rect 201512 229066 201724 229094
rect 201408 213920 201460 213926
rect 201408 213862 201460 213868
rect 201420 213314 201448 213862
rect 201408 213308 201460 213314
rect 201408 213250 201460 213256
rect 201236 212214 201540 212242
rect 201236 212090 201264 212214
rect 201224 212084 201276 212090
rect 201224 212026 201276 212032
rect 201132 210860 201184 210866
rect 201132 210802 201184 210808
rect 201144 209916 201172 210802
rect 201512 209916 201540 212214
rect 199936 209850 199988 209856
rect 199856 209766 199976 209794
rect 199842 209672 199898 209681
rect 199764 209630 199842 209658
rect 199566 209607 199622 209616
rect 199842 209607 199898 209616
rect 199948 209545 199976 209766
rect 199934 209536 199990 209545
rect 199396 209494 199686 209522
rect 197266 209471 197322 209480
rect 199934 209471 199990 209480
rect 201696 209438 201724 229066
rect 202156 211410 202184 300902
rect 202524 238754 202552 307158
rect 202340 238726 202552 238754
rect 202340 234394 202368 238726
rect 202616 234546 202644 311442
rect 202696 302252 202748 302258
rect 202696 302194 202748 302200
rect 202524 234518 202644 234546
rect 202328 234388 202380 234394
rect 202328 234330 202380 234336
rect 202524 231713 202552 234518
rect 202604 234388 202656 234394
rect 202604 234330 202656 234336
rect 202616 233986 202644 234330
rect 202604 233980 202656 233986
rect 202604 233922 202656 233928
rect 202510 231704 202566 231713
rect 202510 231639 202566 231648
rect 202328 228676 202380 228682
rect 202328 228618 202380 228624
rect 202144 211404 202196 211410
rect 202144 211346 202196 211352
rect 202156 209930 202184 211346
rect 202340 211206 202368 228618
rect 202708 212090 202736 302194
rect 202800 219337 202828 321535
rect 206652 319320 206704 319326
rect 206652 319262 206704 319268
rect 206560 318912 206612 318918
rect 206560 318854 206612 318860
rect 205456 312656 205508 312662
rect 205456 312598 205508 312604
rect 204168 311160 204220 311166
rect 204168 311102 204220 311108
rect 204076 305040 204128 305046
rect 204076 304982 204128 304988
rect 203064 297424 203116 297430
rect 203064 297366 203116 297372
rect 202972 297152 203024 297158
rect 202972 297094 203024 297100
rect 202786 219328 202842 219337
rect 202786 219263 202842 219272
rect 202800 218929 202828 219263
rect 202786 218920 202842 218929
rect 202786 218855 202842 218864
rect 202696 212084 202748 212090
rect 202696 212026 202748 212032
rect 202708 211818 202736 212026
rect 202696 211812 202748 211818
rect 202696 211754 202748 211760
rect 202328 211200 202380 211206
rect 202328 211142 202380 211148
rect 202340 209930 202368 211142
rect 202984 209930 203012 297094
rect 203076 229094 203104 297366
rect 203984 296744 204036 296750
rect 203984 296686 204036 296692
rect 203996 235793 204024 296686
rect 203982 235784 204038 235793
rect 203982 235719 204038 235728
rect 203996 235521 204024 235719
rect 203982 235512 204038 235521
rect 203982 235447 204038 235456
rect 203076 229066 203196 229094
rect 202156 209902 202262 209930
rect 202340 209902 202630 209930
rect 202892 209916 203012 209930
rect 202892 209902 202998 209916
rect 202892 209506 202920 209902
rect 203168 209574 203196 229066
rect 204088 212090 204116 304982
rect 204180 218006 204208 311102
rect 204902 307592 204958 307601
rect 204902 307527 204958 307536
rect 204444 300892 204496 300898
rect 204444 300834 204496 300840
rect 204352 299600 204404 299606
rect 204352 299542 204404 299548
rect 204168 218000 204220 218006
rect 204168 217942 204220 217948
rect 204180 217394 204208 217942
rect 204168 217388 204220 217394
rect 204168 217330 204220 217336
rect 203340 212084 203392 212090
rect 203340 212026 203392 212032
rect 204076 212084 204128 212090
rect 204076 212026 204128 212032
rect 203352 209916 203380 212026
rect 204088 211886 204116 212026
rect 204076 211880 204128 211886
rect 204076 211822 204128 211828
rect 203708 211812 203760 211818
rect 203708 211754 203760 211760
rect 203720 211342 203748 211754
rect 203708 211336 203760 211342
rect 203708 211278 203760 211284
rect 203720 209916 203748 211278
rect 204364 210050 204392 299542
rect 204352 210044 204404 210050
rect 204352 209986 204404 209992
rect 204260 209840 204312 209846
rect 204456 209794 204484 300834
rect 204916 241602 204944 307527
rect 205364 303000 205416 303006
rect 205364 302942 205416 302948
rect 205272 300212 205324 300218
rect 205272 300154 205324 300160
rect 204904 241596 204956 241602
rect 204904 241538 204956 241544
rect 204916 238513 204944 241538
rect 204902 238504 204958 238513
rect 204902 238439 204958 238448
rect 205284 230081 205312 300154
rect 205270 230072 205326 230081
rect 205270 230007 205326 230016
rect 205376 228993 205404 302942
rect 205468 231849 205496 312598
rect 205548 305108 205600 305114
rect 205548 305050 205600 305056
rect 205454 231840 205510 231849
rect 205454 231775 205510 231784
rect 205362 228984 205418 228993
rect 205362 228919 205418 228928
rect 205376 228313 205404 228919
rect 205362 228304 205418 228313
rect 205362 228239 205418 228248
rect 205560 212430 205588 305050
rect 206466 304328 206522 304337
rect 206466 304263 206522 304272
rect 206480 248414 206508 304263
rect 206388 248386 206508 248414
rect 206388 240961 206416 248386
rect 206468 243636 206520 243642
rect 206468 243578 206520 243584
rect 206374 240952 206430 240961
rect 206374 240887 206430 240896
rect 206480 238754 206508 243578
rect 206572 243522 206600 318854
rect 206664 243642 206692 319262
rect 206652 243636 206704 243642
rect 206652 243578 206704 243584
rect 206572 243494 206692 243522
rect 206480 238726 206600 238754
rect 206572 233238 206600 238726
rect 206664 238241 206692 243494
rect 206650 238232 206706 238241
rect 206650 238167 206706 238176
rect 206664 237697 206692 238167
rect 206650 237688 206706 237697
rect 206650 237623 206706 237632
rect 205640 233232 205692 233238
rect 205640 233174 205692 233180
rect 206560 233232 206612 233238
rect 206560 233174 206612 233180
rect 205652 232626 205680 233174
rect 205640 232620 205692 232626
rect 205640 232562 205692 232568
rect 206756 229094 206784 321642
rect 217966 321056 218022 321065
rect 217966 320991 218022 321000
rect 206926 320920 206982 320929
rect 206926 320855 206982 320864
rect 206834 316704 206890 316713
rect 206834 316639 206890 316648
rect 206664 229066 206784 229094
rect 206664 223553 206692 229066
rect 206848 223938 206876 316639
rect 206940 224058 206968 320855
rect 210974 320784 211030 320793
rect 210974 320719 211030 320728
rect 207938 319560 207994 319569
rect 207938 319495 207994 319504
rect 207848 301504 207900 301510
rect 207848 301446 207900 301452
rect 207756 298852 207808 298858
rect 207756 298794 207808 298800
rect 207768 240854 207796 298794
rect 207756 240848 207808 240854
rect 207756 240790 207808 240796
rect 207860 239465 207888 301446
rect 207846 239456 207902 239465
rect 207846 239391 207902 239400
rect 207952 238754 207980 319495
rect 208030 319424 208086 319433
rect 208030 319359 208086 319368
rect 207860 238726 207980 238754
rect 207664 238604 207716 238610
rect 207664 238546 207716 238552
rect 206928 224052 206980 224058
rect 206928 223994 206980 224000
rect 206848 223910 206968 223938
rect 206836 223848 206888 223854
rect 206836 223790 206888 223796
rect 205638 223544 205694 223553
rect 205638 223479 205694 223488
rect 206650 223544 206706 223553
rect 206650 223479 206706 223488
rect 205652 222970 205680 223479
rect 205640 222964 205692 222970
rect 205640 222906 205692 222912
rect 205640 216640 205692 216646
rect 205640 216582 205692 216588
rect 205652 216034 205680 216582
rect 205640 216028 205692 216034
rect 205640 215970 205692 215976
rect 206848 215286 206876 223790
rect 206940 216646 206968 223910
rect 206928 216640 206980 216646
rect 206928 216582 206980 216588
rect 205640 215280 205692 215286
rect 205640 215222 205692 215228
rect 206836 215280 206888 215286
rect 206836 215222 206888 215228
rect 205652 214674 205680 215222
rect 205640 214668 205692 214674
rect 205640 214610 205692 214616
rect 205548 212424 205600 212430
rect 205548 212366 205600 212372
rect 204812 212084 204864 212090
rect 204812 212026 204864 212032
rect 204824 209916 204852 212026
rect 205560 211154 205588 212366
rect 205560 211126 205680 211154
rect 205272 210452 205324 210458
rect 205272 210394 205324 210400
rect 204312 209788 204484 209794
rect 204260 209782 204484 209788
rect 204272 209780 204484 209782
rect 204272 209766 204470 209780
rect 203156 209568 203208 209574
rect 203156 209510 203208 209516
rect 203892 209568 203944 209574
rect 203944 209516 204102 209522
rect 203892 209510 204102 209516
rect 202880 209500 202932 209506
rect 203904 209494 204102 209510
rect 202880 209442 202932 209448
rect 163596 209432 163648 209438
rect 201684 209432 201736 209438
rect 163648 209380 163990 209386
rect 163596 209374 163990 209380
rect 204996 209432 205048 209438
rect 201736 209380 201894 209386
rect 201684 209374 201894 209380
rect 205284 209386 205312 210394
rect 205364 210044 205416 210050
rect 205364 209986 205416 209992
rect 205376 209930 205404 209986
rect 205652 209930 205680 211126
rect 205376 209902 205574 209930
rect 205652 209902 205942 209930
rect 205048 209380 205312 209386
rect 204996 209374 205312 209380
rect 163608 209358 163990 209374
rect 201696 209358 201894 209374
rect 205008 209358 205312 209374
rect 207570 170368 207626 170377
rect 207570 170303 207626 170312
rect 162400 161560 162452 161566
rect 162452 161508 162532 161514
rect 162400 161502 162532 161508
rect 162412 161486 162532 161502
rect 162504 160684 162532 161486
rect 207480 161152 207532 161158
rect 207480 161094 207532 161100
rect 162596 159186 162624 160140
rect 162688 159934 162716 160140
rect 162676 159928 162728 159934
rect 162676 159870 162728 159876
rect 162584 159180 162636 159186
rect 162584 159122 162636 159128
rect 162308 158500 162360 158506
rect 162308 158442 162360 158448
rect 162216 158296 162268 158302
rect 162216 158238 162268 158244
rect 162780 158030 162808 160140
rect 162768 158024 162820 158030
rect 162768 157966 162820 157972
rect 162872 157418 162900 160140
rect 162964 159934 162992 160140
rect 162952 159928 163004 159934
rect 163056 159905 163084 160140
rect 162952 159870 163004 159876
rect 163042 159896 163098 159905
rect 163148 159866 163176 160140
rect 163042 159831 163098 159840
rect 163136 159860 163188 159866
rect 163136 159802 163188 159808
rect 162950 159760 163006 159769
rect 163240 159746 163268 160140
rect 163332 159934 163360 160140
rect 163320 159928 163372 159934
rect 163424 159905 163452 160140
rect 163320 159870 163372 159876
rect 163410 159896 163466 159905
rect 163006 159718 163268 159746
rect 162950 159695 163006 159704
rect 162964 159089 162992 159695
rect 163044 159656 163096 159662
rect 163044 159598 163096 159604
rect 162950 159080 163006 159089
rect 162950 159015 163006 159024
rect 163056 158681 163084 159598
rect 163136 158976 163188 158982
rect 163136 158918 163188 158924
rect 163042 158672 163098 158681
rect 163042 158607 163098 158616
rect 163044 158568 163096 158574
rect 163044 158510 163096 158516
rect 162860 157412 162912 157418
rect 162860 157354 162912 157360
rect 162124 157208 162176 157214
rect 162124 157150 162176 157156
rect 162860 157208 162912 157214
rect 162860 157150 162912 157156
rect 162216 157140 162268 157146
rect 162216 157082 162268 157088
rect 162124 156868 162176 156874
rect 162124 156810 162176 156816
rect 162136 156602 162164 156810
rect 162124 156596 162176 156602
rect 162124 156538 162176 156544
rect 161848 155712 161900 155718
rect 161848 155654 161900 155660
rect 162228 147674 162256 157082
rect 162136 147646 162256 147674
rect 161756 135924 161808 135930
rect 161756 135866 161808 135872
rect 162136 3602 162164 147646
rect 162872 134570 162900 157150
rect 162860 134564 162912 134570
rect 162860 134506 162912 134512
rect 162860 118040 162912 118046
rect 162860 117982 162912 117988
rect 162872 16574 162900 117982
rect 163056 117978 163084 158510
rect 163044 117972 163096 117978
rect 163044 117914 163096 117920
rect 163148 105602 163176 158918
rect 163332 157334 163360 159870
rect 163410 159831 163466 159840
rect 163516 159746 163544 160140
rect 163608 159905 163636 160140
rect 163594 159896 163650 159905
rect 163594 159831 163650 159840
rect 163424 159718 163544 159746
rect 163424 159633 163452 159718
rect 163410 159624 163466 159633
rect 163410 159559 163466 159568
rect 163424 158982 163452 159559
rect 163412 158976 163464 158982
rect 163412 158918 163464 158924
rect 163504 158024 163556 158030
rect 163502 157992 163504 158001
rect 163556 157992 163558 158001
rect 163502 157927 163558 157936
rect 163504 157480 163556 157486
rect 163502 157448 163504 157457
rect 163556 157448 163558 157457
rect 163502 157383 163558 157392
rect 163332 157306 163452 157334
rect 163228 155712 163280 155718
rect 163228 155654 163280 155660
rect 163240 152538 163268 155654
rect 163240 152510 163360 152538
rect 163228 152448 163280 152454
rect 163228 152390 163280 152396
rect 163240 119406 163268 152390
rect 163332 147674 163360 152510
rect 163424 148374 163452 157306
rect 163502 156496 163558 156505
rect 163502 156431 163504 156440
rect 163556 156431 163558 156440
rect 163504 156402 163556 156408
rect 163412 148368 163464 148374
rect 163412 148310 163464 148316
rect 163332 147646 163452 147674
rect 163228 119400 163280 119406
rect 163228 119342 163280 119348
rect 163424 112470 163452 147646
rect 163516 140078 163544 156402
rect 163608 147674 163636 159831
rect 163700 159662 163728 160140
rect 163688 159656 163740 159662
rect 163688 159598 163740 159604
rect 163792 158642 163820 160140
rect 163780 158636 163832 158642
rect 163780 158578 163832 158584
rect 163686 157856 163742 157865
rect 163686 157791 163742 157800
rect 163700 157554 163728 157791
rect 163688 157548 163740 157554
rect 163688 157490 163740 157496
rect 163792 152454 163820 158578
rect 163884 158545 163912 160140
rect 163870 158536 163926 158545
rect 163870 158471 163926 158480
rect 163976 158409 164004 160140
rect 163962 158400 164018 158409
rect 163962 158335 164018 158344
rect 163976 158166 164004 158335
rect 163964 158160 164016 158166
rect 163964 158102 164016 158108
rect 164068 157185 164096 160140
rect 164160 159866 164188 160140
rect 164252 159905 164280 160140
rect 164238 159896 164294 159905
rect 164148 159860 164200 159866
rect 164238 159831 164294 159840
rect 164148 159802 164200 159808
rect 164160 158778 164188 159802
rect 164240 159316 164292 159322
rect 164240 159258 164292 159264
rect 164148 158772 164200 158778
rect 164148 158714 164200 158720
rect 164252 158409 164280 159258
rect 164344 158982 164372 160140
rect 164436 159866 164464 160140
rect 164424 159860 164476 159866
rect 164424 159802 164476 159808
rect 164424 159588 164476 159594
rect 164424 159530 164476 159536
rect 164436 159254 164464 159530
rect 164424 159248 164476 159254
rect 164424 159190 164476 159196
rect 164332 158976 164384 158982
rect 164332 158918 164384 158924
rect 164330 158808 164386 158817
rect 164330 158743 164386 158752
rect 164424 158772 164476 158778
rect 164344 158710 164372 158743
rect 164424 158714 164476 158720
rect 164332 158704 164384 158710
rect 164332 158646 164384 158652
rect 164332 158568 164384 158574
rect 164332 158510 164384 158516
rect 164238 158400 164294 158409
rect 164344 158370 164372 158510
rect 164238 158335 164294 158344
rect 164332 158364 164384 158370
rect 164332 158306 164384 158312
rect 164344 158273 164372 158306
rect 164330 158264 164386 158273
rect 164330 158199 164386 158208
rect 164240 157888 164292 157894
rect 164240 157830 164292 157836
rect 164330 157856 164386 157865
rect 164146 157448 164202 157457
rect 164252 157418 164280 157830
rect 164330 157791 164386 157800
rect 164146 157383 164148 157392
rect 164200 157383 164202 157392
rect 164240 157412 164292 157418
rect 164148 157354 164200 157360
rect 164240 157354 164292 157360
rect 164054 157176 164110 157185
rect 164054 157111 164110 157120
rect 164240 156256 164292 156262
rect 164240 156198 164292 156204
rect 163780 152448 163832 152454
rect 163780 152390 163832 152396
rect 163608 147646 163820 147674
rect 163504 140072 163556 140078
rect 163504 140014 163556 140020
rect 163412 112464 163464 112470
rect 163412 112406 163464 112412
rect 163136 105596 163188 105602
rect 163136 105538 163188 105544
rect 162872 16546 163728 16574
rect 162124 3596 162176 3602
rect 162124 3538 162176 3544
rect 162492 3324 162544 3330
rect 162492 3266 162544 3272
rect 161480 3256 161532 3262
rect 161480 3198 161532 3204
rect 162504 480 162532 3266
rect 163700 480 163728 16546
rect 163792 11762 163820 147646
rect 164252 142866 164280 156198
rect 164344 155310 164372 157791
rect 164332 155304 164384 155310
rect 164332 155246 164384 155252
rect 164240 142860 164292 142866
rect 164240 142802 164292 142808
rect 164436 137290 164464 158714
rect 164528 143342 164556 160140
rect 164620 158642 164648 160140
rect 164712 159939 164740 160140
rect 164698 159930 164754 159939
rect 164698 159865 164754 159874
rect 164700 159792 164752 159798
rect 164700 159734 164752 159740
rect 164712 158778 164740 159734
rect 164700 158772 164752 158778
rect 164700 158714 164752 158720
rect 164698 158672 164754 158681
rect 164608 158636 164660 158642
rect 164698 158607 164754 158616
rect 164608 158578 164660 158584
rect 164606 158536 164662 158545
rect 164606 158471 164662 158480
rect 164620 158001 164648 158471
rect 164606 157992 164662 158001
rect 164606 157927 164662 157936
rect 164516 143336 164568 143342
rect 164516 143278 164568 143284
rect 164528 141438 164556 143278
rect 164516 141432 164568 141438
rect 164516 141374 164568 141380
rect 164424 137284 164476 137290
rect 164424 137226 164476 137232
rect 164620 102814 164648 157927
rect 164712 116618 164740 158607
rect 164804 157321 164832 160140
rect 164896 158545 164924 160140
rect 164882 158536 164938 158545
rect 164882 158471 164938 158480
rect 164882 158400 164938 158409
rect 164882 158335 164938 158344
rect 164790 157312 164846 157321
rect 164790 157247 164846 157256
rect 164792 155644 164844 155650
rect 164792 155586 164844 155592
rect 164700 116612 164752 116618
rect 164700 116554 164752 116560
rect 164608 102808 164660 102814
rect 164608 102750 164660 102756
rect 163780 11756 163832 11762
rect 163780 11698 163832 11704
rect 164804 6914 164832 155586
rect 164896 147674 164924 158335
rect 164988 157282 165016 160140
rect 164976 157276 165028 157282
rect 164976 157218 165028 157224
rect 164988 156262 165016 157218
rect 164976 156256 165028 156262
rect 164976 156198 165028 156204
rect 165080 155922 165108 160140
rect 165172 159769 165200 160140
rect 165158 159760 165214 159769
rect 165158 159695 165214 159704
rect 165264 159644 165292 160140
rect 165356 159905 165384 160140
rect 165342 159896 165398 159905
rect 165342 159831 165398 159840
rect 165344 159792 165396 159798
rect 165344 159734 165396 159740
rect 165448 159746 165476 160140
rect 165540 159934 165568 160140
rect 165528 159928 165580 159934
rect 165632 159905 165660 160140
rect 165528 159870 165580 159876
rect 165618 159896 165674 159905
rect 165618 159831 165674 159840
rect 165620 159792 165672 159798
rect 165526 159760 165582 159769
rect 165172 159616 165292 159644
rect 165172 158953 165200 159616
rect 165356 159322 165384 159734
rect 165448 159718 165526 159746
rect 165344 159316 165396 159322
rect 165344 159258 165396 159264
rect 165252 158976 165304 158982
rect 165158 158944 165214 158953
rect 165252 158918 165304 158924
rect 165158 158879 165214 158888
rect 165158 158536 165214 158545
rect 165158 158471 165214 158480
rect 165172 157962 165200 158471
rect 165160 157956 165212 157962
rect 165160 157898 165212 157904
rect 165264 157865 165292 158918
rect 165344 157888 165396 157894
rect 165250 157856 165306 157865
rect 165344 157830 165396 157836
rect 165250 157791 165306 157800
rect 165068 155916 165120 155922
rect 165068 155858 165120 155864
rect 164896 147646 165200 147674
rect 164884 147008 164936 147014
rect 164884 146950 164936 146956
rect 164896 13122 164924 146950
rect 165172 140146 165200 147646
rect 165264 147014 165292 157791
rect 165356 157690 165384 157830
rect 165344 157684 165396 157690
rect 165344 157626 165396 157632
rect 165252 147008 165304 147014
rect 165252 146950 165304 146956
rect 165160 140140 165212 140146
rect 165160 140082 165212 140088
rect 165448 17270 165476 159718
rect 165620 159734 165672 159740
rect 165526 159695 165582 159704
rect 165632 159633 165660 159734
rect 165618 159624 165674 159633
rect 165618 159559 165674 159568
rect 165528 159452 165580 159458
rect 165528 159394 165580 159400
rect 165540 158642 165568 159394
rect 165632 158953 165660 159559
rect 165618 158944 165674 158953
rect 165618 158879 165674 158888
rect 165724 158794 165752 160140
rect 165632 158766 165752 158794
rect 165528 158636 165580 158642
rect 165528 158578 165580 158584
rect 165632 158438 165660 158766
rect 165710 158672 165766 158681
rect 165710 158607 165766 158616
rect 165620 158432 165672 158438
rect 165620 158374 165672 158380
rect 165620 152244 165672 152250
rect 165620 152186 165672 152192
rect 165632 109750 165660 152186
rect 165724 142934 165752 158607
rect 165816 157334 165844 160140
rect 165908 159089 165936 160140
rect 165894 159080 165950 159089
rect 165894 159015 165950 159024
rect 166000 158930 166028 160140
rect 165908 158902 166028 158930
rect 165908 158370 165936 158902
rect 166092 158794 166120 160140
rect 166184 159866 166212 160140
rect 166276 159905 166304 160140
rect 166262 159896 166318 159905
rect 166172 159860 166224 159866
rect 166262 159831 166318 159840
rect 166172 159802 166224 159808
rect 166170 159760 166226 159769
rect 166170 159695 166226 159704
rect 166000 158766 166120 158794
rect 165896 158364 165948 158370
rect 165896 158306 165948 158312
rect 165816 157306 165936 157334
rect 165804 152516 165856 152522
rect 165804 152458 165856 152464
rect 165712 142928 165764 142934
rect 165712 142870 165764 142876
rect 165816 138718 165844 152458
rect 165908 147014 165936 157306
rect 166000 157049 166028 158766
rect 166184 158658 166212 159695
rect 166276 158681 166304 159831
rect 166368 159633 166396 160140
rect 166354 159624 166410 159633
rect 166354 159559 166410 159568
rect 166460 159225 166488 160140
rect 166552 159254 166580 160140
rect 166540 159248 166592 159254
rect 166446 159216 166502 159225
rect 166540 159190 166592 159196
rect 166446 159151 166502 159160
rect 166354 158944 166410 158953
rect 166354 158879 166410 158888
rect 166092 158630 166212 158658
rect 166262 158672 166318 158681
rect 165986 157040 166042 157049
rect 165986 156975 166042 156984
rect 165896 147008 165948 147014
rect 165896 146950 165948 146956
rect 165804 138712 165856 138718
rect 165804 138654 165856 138660
rect 166092 124914 166120 158630
rect 166262 158607 166318 158616
rect 166368 158522 166396 158879
rect 166184 158494 166396 158522
rect 166184 133210 166212 158494
rect 166356 158364 166408 158370
rect 166356 158306 166408 158312
rect 166262 158128 166318 158137
rect 166262 158063 166318 158072
rect 166276 157593 166304 158063
rect 166262 157584 166318 157593
rect 166368 157554 166396 158306
rect 166262 157519 166318 157528
rect 166356 157548 166408 157554
rect 166356 157490 166408 157496
rect 166368 155990 166396 157490
rect 166356 155984 166408 155990
rect 166356 155926 166408 155932
rect 166460 152522 166488 159151
rect 166448 152516 166500 152522
rect 166448 152458 166500 152464
rect 166552 152250 166580 159190
rect 166644 155786 166672 160140
rect 166736 159905 166764 160140
rect 166722 159896 166778 159905
rect 166722 159831 166778 159840
rect 166736 158545 166764 159831
rect 166828 159769 166856 160140
rect 166814 159760 166870 159769
rect 166814 159695 166870 159704
rect 166920 159610 166948 160140
rect 166828 159582 166948 159610
rect 166828 158778 166856 159582
rect 166908 159452 166960 159458
rect 166908 159394 166960 159400
rect 166816 158772 166868 158778
rect 166816 158714 166868 158720
rect 166814 158672 166870 158681
rect 166814 158607 166870 158616
rect 166722 158536 166778 158545
rect 166722 158471 166778 158480
rect 166724 158296 166776 158302
rect 166724 158238 166776 158244
rect 166736 157486 166764 158238
rect 166724 157480 166776 157486
rect 166724 157422 166776 157428
rect 166632 155780 166684 155786
rect 166632 155722 166684 155728
rect 166540 152244 166592 152250
rect 166540 152186 166592 152192
rect 166264 147008 166316 147014
rect 166264 146950 166316 146956
rect 166276 141506 166304 146950
rect 166264 141500 166316 141506
rect 166264 141442 166316 141448
rect 166172 133204 166224 133210
rect 166172 133146 166224 133152
rect 166264 133204 166316 133210
rect 166264 133146 166316 133152
rect 166080 124908 166132 124914
rect 166080 124850 166132 124856
rect 165620 109744 165672 109750
rect 165620 109686 165672 109692
rect 165436 17264 165488 17270
rect 165436 17206 165488 17212
rect 164884 13116 164936 13122
rect 164884 13058 164936 13064
rect 164804 6886 164924 6914
rect 164896 480 164924 6886
rect 166080 3460 166132 3466
rect 166080 3402 166132 3408
rect 166092 480 166120 3402
rect 166276 3330 166304 133146
rect 166828 115258 166856 158607
rect 166920 158234 166948 159394
rect 166908 158228 166960 158234
rect 166908 158170 166960 158176
rect 167012 157729 167040 160140
rect 167104 158681 167132 160140
rect 167196 159905 167224 160140
rect 167182 159896 167238 159905
rect 167182 159831 167238 159840
rect 167196 159458 167224 159831
rect 167184 159452 167236 159458
rect 167184 159394 167236 159400
rect 167182 159352 167238 159361
rect 167182 159287 167238 159296
rect 167196 158982 167224 159287
rect 167184 158976 167236 158982
rect 167184 158918 167236 158924
rect 167090 158672 167146 158681
rect 167090 158607 167146 158616
rect 166998 157720 167054 157729
rect 166998 157655 167054 157664
rect 167104 120766 167132 158607
rect 167184 156120 167236 156126
rect 167184 156062 167236 156068
rect 167196 151814 167224 156062
rect 167288 155972 167316 160140
rect 167380 159712 167408 160140
rect 167472 159905 167500 160140
rect 167458 159896 167514 159905
rect 167458 159831 167514 159840
rect 167564 159798 167592 160140
rect 167656 159905 167684 160140
rect 167748 159934 167776 160140
rect 167736 159928 167788 159934
rect 167642 159896 167698 159905
rect 167736 159870 167788 159876
rect 167642 159831 167698 159840
rect 167552 159792 167604 159798
rect 167552 159734 167604 159740
rect 167460 159724 167512 159730
rect 167380 159684 167460 159712
rect 167460 159666 167512 159672
rect 167368 159316 167420 159322
rect 167368 159258 167420 159264
rect 167380 158438 167408 159258
rect 167368 158432 167420 158438
rect 167368 158374 167420 158380
rect 167458 158400 167514 158409
rect 167458 158335 167514 158344
rect 167288 155944 167408 155972
rect 167196 151786 167316 151814
rect 167288 140622 167316 151786
rect 167276 140616 167328 140622
rect 167276 140558 167328 140564
rect 167288 139466 167316 140558
rect 167380 140486 167408 155944
rect 167368 140480 167420 140486
rect 167368 140422 167420 140428
rect 167276 139460 167328 139466
rect 167276 139402 167328 139408
rect 167380 138786 167408 140422
rect 167368 138780 167420 138786
rect 167368 138722 167420 138728
rect 167092 120760 167144 120766
rect 167092 120702 167144 120708
rect 166816 115252 166868 115258
rect 166816 115194 166868 115200
rect 167472 108322 167500 158335
rect 167564 154834 167592 159734
rect 167656 157010 167684 159831
rect 167736 159724 167788 159730
rect 167736 159666 167788 159672
rect 167748 159322 167776 159666
rect 167736 159316 167788 159322
rect 167736 159258 167788 159264
rect 167644 157004 167696 157010
rect 167644 156946 167696 156952
rect 167552 154828 167604 154834
rect 167552 154770 167604 154776
rect 167748 154574 167776 159258
rect 167840 155972 167868 160140
rect 167932 159633 167960 160140
rect 167918 159624 167974 159633
rect 167918 159559 167974 159568
rect 168024 156641 168052 160140
rect 168010 156632 168066 156641
rect 168010 156567 168066 156576
rect 168116 156126 168144 160140
rect 168208 159769 168236 160140
rect 168300 159905 168328 160140
rect 168286 159896 168342 159905
rect 168286 159831 168342 159840
rect 168194 159760 168250 159769
rect 168194 159695 168250 159704
rect 168208 156670 168236 159695
rect 168392 159610 168420 160140
rect 168484 159769 168512 160140
rect 168470 159760 168526 159769
rect 168470 159695 168526 159704
rect 168288 159588 168340 159594
rect 168392 159582 168512 159610
rect 168288 159530 168340 159536
rect 168300 158506 168328 159530
rect 168288 158500 168340 158506
rect 168288 158442 168340 158448
rect 168378 158400 168434 158409
rect 168378 158335 168434 158344
rect 168286 158264 168342 158273
rect 168286 158199 168288 158208
rect 168340 158199 168342 158208
rect 168288 158170 168340 158176
rect 168196 156664 168248 156670
rect 168196 156606 168248 156612
rect 168104 156120 168156 156126
rect 168104 156062 168156 156068
rect 167840 155944 168144 155972
rect 167564 154546 167776 154574
rect 167564 151814 167592 154546
rect 167564 151786 167960 151814
rect 167644 139460 167696 139466
rect 167644 139402 167696 139408
rect 167460 108316 167512 108322
rect 167460 108258 167512 108264
rect 167656 7614 167684 139402
rect 167736 138032 167788 138038
rect 167736 137974 167788 137980
rect 167748 127634 167776 137974
rect 167736 127628 167788 127634
rect 167736 127570 167788 127576
rect 167644 7608 167696 7614
rect 167644 7550 167696 7556
rect 167932 4826 167960 151786
rect 168116 139194 168144 155944
rect 168288 154828 168340 154834
rect 168288 154770 168340 154776
rect 168104 139188 168156 139194
rect 168104 139130 168156 139136
rect 168116 138038 168144 139130
rect 168104 138032 168156 138038
rect 168104 137974 168156 137980
rect 168300 129062 168328 154770
rect 168392 134638 168420 158335
rect 168484 158273 168512 159582
rect 168576 159050 168604 160140
rect 168564 159044 168616 159050
rect 168564 158986 168616 158992
rect 168562 158944 168618 158953
rect 168562 158879 168618 158888
rect 168470 158264 168526 158273
rect 168470 158199 168526 158208
rect 168470 158128 168526 158137
rect 168470 158063 168526 158072
rect 168484 157729 168512 158063
rect 168470 157720 168526 157729
rect 168470 157655 168526 157664
rect 168576 157570 168604 158879
rect 168668 158681 168696 160140
rect 168760 159905 168788 160140
rect 168746 159896 168802 159905
rect 168746 159831 168802 159840
rect 168654 158672 168710 158681
rect 168654 158607 168710 158616
rect 168484 157542 168604 157570
rect 168484 155718 168512 157542
rect 168760 156738 168788 159831
rect 168852 156777 168880 160140
rect 168944 159118 168972 160140
rect 169036 159769 169064 160140
rect 169022 159760 169078 159769
rect 169022 159695 169078 159704
rect 168932 159112 168984 159118
rect 168932 159054 168984 159060
rect 168944 158137 168972 159054
rect 168930 158128 168986 158137
rect 168930 158063 168986 158072
rect 168932 157956 168984 157962
rect 168932 157898 168984 157904
rect 168838 156768 168894 156777
rect 168748 156732 168800 156738
rect 168838 156703 168894 156712
rect 168748 156674 168800 156680
rect 168656 155984 168708 155990
rect 168656 155926 168708 155932
rect 168472 155712 168524 155718
rect 168472 155654 168524 155660
rect 168668 145586 168696 155926
rect 168656 145580 168708 145586
rect 168656 145522 168708 145528
rect 168380 134632 168432 134638
rect 168380 134574 168432 134580
rect 168288 129056 168340 129062
rect 168288 128998 168340 129004
rect 168944 14482 168972 157898
rect 169036 156806 169064 159695
rect 169024 156800 169076 156806
rect 169024 156742 169076 156748
rect 169128 155990 169156 160140
rect 169220 159905 169248 160140
rect 169206 159896 169262 159905
rect 169206 159831 169262 159840
rect 169312 159633 169340 160140
rect 169298 159624 169354 159633
rect 169298 159559 169354 159568
rect 169208 158636 169260 158642
rect 169208 158578 169260 158584
rect 169116 155984 169168 155990
rect 169116 155926 169168 155932
rect 169220 155802 169248 158578
rect 169312 157962 169340 159559
rect 169404 159497 169432 160140
rect 169496 159905 169524 160140
rect 169482 159896 169538 159905
rect 169482 159831 169538 159840
rect 169390 159488 169446 159497
rect 169390 159423 169446 159432
rect 169390 158672 169446 158681
rect 169390 158607 169446 158616
rect 169300 157956 169352 157962
rect 169300 157898 169352 157904
rect 169300 155916 169352 155922
rect 169300 155858 169352 155864
rect 169128 155774 169248 155802
rect 169128 144294 169156 155774
rect 169208 155712 169260 155718
rect 169208 155654 169260 155660
rect 169116 144288 169168 144294
rect 169116 144230 169168 144236
rect 169024 130416 169076 130422
rect 169024 130358 169076 130364
rect 168932 14476 168984 14482
rect 168932 14418 168984 14424
rect 167920 4820 167972 4826
rect 167920 4762 167972 4768
rect 168380 3528 168432 3534
rect 168380 3470 168432 3476
rect 166264 3324 166316 3330
rect 166264 3266 166316 3272
rect 167184 3052 167236 3058
rect 167184 2994 167236 3000
rect 167196 480 167224 2994
rect 168392 480 168420 3470
rect 169036 3058 169064 130358
rect 169220 106962 169248 155654
rect 169312 146266 169340 155858
rect 169404 151814 169432 158607
rect 169496 158409 169524 159831
rect 169588 159458 169616 160140
rect 169576 159452 169628 159458
rect 169576 159394 169628 159400
rect 169482 158400 169538 158409
rect 169482 158335 169538 158344
rect 169484 157956 169536 157962
rect 169484 157898 169536 157904
rect 169496 157418 169524 157898
rect 169484 157412 169536 157418
rect 169484 157354 169536 157360
rect 169588 153950 169616 159394
rect 169680 155922 169708 160140
rect 169772 159934 169800 160140
rect 169760 159928 169812 159934
rect 169760 159870 169812 159876
rect 169772 158642 169800 159870
rect 169864 159497 169892 160140
rect 169850 159488 169906 159497
rect 169850 159423 169906 159432
rect 169760 158636 169812 158642
rect 169760 158578 169812 158584
rect 169760 158092 169812 158098
rect 169760 158034 169812 158040
rect 169772 156602 169800 158034
rect 169760 156596 169812 156602
rect 169760 156538 169812 156544
rect 169668 155916 169720 155922
rect 169668 155858 169720 155864
rect 169576 153944 169628 153950
rect 169576 153886 169628 153892
rect 169404 151786 169524 151814
rect 169300 146260 169352 146266
rect 169300 146202 169352 146208
rect 169496 123486 169524 151786
rect 169760 143200 169812 143206
rect 169760 143142 169812 143148
rect 169772 143002 169800 143142
rect 169760 142996 169812 143002
rect 169760 142938 169812 142944
rect 169760 140344 169812 140350
rect 169760 140286 169812 140292
rect 169772 133278 169800 140286
rect 169760 133272 169812 133278
rect 169760 133214 169812 133220
rect 169484 123480 169536 123486
rect 169484 123422 169536 123428
rect 169208 106956 169260 106962
rect 169208 106898 169260 106904
rect 169864 104174 169892 159423
rect 169956 158982 169984 160140
rect 169944 158976 169996 158982
rect 169944 158918 169996 158924
rect 169944 155984 169996 155990
rect 169944 155926 169996 155932
rect 169956 140418 169984 155926
rect 169944 140412 169996 140418
rect 169944 140354 169996 140360
rect 170048 140350 170076 160140
rect 170140 158098 170168 160140
rect 170128 158092 170180 158098
rect 170128 158034 170180 158040
rect 170232 157622 170260 160140
rect 170220 157616 170272 157622
rect 170220 157558 170272 157564
rect 170126 157312 170182 157321
rect 170126 157247 170182 157256
rect 170140 143206 170168 157247
rect 170324 155990 170352 160140
rect 170416 159905 170444 160140
rect 170402 159896 170458 159905
rect 170402 159831 170458 159840
rect 170312 155984 170364 155990
rect 170312 155926 170364 155932
rect 170416 155530 170444 159831
rect 170508 158273 170536 160140
rect 170600 159769 170628 160140
rect 170586 159760 170642 159769
rect 170692 159730 170720 160140
rect 170784 159769 170812 160140
rect 170770 159760 170826 159769
rect 170586 159695 170642 159704
rect 170680 159724 170732 159730
rect 170770 159695 170826 159704
rect 170680 159666 170732 159672
rect 170680 159588 170732 159594
rect 170680 159530 170732 159536
rect 170586 158944 170642 158953
rect 170586 158879 170642 158888
rect 170600 158438 170628 158879
rect 170588 158432 170640 158438
rect 170588 158374 170640 158380
rect 170494 158264 170550 158273
rect 170494 158199 170550 158208
rect 170692 158137 170720 159530
rect 170772 159044 170824 159050
rect 170876 159032 170904 160140
rect 170968 159905 170996 160140
rect 170954 159896 171010 159905
rect 170954 159831 171010 159840
rect 170956 159792 171008 159798
rect 170954 159760 170956 159769
rect 171008 159760 171010 159769
rect 170954 159695 171010 159704
rect 171060 159186 171088 160140
rect 171152 159905 171180 160140
rect 171138 159896 171194 159905
rect 171138 159831 171194 159840
rect 171048 159180 171100 159186
rect 171048 159122 171100 159128
rect 170824 159004 170904 159032
rect 170772 158986 170824 158992
rect 170678 158128 170734 158137
rect 170678 158063 170734 158072
rect 170692 156942 170720 158063
rect 170784 157593 170812 158986
rect 171060 158681 171088 159122
rect 171046 158672 171102 158681
rect 171046 158607 171102 158616
rect 170862 158264 170918 158273
rect 170862 158199 170918 158208
rect 170770 157584 170826 157593
rect 170770 157519 170826 157528
rect 170680 156936 170732 156942
rect 170680 156878 170732 156884
rect 170416 155502 170812 155530
rect 170128 143200 170180 143206
rect 170128 143142 170180 143148
rect 170404 140412 170456 140418
rect 170404 140354 170456 140360
rect 170036 140344 170088 140350
rect 170036 140286 170088 140292
rect 170416 124982 170444 140354
rect 170404 124976 170456 124982
rect 170404 124918 170456 124924
rect 169852 104168 169904 104174
rect 169852 104110 169904 104116
rect 170784 8974 170812 155502
rect 170876 152590 170904 158199
rect 170954 158128 171010 158137
rect 170954 158063 171010 158072
rect 170864 152584 170916 152590
rect 170864 152526 170916 152532
rect 170968 142154 170996 158063
rect 171152 156670 171180 159831
rect 171244 159730 171272 160140
rect 171232 159724 171284 159730
rect 171232 159666 171284 159672
rect 171230 159624 171286 159633
rect 171230 159559 171286 159568
rect 171244 158166 171272 159559
rect 171336 158681 171364 160140
rect 171428 159769 171456 160140
rect 171414 159760 171470 159769
rect 171414 159695 171470 159704
rect 171322 158672 171378 158681
rect 171322 158607 171378 158616
rect 171232 158160 171284 158166
rect 171232 158102 171284 158108
rect 171140 156664 171192 156670
rect 171140 156606 171192 156612
rect 171232 155984 171284 155990
rect 171232 155926 171284 155932
rect 171140 155712 171192 155718
rect 171140 155654 171192 155660
rect 170876 142126 170996 142154
rect 170876 131782 170904 142126
rect 170864 131776 170916 131782
rect 170864 131718 170916 131724
rect 171152 16574 171180 155654
rect 171244 141914 171272 155926
rect 171428 142154 171456 159695
rect 171520 159633 171548 160140
rect 171506 159624 171562 159633
rect 171506 159559 171562 159568
rect 171508 158976 171560 158982
rect 171508 158918 171560 158924
rect 171520 158284 171548 158918
rect 171612 158409 171640 160140
rect 171704 159594 171732 160140
rect 171796 159905 171824 160140
rect 171782 159896 171838 159905
rect 171782 159831 171838 159840
rect 171784 159724 171836 159730
rect 171784 159666 171836 159672
rect 171692 159588 171744 159594
rect 171692 159530 171744 159536
rect 171598 158400 171654 158409
rect 171704 158370 171732 159530
rect 171598 158335 171654 158344
rect 171692 158364 171744 158370
rect 171692 158306 171744 158312
rect 171520 158256 171640 158284
rect 171508 158160 171560 158166
rect 171508 158102 171560 158108
rect 171520 156754 171548 158102
rect 171612 157146 171640 158256
rect 171796 157486 171824 159666
rect 171784 157480 171836 157486
rect 171784 157422 171836 157428
rect 171600 157140 171652 157146
rect 171600 157082 171652 157088
rect 171520 156726 171640 156754
rect 171508 156664 171560 156670
rect 171508 156606 171560 156612
rect 171336 142126 171456 142154
rect 171232 141908 171284 141914
rect 171232 141850 171284 141856
rect 171336 138854 171364 142126
rect 171324 138848 171376 138854
rect 171324 138790 171376 138796
rect 171520 98666 171548 156606
rect 171612 151814 171640 156726
rect 171796 155802 171824 157422
rect 171888 155990 171916 160140
rect 171980 158137 172008 160140
rect 172072 158982 172100 160140
rect 172060 158976 172112 158982
rect 172060 158918 172112 158924
rect 172164 158778 172192 160140
rect 172152 158772 172204 158778
rect 172152 158714 172204 158720
rect 172150 158672 172206 158681
rect 172150 158607 172206 158616
rect 172060 158364 172112 158370
rect 172060 158306 172112 158312
rect 171966 158128 172022 158137
rect 171966 158063 172022 158072
rect 171876 155984 171928 155990
rect 171876 155926 171928 155932
rect 171796 155774 171916 155802
rect 171612 151786 171824 151814
rect 171796 129130 171824 151786
rect 171888 140214 171916 155774
rect 171980 148510 172008 158063
rect 171968 148504 172020 148510
rect 171968 148446 172020 148452
rect 172072 145722 172100 158306
rect 172164 151814 172192 158607
rect 172256 153105 172284 160140
rect 172348 158302 172376 160140
rect 172336 158296 172388 158302
rect 172336 158238 172388 158244
rect 172440 158234 172468 160140
rect 172532 159633 172560 160140
rect 172624 159905 172652 160140
rect 172610 159896 172666 159905
rect 172716 159866 172744 160140
rect 172610 159831 172666 159840
rect 172704 159860 172756 159866
rect 172704 159802 172756 159808
rect 172702 159760 172758 159769
rect 172702 159695 172758 159704
rect 172518 159624 172574 159633
rect 172518 159559 172574 159568
rect 172612 159384 172664 159390
rect 172612 159326 172664 159332
rect 172624 159066 172652 159326
rect 172532 159038 172652 159066
rect 172428 158228 172480 158234
rect 172428 158170 172480 158176
rect 172532 154018 172560 159038
rect 172716 158522 172744 159695
rect 172808 158710 172836 160140
rect 172900 159905 172928 160140
rect 172886 159896 172942 159905
rect 172886 159831 172942 159840
rect 172888 159792 172940 159798
rect 172888 159734 172940 159740
rect 172796 158704 172848 158710
rect 172796 158646 172848 158652
rect 172716 158494 172836 158522
rect 172612 158432 172664 158438
rect 172612 158374 172664 158380
rect 172624 158098 172652 158374
rect 172702 158264 172758 158273
rect 172702 158199 172758 158208
rect 172612 158092 172664 158098
rect 172612 158034 172664 158040
rect 172520 154012 172572 154018
rect 172520 153954 172572 153960
rect 172612 153196 172664 153202
rect 172612 153138 172664 153144
rect 172242 153096 172298 153105
rect 172242 153031 172298 153040
rect 172164 151786 172468 151814
rect 172060 145716 172112 145722
rect 172060 145658 172112 145664
rect 171876 140208 171928 140214
rect 171876 140150 171928 140156
rect 171784 129124 171836 129130
rect 171784 129066 171836 129072
rect 172440 127702 172468 151786
rect 172624 142154 172652 153138
rect 172716 151094 172744 158199
rect 172808 151814 172836 158494
rect 172900 156330 172928 159734
rect 172992 158574 173020 160140
rect 173084 158681 173112 160140
rect 173176 159390 173204 160140
rect 173268 159769 173296 160140
rect 173254 159760 173310 159769
rect 173254 159695 173310 159704
rect 173256 159656 173308 159662
rect 173256 159598 173308 159604
rect 173268 159458 173296 159598
rect 173256 159452 173308 159458
rect 173256 159394 173308 159400
rect 173164 159384 173216 159390
rect 173164 159326 173216 159332
rect 173070 158672 173126 158681
rect 173070 158607 173126 158616
rect 172980 158568 173032 158574
rect 172980 158510 173032 158516
rect 172992 157214 173020 158510
rect 173360 157321 173388 160140
rect 173452 159769 173480 160140
rect 173438 159760 173494 159769
rect 173438 159695 173494 159704
rect 173438 159624 173494 159633
rect 173438 159559 173494 159568
rect 173452 158953 173480 159559
rect 173438 158944 173494 158953
rect 173438 158879 173494 158888
rect 173440 158704 173492 158710
rect 173440 158646 173492 158652
rect 173346 157312 173402 157321
rect 173346 157247 173402 157256
rect 172980 157208 173032 157214
rect 172980 157150 173032 157156
rect 172888 156324 172940 156330
rect 172888 156266 172940 156272
rect 173348 155576 173400 155582
rect 173348 155518 173400 155524
rect 173256 152380 173308 152386
rect 173256 152322 173308 152328
rect 172808 151786 173112 151814
rect 172704 151088 172756 151094
rect 172704 151030 172756 151036
rect 172532 142126 172652 142154
rect 172428 127696 172480 127702
rect 172428 127638 172480 127644
rect 171508 98660 171560 98666
rect 171508 98602 171560 98608
rect 172532 16574 172560 142126
rect 173084 111110 173112 151786
rect 173162 149152 173218 149161
rect 173162 149087 173218 149096
rect 173072 111104 173124 111110
rect 173072 111046 173124 111052
rect 171152 16546 172008 16574
rect 172532 16546 172744 16574
rect 170772 8968 170824 8974
rect 170772 8910 170824 8916
rect 170772 3664 170824 3670
rect 170772 3606 170824 3612
rect 169576 3596 169628 3602
rect 169576 3538 169628 3544
rect 169024 3052 169076 3058
rect 169024 2994 169076 3000
rect 169588 480 169616 3538
rect 170784 480 170812 3606
rect 171980 480 172008 16546
rect 156574 354 156686 480
rect 156156 326 156686 354
rect 156574 -960 156686 326
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 172716 354 172744 16546
rect 173176 3466 173204 149087
rect 173268 137358 173296 152322
rect 173360 143070 173388 155518
rect 173452 154290 173480 158646
rect 173544 155582 173572 160140
rect 173532 155576 173584 155582
rect 173532 155518 173584 155524
rect 173440 154284 173492 154290
rect 173440 154226 173492 154232
rect 173636 147286 173664 160140
rect 173728 159905 173756 160140
rect 173714 159896 173770 159905
rect 173714 159831 173770 159840
rect 173728 155378 173756 159831
rect 173716 155372 173768 155378
rect 173716 155314 173768 155320
rect 173716 154284 173768 154290
rect 173716 154226 173768 154232
rect 173728 152658 173756 154226
rect 173716 152652 173768 152658
rect 173716 152594 173768 152600
rect 173820 152386 173848 160140
rect 173912 159798 173940 160140
rect 174004 159905 174032 160140
rect 173990 159896 174046 159905
rect 174096 159866 174124 160140
rect 173990 159831 174046 159840
rect 174084 159860 174136 159866
rect 173900 159792 173952 159798
rect 173900 159734 173952 159740
rect 174004 159746 174032 159831
rect 174084 159802 174136 159808
rect 174004 159718 174124 159746
rect 173992 159656 174044 159662
rect 173898 159624 173954 159633
rect 173992 159598 174044 159604
rect 173898 159559 173954 159568
rect 173808 152380 173860 152386
rect 173808 152322 173860 152328
rect 173912 148578 173940 159559
rect 174004 158409 174032 159598
rect 173990 158400 174046 158409
rect 173990 158335 174046 158344
rect 173990 158264 174046 158273
rect 173990 158199 174046 158208
rect 173900 148572 173952 148578
rect 173900 148514 173952 148520
rect 173900 147688 173952 147694
rect 173900 147630 173952 147636
rect 173624 147280 173676 147286
rect 173624 147222 173676 147228
rect 173348 143064 173400 143070
rect 173348 143006 173400 143012
rect 173256 137352 173308 137358
rect 173256 137294 173308 137300
rect 173164 3460 173216 3466
rect 173164 3402 173216 3408
rect 173134 354 173246 480
rect 172716 326 173246 354
rect 173912 354 173940 147630
rect 174004 118046 174032 158199
rect 174096 151162 174124 159718
rect 174084 151156 174136 151162
rect 174084 151098 174136 151104
rect 174188 149122 174216 160140
rect 174280 159769 174308 160140
rect 174266 159760 174322 159769
rect 174266 159695 174322 159704
rect 174268 159656 174320 159662
rect 174268 159598 174320 159604
rect 174280 158030 174308 159598
rect 174268 158024 174320 158030
rect 174268 157966 174320 157972
rect 174372 157078 174400 160140
rect 174464 157729 174492 160140
rect 174556 159905 174584 160140
rect 174542 159896 174598 159905
rect 174542 159831 174598 159840
rect 174450 157720 174506 157729
rect 174450 157655 174506 157664
rect 174360 157072 174412 157078
rect 174360 157014 174412 157020
rect 174372 155446 174400 157014
rect 174360 155440 174412 155446
rect 174360 155382 174412 155388
rect 174556 155242 174584 159831
rect 174648 158681 174676 160140
rect 174740 159089 174768 160140
rect 174832 159866 174860 160140
rect 174820 159860 174872 159866
rect 174820 159802 174872 159808
rect 174818 159760 174874 159769
rect 174818 159695 174874 159704
rect 174726 159080 174782 159089
rect 174726 159015 174782 159024
rect 174832 158817 174860 159695
rect 174818 158808 174874 158817
rect 174818 158743 174874 158752
rect 174634 158672 174690 158681
rect 174634 158607 174690 158616
rect 174636 158364 174688 158370
rect 174636 158306 174688 158312
rect 174544 155236 174596 155242
rect 174544 155178 174596 155184
rect 174648 152726 174676 158306
rect 174924 156398 174952 160140
rect 174912 156392 174964 156398
rect 174912 156334 174964 156340
rect 175016 154086 175044 160140
rect 175108 159633 175136 160140
rect 175094 159624 175150 159633
rect 175094 159559 175150 159568
rect 175096 159520 175148 159526
rect 175096 159462 175148 159468
rect 175108 158982 175136 159462
rect 175096 158976 175148 158982
rect 175096 158918 175148 158924
rect 175200 155650 175228 160140
rect 175292 158409 175320 160140
rect 175278 158400 175334 158409
rect 175278 158335 175334 158344
rect 175278 158264 175334 158273
rect 175278 158199 175334 158208
rect 175188 155644 175240 155650
rect 175188 155586 175240 155592
rect 175004 154080 175056 154086
rect 175004 154022 175056 154028
rect 174636 152720 174688 152726
rect 174636 152662 174688 152668
rect 174648 151814 174676 152662
rect 174556 151786 174676 151814
rect 174176 149116 174228 149122
rect 174176 149058 174228 149064
rect 174188 148306 174216 149058
rect 174176 148300 174228 148306
rect 174176 148242 174228 148248
rect 173992 118040 174044 118046
rect 173992 117982 174044 117988
rect 174556 3602 174584 151786
rect 174636 144084 174688 144090
rect 174636 144026 174688 144032
rect 174648 3670 174676 144026
rect 175016 142154 175044 154022
rect 175292 153082 175320 158199
rect 175384 153218 175412 160140
rect 175476 155922 175504 160140
rect 175568 158370 175596 160140
rect 175660 158681 175688 160140
rect 175646 158672 175702 158681
rect 175646 158607 175702 158616
rect 175556 158364 175608 158370
rect 175556 158306 175608 158312
rect 175752 157010 175780 160140
rect 175740 157004 175792 157010
rect 175740 156946 175792 156952
rect 175464 155916 175516 155922
rect 175464 155858 175516 155864
rect 175752 155718 175780 156946
rect 175740 155712 175792 155718
rect 175740 155654 175792 155660
rect 175844 154358 175872 160140
rect 175936 159905 175964 160140
rect 175922 159896 175978 159905
rect 175922 159831 175978 159840
rect 175936 158273 175964 159831
rect 176028 158846 176056 160140
rect 176016 158840 176068 158846
rect 176016 158782 176068 158788
rect 175922 158264 175978 158273
rect 175922 158199 175978 158208
rect 175832 154352 175884 154358
rect 175832 154294 175884 154300
rect 175384 153190 175596 153218
rect 175464 153128 175516 153134
rect 175292 153054 175412 153082
rect 175464 153070 175516 153076
rect 175280 152992 175332 152998
rect 175280 152934 175332 152940
rect 174740 142126 175044 142154
rect 174740 133210 174768 142126
rect 174728 133204 174780 133210
rect 174728 133146 174780 133152
rect 175292 16574 175320 152934
rect 175384 147694 175412 153054
rect 175372 147688 175424 147694
rect 175372 147630 175424 147636
rect 175476 144906 175504 153070
rect 175568 146266 175596 153190
rect 176028 152998 176056 158782
rect 176120 157962 176148 160140
rect 176212 159118 176240 160140
rect 176200 159112 176252 159118
rect 176200 159054 176252 159060
rect 176108 157956 176160 157962
rect 176108 157898 176160 157904
rect 176016 152992 176068 152998
rect 176016 152934 176068 152940
rect 176120 151814 176148 157898
rect 176212 155122 176240 159054
rect 176304 155514 176332 160140
rect 176396 159934 176424 160140
rect 176384 159928 176436 159934
rect 176384 159870 176436 159876
rect 176396 158817 176424 159870
rect 176382 158808 176438 158817
rect 176382 158743 176438 158752
rect 176382 158672 176438 158681
rect 176382 158607 176438 158616
rect 176396 157865 176424 158607
rect 176382 157856 176438 157865
rect 176382 157791 176438 157800
rect 176384 155916 176436 155922
rect 176384 155858 176436 155864
rect 176292 155508 176344 155514
rect 176292 155450 176344 155456
rect 176212 155094 176332 155122
rect 176198 153096 176254 153105
rect 176198 153031 176254 153040
rect 176028 151786 176148 151814
rect 175556 146260 175608 146266
rect 175556 146202 175608 146208
rect 175464 144900 175516 144906
rect 175464 144842 175516 144848
rect 176028 28966 176056 151786
rect 176108 146260 176160 146266
rect 176108 146202 176160 146208
rect 176120 145858 176148 146202
rect 176108 145852 176160 145858
rect 176108 145794 176160 145800
rect 176120 130422 176148 145794
rect 176212 144498 176240 153031
rect 176200 144492 176252 144498
rect 176200 144434 176252 144440
rect 176212 144090 176240 144434
rect 176200 144084 176252 144090
rect 176200 144026 176252 144032
rect 176108 130416 176160 130422
rect 176108 130358 176160 130364
rect 176016 28960 176068 28966
rect 176016 28902 176068 28908
rect 175292 16546 175504 16574
rect 174636 3664 174688 3670
rect 174636 3606 174688 3612
rect 174544 3596 174596 3602
rect 174544 3538 174596 3544
rect 175476 480 175504 16546
rect 176304 5574 176332 155094
rect 176292 5568 176344 5574
rect 176292 5510 176344 5516
rect 176396 3534 176424 155858
rect 176488 153134 176516 160140
rect 176580 158642 176608 160140
rect 176568 158636 176620 158642
rect 176568 158578 176620 158584
rect 176580 157622 176608 158578
rect 176568 157616 176620 157622
rect 176568 157558 176620 157564
rect 176568 154352 176620 154358
rect 176568 154294 176620 154300
rect 176580 153202 176608 154294
rect 176568 153196 176620 153202
rect 176568 153138 176620 153144
rect 176476 153128 176528 153134
rect 176476 153070 176528 153076
rect 176672 152640 176700 160140
rect 176764 152862 176792 160140
rect 176856 159118 176884 160140
rect 176844 159112 176896 159118
rect 176844 159054 176896 159060
rect 176856 158642 176884 159054
rect 176844 158636 176896 158642
rect 176844 158578 176896 158584
rect 176844 158500 176896 158506
rect 176844 158442 176896 158448
rect 176856 157758 176884 158442
rect 176844 157752 176896 157758
rect 176844 157694 176896 157700
rect 176752 152856 176804 152862
rect 176752 152798 176804 152804
rect 176580 152612 176700 152640
rect 176580 149734 176608 152612
rect 176660 152516 176712 152522
rect 176660 152458 176712 152464
rect 176568 149728 176620 149734
rect 176568 149670 176620 149676
rect 176568 144900 176620 144906
rect 176568 144842 176620 144848
rect 176580 144362 176608 144842
rect 176568 144356 176620 144362
rect 176568 144298 176620 144304
rect 176580 125594 176608 144298
rect 176568 125588 176620 125594
rect 176568 125530 176620 125536
rect 176672 68338 176700 152458
rect 176948 152454 176976 160140
rect 177040 159769 177068 160140
rect 177026 159760 177082 159769
rect 177026 159695 177082 159704
rect 177040 152522 177068 159695
rect 177132 158642 177160 160140
rect 177120 158636 177172 158642
rect 177120 158578 177172 158584
rect 177120 158500 177172 158506
rect 177120 158442 177172 158448
rect 177132 157894 177160 158442
rect 177120 157888 177172 157894
rect 177224 157865 177252 160140
rect 177316 159905 177344 160140
rect 177302 159896 177358 159905
rect 177302 159831 177358 159840
rect 177120 157830 177172 157836
rect 177210 157856 177266 157865
rect 177132 155990 177160 157830
rect 177210 157791 177266 157800
rect 177120 155984 177172 155990
rect 177120 155926 177172 155932
rect 177316 152522 177344 159831
rect 177408 158506 177436 160140
rect 177396 158500 177448 158506
rect 177396 158442 177448 158448
rect 177396 158228 177448 158234
rect 177396 158170 177448 158176
rect 177028 152516 177080 152522
rect 177028 152458 177080 152464
rect 177304 152516 177356 152522
rect 177304 152458 177356 152464
rect 176936 152448 176988 152454
rect 176936 152390 176988 152396
rect 177408 149546 177436 158170
rect 177500 157690 177528 160140
rect 177592 158681 177620 160140
rect 177684 159934 177712 160140
rect 177672 159928 177724 159934
rect 177672 159870 177724 159876
rect 177578 158672 177634 158681
rect 177578 158607 177634 158616
rect 177684 158234 177712 159870
rect 177672 158228 177724 158234
rect 177672 158170 177724 158176
rect 177776 158137 177804 160140
rect 177762 158128 177818 158137
rect 177762 158063 177818 158072
rect 177868 158001 177896 160140
rect 177854 157992 177910 158001
rect 177854 157927 177910 157936
rect 177672 157752 177724 157758
rect 177672 157694 177724 157700
rect 177488 157684 177540 157690
rect 177488 157626 177540 157632
rect 176856 149518 177436 149546
rect 176856 147626 176884 149518
rect 176844 147620 176896 147626
rect 176844 147562 176896 147568
rect 177500 142154 177528 157626
rect 177684 154834 177712 157694
rect 177960 157334 177988 160140
rect 177776 157306 177988 157334
rect 177672 154828 177724 154834
rect 177672 154770 177724 154776
rect 177776 152538 177804 157306
rect 178052 155786 178080 160140
rect 178144 157334 178172 160140
rect 178236 158914 178264 160140
rect 178224 158908 178276 158914
rect 178224 158850 178276 158856
rect 178144 157306 178264 157334
rect 178040 155780 178092 155786
rect 178040 155722 178092 155728
rect 178040 155508 178092 155514
rect 178040 155450 178092 155456
rect 178052 155242 178080 155450
rect 178040 155236 178092 155242
rect 178040 155178 178092 155184
rect 177316 142126 177528 142154
rect 177592 152510 177804 152538
rect 177948 152516 178000 152522
rect 177316 108322 177344 142126
rect 177592 141506 177620 152510
rect 177948 152458 178000 152464
rect 177764 152448 177816 152454
rect 177764 152390 177816 152396
rect 177776 152114 177804 152390
rect 177764 152108 177816 152114
rect 177764 152050 177816 152056
rect 177580 141500 177632 141506
rect 177580 141442 177632 141448
rect 177776 131782 177804 152050
rect 177764 131776 177816 131782
rect 177764 131718 177816 131724
rect 177304 108316 177356 108322
rect 177304 108258 177356 108264
rect 176660 68332 176712 68338
rect 176660 68274 176712 68280
rect 177960 58682 177988 152458
rect 177948 58676 178000 58682
rect 177948 58618 178000 58624
rect 176660 28960 176712 28966
rect 176660 28902 176712 28908
rect 176384 3528 176436 3534
rect 176384 3470 176436 3476
rect 176672 480 176700 28902
rect 178052 16574 178080 155178
rect 178236 141574 178264 157306
rect 178328 154426 178356 160140
rect 178316 154420 178368 154426
rect 178316 154362 178368 154368
rect 178420 147674 178448 160140
rect 178512 156738 178540 160140
rect 178500 156732 178552 156738
rect 178500 156674 178552 156680
rect 178604 153882 178632 160140
rect 178592 153876 178644 153882
rect 178592 153818 178644 153824
rect 178696 152250 178724 160140
rect 178788 156670 178816 160140
rect 178776 156664 178828 156670
rect 178776 156606 178828 156612
rect 178684 152244 178736 152250
rect 178684 152186 178736 152192
rect 178880 149870 178908 160140
rect 178972 159905 179000 160140
rect 178958 159896 179014 159905
rect 178958 159831 179014 159840
rect 178960 159792 179012 159798
rect 178960 159734 179012 159740
rect 178972 159526 179000 159734
rect 178960 159520 179012 159526
rect 178960 159462 179012 159468
rect 178960 159112 179012 159118
rect 178960 159054 179012 159060
rect 178972 157962 179000 159054
rect 178960 157956 179012 157962
rect 178960 157898 179012 157904
rect 179064 157826 179092 160140
rect 179156 158681 179184 160140
rect 179248 159769 179276 160140
rect 179234 159760 179290 159769
rect 179234 159695 179290 159704
rect 179142 158672 179198 158681
rect 179142 158607 179198 158616
rect 179052 157820 179104 157826
rect 179052 157762 179104 157768
rect 179064 156641 179092 157762
rect 179050 156632 179106 156641
rect 179050 156567 179106 156576
rect 179340 155378 179368 160140
rect 179328 155372 179380 155378
rect 179328 155314 179380 155320
rect 179328 152856 179380 152862
rect 179328 152798 179380 152804
rect 178868 149864 178920 149870
rect 178868 149806 178920 149812
rect 178420 147646 179184 147674
rect 179156 141642 179184 147646
rect 179340 145450 179368 152798
rect 179432 152182 179460 160140
rect 179524 152590 179552 160140
rect 179616 156806 179644 160140
rect 179604 156800 179656 156806
rect 179604 156742 179656 156748
rect 179512 152584 179564 152590
rect 179512 152526 179564 152532
rect 179512 152312 179564 152318
rect 179708 152266 179736 160140
rect 179800 159769 179828 160140
rect 179786 159760 179842 159769
rect 179786 159695 179842 159704
rect 179892 155038 179920 160140
rect 179880 155032 179932 155038
rect 179880 154974 179932 154980
rect 179984 152318 180012 160140
rect 180076 159905 180104 160140
rect 180062 159896 180118 159905
rect 180062 159831 180118 159840
rect 180168 155514 180196 160140
rect 180260 158030 180288 160140
rect 180352 159905 180380 160140
rect 180338 159896 180394 159905
rect 180338 159831 180394 159840
rect 180338 159760 180394 159769
rect 180338 159695 180394 159704
rect 180248 158024 180300 158030
rect 180248 157966 180300 157972
rect 180352 157334 180380 159695
rect 180444 157978 180472 160140
rect 180536 158098 180564 160140
rect 180628 159905 180656 160140
rect 180614 159896 180670 159905
rect 180614 159831 180670 159840
rect 180524 158092 180576 158098
rect 180524 158034 180576 158040
rect 180444 157950 180656 157978
rect 180352 157306 180564 157334
rect 180156 155508 180208 155514
rect 180156 155450 180208 155456
rect 180064 154828 180116 154834
rect 180064 154770 180116 154776
rect 179512 152254 179564 152260
rect 179420 152176 179472 152182
rect 179420 152118 179472 152124
rect 179328 145444 179380 145450
rect 179328 145386 179380 145392
rect 179144 141636 179196 141642
rect 179144 141578 179196 141584
rect 178224 141568 178276 141574
rect 178224 141510 178276 141516
rect 179052 141568 179104 141574
rect 179052 141510 179104 141516
rect 179064 105670 179092 141510
rect 179052 105664 179104 105670
rect 179052 105606 179104 105612
rect 179156 86290 179184 141578
rect 179236 141500 179288 141506
rect 179236 141442 179288 141448
rect 179144 86284 179196 86290
rect 179144 86226 179196 86232
rect 178052 16546 178632 16574
rect 177856 5568 177908 5574
rect 177856 5510 177908 5516
rect 177868 480 177896 5510
rect 174238 354 174350 480
rect 173912 326 174350 354
rect 173134 -960 173246 326
rect 174238 -960 174350 326
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 178604 354 178632 16546
rect 179248 3670 179276 141442
rect 179236 3664 179288 3670
rect 179236 3606 179288 3612
rect 179340 3602 179368 145386
rect 179524 139126 179552 152254
rect 179616 152238 179736 152266
rect 179972 152312 180024 152318
rect 179972 152254 180024 152260
rect 179616 144430 179644 152238
rect 179696 152176 179748 152182
rect 179696 152118 179748 152124
rect 179708 145518 179736 152118
rect 179696 145512 179748 145518
rect 179696 145454 179748 145460
rect 179604 144424 179656 144430
rect 179604 144366 179656 144372
rect 179512 139120 179564 139126
rect 179512 139062 179564 139068
rect 179418 98696 179474 98705
rect 179418 98631 179474 98640
rect 179432 16574 179460 98631
rect 179432 16546 180012 16574
rect 179328 3596 179380 3602
rect 179328 3538 179380 3544
rect 179984 3482 180012 16546
rect 180076 3874 180104 154770
rect 180432 152584 180484 152590
rect 180432 152526 180484 152532
rect 180156 152312 180208 152318
rect 180156 152254 180208 152260
rect 180168 152114 180196 152254
rect 180156 152108 180208 152114
rect 180156 152050 180208 152056
rect 180444 137290 180472 152526
rect 180432 137284 180484 137290
rect 180432 137226 180484 137232
rect 180536 135930 180564 157306
rect 180628 153950 180656 157950
rect 180616 153944 180668 153950
rect 180616 153886 180668 153892
rect 180720 153746 180748 160140
rect 180708 153740 180760 153746
rect 180708 153682 180760 153688
rect 180812 151230 180840 160140
rect 180904 159769 180932 160140
rect 180890 159760 180946 159769
rect 180890 159695 180946 159704
rect 180904 152522 180932 159695
rect 180996 152590 181024 160140
rect 181088 156942 181116 160140
rect 181180 159905 181208 160140
rect 181166 159896 181222 159905
rect 181166 159831 181222 159840
rect 181076 156936 181128 156942
rect 181076 156878 181128 156884
rect 180984 152584 181036 152590
rect 180984 152526 181036 152532
rect 180892 152516 180944 152522
rect 180892 152458 180944 152464
rect 181180 152454 181208 159831
rect 181168 152448 181220 152454
rect 181168 152390 181220 152396
rect 181272 151774 181300 160140
rect 181364 158166 181392 160140
rect 181456 158681 181484 160140
rect 181442 158672 181498 158681
rect 181442 158607 181498 158616
rect 181352 158160 181404 158166
rect 181352 158102 181404 158108
rect 181444 155984 181496 155990
rect 181444 155926 181496 155932
rect 181260 151768 181312 151774
rect 181260 151710 181312 151716
rect 180800 151224 180852 151230
rect 180800 151166 180852 151172
rect 180524 135924 180576 135930
rect 180524 135866 180576 135872
rect 180156 125588 180208 125594
rect 180156 125530 180208 125536
rect 180168 3942 180196 125530
rect 181456 16574 181484 155926
rect 181548 150006 181576 160140
rect 181640 151502 181668 160140
rect 181732 159769 181760 160140
rect 181718 159760 181774 159769
rect 181718 159695 181774 159704
rect 181720 159384 181772 159390
rect 181720 159326 181772 159332
rect 181732 159118 181760 159326
rect 181720 159112 181772 159118
rect 181720 159054 181772 159060
rect 181824 152862 181852 160140
rect 181916 159905 181944 160140
rect 181902 159896 181958 159905
rect 181902 159831 181958 159840
rect 181904 159044 181956 159050
rect 181904 158986 181956 158992
rect 181916 158953 181944 158986
rect 181902 158944 181958 158953
rect 181902 158879 181958 158888
rect 182008 158137 182036 160140
rect 181994 158128 182050 158137
rect 181994 158063 182050 158072
rect 182100 157334 182128 160140
rect 181916 157306 182128 157334
rect 181812 152856 181864 152862
rect 181812 152798 181864 152804
rect 181916 152538 181944 157306
rect 182192 154154 182220 160140
rect 182284 159905 182312 160140
rect 182270 159896 182326 159905
rect 182270 159831 182326 159840
rect 182376 158778 182404 160140
rect 182364 158772 182416 158778
rect 182364 158714 182416 158720
rect 182272 158704 182324 158710
rect 182272 158646 182324 158652
rect 182180 154148 182232 154154
rect 182180 154090 182232 154096
rect 181824 152510 181944 152538
rect 181996 152516 182048 152522
rect 181628 151496 181680 151502
rect 181628 151438 181680 151444
rect 181536 150000 181588 150006
rect 181536 149942 181588 149948
rect 181824 146878 181852 152510
rect 181996 152458 182048 152464
rect 182180 152516 182232 152522
rect 182180 152458 182232 152464
rect 181904 152448 181956 152454
rect 181904 152390 181956 152396
rect 181812 146872 181864 146878
rect 181812 146814 181864 146820
rect 181916 134638 181944 152390
rect 181904 134632 181956 134638
rect 181904 134574 181956 134580
rect 182008 129062 182036 152458
rect 182088 149728 182140 149734
rect 182088 149670 182140 149676
rect 181996 129056 182048 129062
rect 181996 128998 182048 129004
rect 181456 16546 181576 16574
rect 180156 3936 180208 3942
rect 180156 3878 180208 3884
rect 181444 3936 181496 3942
rect 181444 3878 181496 3884
rect 180064 3868 180116 3874
rect 180064 3810 180116 3816
rect 179984 3454 180288 3482
rect 180260 480 180288 3454
rect 181456 480 181484 3878
rect 181548 3466 181576 16546
rect 182100 3534 182128 149670
rect 182088 3528 182140 3534
rect 182088 3470 182140 3476
rect 181536 3460 181588 3466
rect 181536 3402 181588 3408
rect 179022 354 179134 480
rect 178604 326 179134 354
rect 179022 -960 179134 326
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182192 354 182220 152458
rect 182284 143070 182312 158646
rect 182468 154970 182496 160140
rect 182560 159594 182588 160140
rect 182548 159588 182600 159594
rect 182548 159530 182600 159536
rect 182560 158681 182588 159530
rect 182546 158672 182602 158681
rect 182546 158607 182602 158616
rect 182456 154964 182508 154970
rect 182456 154906 182508 154912
rect 182652 151638 182680 160140
rect 182744 158506 182772 160140
rect 182836 159905 182864 160140
rect 182822 159896 182878 159905
rect 182822 159831 182878 159840
rect 182732 158500 182784 158506
rect 182732 158442 182784 158448
rect 182836 158137 182864 159831
rect 182822 158128 182878 158137
rect 182822 158063 182878 158072
rect 182732 157616 182784 157622
rect 182732 157558 182784 157564
rect 182744 152522 182772 157558
rect 182928 154222 182956 160140
rect 182916 154216 182968 154222
rect 182916 154158 182968 154164
rect 182732 152516 182784 152522
rect 182732 152458 182784 152464
rect 182640 151632 182692 151638
rect 182640 151574 182692 151580
rect 183020 149530 183048 160140
rect 183112 158681 183140 160140
rect 183098 158672 183154 158681
rect 183098 158607 183154 158616
rect 183204 157334 183232 160140
rect 183296 159905 183324 160140
rect 183282 159896 183338 159905
rect 183282 159831 183338 159840
rect 183388 159769 183416 160140
rect 183374 159760 183430 159769
rect 183374 159695 183430 159704
rect 183284 158772 183336 158778
rect 183284 158714 183336 158720
rect 183112 157306 183232 157334
rect 183008 149524 183060 149530
rect 183008 149466 183060 149472
rect 183112 149410 183140 157306
rect 183192 154148 183244 154154
rect 183192 154090 183244 154096
rect 183204 150958 183232 154090
rect 183296 152930 183324 158714
rect 183480 158710 183508 160140
rect 183468 158704 183520 158710
rect 183468 158646 183520 158652
rect 183466 158128 183522 158137
rect 183466 158063 183522 158072
rect 183284 152924 183336 152930
rect 183284 152866 183336 152872
rect 183192 150952 183244 150958
rect 183192 150894 183244 150900
rect 182376 149382 183140 149410
rect 182376 147422 182404 149382
rect 182824 147620 182876 147626
rect 182824 147562 182876 147568
rect 182364 147416 182416 147422
rect 182364 147358 182416 147364
rect 182272 143064 182324 143070
rect 182272 143006 182324 143012
rect 182836 3398 182864 147562
rect 183480 111110 183508 158063
rect 183572 151434 183600 160140
rect 183664 158778 183692 160140
rect 183652 158772 183704 158778
rect 183652 158714 183704 158720
rect 183756 155106 183784 160140
rect 183744 155100 183796 155106
rect 183744 155042 183796 155048
rect 183848 153678 183876 160140
rect 183940 159905 183968 160140
rect 183926 159896 183982 159905
rect 183926 159831 183982 159840
rect 183836 153672 183888 153678
rect 183836 153614 183888 153620
rect 183744 152516 183796 152522
rect 183744 152458 183796 152464
rect 183652 152448 183704 152454
rect 183652 152390 183704 152396
rect 183560 151428 183612 151434
rect 183560 151370 183612 151376
rect 183664 141846 183692 152390
rect 183756 146062 183784 152458
rect 184032 150278 184060 160140
rect 184124 158234 184152 160140
rect 184216 159905 184244 160140
rect 184202 159896 184258 159905
rect 184202 159831 184258 159840
rect 184204 158908 184256 158914
rect 184204 158850 184256 158856
rect 184216 158778 184244 158850
rect 184204 158772 184256 158778
rect 184204 158714 184256 158720
rect 184112 158228 184164 158234
rect 184112 158170 184164 158176
rect 184112 157956 184164 157962
rect 184112 157898 184164 157904
rect 184020 150272 184072 150278
rect 184020 150214 184072 150220
rect 184124 147674 184152 157898
rect 184216 152538 184244 158714
rect 184308 157334 184336 160140
rect 184400 158710 184428 160140
rect 184492 159769 184520 160140
rect 184478 159760 184534 159769
rect 184478 159695 184534 159704
rect 184388 158704 184440 158710
rect 184388 158646 184440 158652
rect 184308 157306 184428 157334
rect 184216 152510 184336 152538
rect 184308 147674 184336 152510
rect 184400 148850 184428 157306
rect 184584 152522 184612 160140
rect 184572 152516 184624 152522
rect 184572 152458 184624 152464
rect 184388 148844 184440 148850
rect 184388 148786 184440 148792
rect 184676 148714 184704 160140
rect 184768 159497 184796 160140
rect 184754 159488 184810 159497
rect 184754 159423 184810 159432
rect 184756 158636 184808 158642
rect 184756 158578 184808 158584
rect 184768 157962 184796 158578
rect 184756 157956 184808 157962
rect 184756 157898 184808 157904
rect 184860 152454 184888 160140
rect 184952 153474 184980 160140
rect 185044 158681 185072 160140
rect 185030 158672 185086 158681
rect 185030 158607 185086 158616
rect 185136 157334 185164 160140
rect 185228 157826 185256 160140
rect 185216 157820 185268 157826
rect 185216 157762 185268 157768
rect 185320 157334 185348 160140
rect 185412 159662 185440 160140
rect 185400 159656 185452 159662
rect 185400 159598 185452 159604
rect 185044 157306 185164 157334
rect 185228 157306 185348 157334
rect 184940 153468 184992 153474
rect 184940 153410 184992 153416
rect 184848 152448 184900 152454
rect 184848 152390 184900 152396
rect 184940 152448 184992 152454
rect 184940 152390 184992 152396
rect 184664 148708 184716 148714
rect 184664 148650 184716 148656
rect 184124 147646 184244 147674
rect 184308 147646 184612 147674
rect 183744 146056 183796 146062
rect 183744 145998 183796 146004
rect 183652 141840 183704 141846
rect 183652 141782 183704 141788
rect 183468 111104 183520 111110
rect 183468 111046 183520 111052
rect 183744 3528 183796 3534
rect 183744 3470 183796 3476
rect 182824 3392 182876 3398
rect 182824 3334 182876 3340
rect 183756 480 183784 3470
rect 184216 3058 184244 147646
rect 184584 119406 184612 147646
rect 184952 140554 184980 152390
rect 185044 143478 185072 157306
rect 185228 152538 185256 157306
rect 185504 154018 185532 160140
rect 185492 154012 185544 154018
rect 185492 153954 185544 153960
rect 185136 152510 185256 152538
rect 185136 143546 185164 152510
rect 185596 148646 185624 160140
rect 185688 151570 185716 160140
rect 185780 157486 185808 160140
rect 185872 158681 185900 160140
rect 185858 158672 185914 158681
rect 185858 158607 185914 158616
rect 185768 157480 185820 157486
rect 185768 157422 185820 157428
rect 185964 157334 185992 160140
rect 185780 157306 185992 157334
rect 185676 151564 185728 151570
rect 185676 151506 185728 151512
rect 185584 148640 185636 148646
rect 185584 148582 185636 148588
rect 185780 148458 185808 157306
rect 186056 156602 186084 160140
rect 186044 156596 186096 156602
rect 186044 156538 186096 156544
rect 185860 153468 185912 153474
rect 185860 153410 185912 153416
rect 185872 149598 185900 153410
rect 185860 149592 185912 149598
rect 185860 149534 185912 149540
rect 185228 148430 185808 148458
rect 185228 144838 185256 148430
rect 186148 147674 186176 160140
rect 186240 152454 186268 160140
rect 186332 158817 186360 160140
rect 186318 158808 186374 158817
rect 186318 158743 186374 158752
rect 186320 158704 186372 158710
rect 186320 158646 186372 158652
rect 186332 158302 186360 158646
rect 186320 158296 186372 158302
rect 186320 158238 186372 158244
rect 186320 152652 186372 152658
rect 186320 152594 186372 152600
rect 186228 152448 186280 152454
rect 186228 152390 186280 152396
rect 185320 147646 186176 147674
rect 185320 145926 185348 147646
rect 185308 145920 185360 145926
rect 185308 145862 185360 145868
rect 185216 144832 185268 144838
rect 185216 144774 185268 144780
rect 185124 143540 185176 143546
rect 185124 143482 185176 143488
rect 186228 143540 186280 143546
rect 186228 143482 186280 143488
rect 185032 143472 185084 143478
rect 185032 143414 185084 143420
rect 186240 143138 186268 143482
rect 186228 143132 186280 143138
rect 186228 143074 186280 143080
rect 186134 141264 186190 141273
rect 186134 141199 186190 141208
rect 186148 140865 186176 141199
rect 186134 140856 186190 140865
rect 186134 140791 186190 140800
rect 184940 140548 184992 140554
rect 184940 140490 184992 140496
rect 184572 119400 184624 119406
rect 184572 119342 184624 119348
rect 184296 108316 184348 108322
rect 184296 108258 184348 108264
rect 184308 3942 184336 108258
rect 186148 6914 186176 140791
rect 186056 6886 186176 6914
rect 184296 3936 184348 3942
rect 184296 3878 184348 3884
rect 186056 3738 186084 6886
rect 186044 3732 186096 3738
rect 186044 3674 186096 3680
rect 186240 3602 186268 143074
rect 186332 133754 186360 152594
rect 186320 133748 186372 133754
rect 186320 133690 186372 133696
rect 186320 131776 186372 131782
rect 186320 131718 186372 131724
rect 186332 16574 186360 131718
rect 186424 126954 186452 160140
rect 186516 159934 186544 160140
rect 186504 159928 186556 159934
rect 186504 159870 186556 159876
rect 186504 157956 186556 157962
rect 186504 157898 186556 157904
rect 186516 152590 186544 157898
rect 186608 152674 186636 160140
rect 186700 158681 186728 160140
rect 186686 158672 186742 158681
rect 186686 158607 186742 158616
rect 186608 152646 186728 152674
rect 186504 152584 186556 152590
rect 186504 152526 186556 152532
rect 186596 152448 186648 152454
rect 186596 152390 186648 152396
rect 186504 152176 186556 152182
rect 186504 152118 186556 152124
rect 186516 132326 186544 152118
rect 186608 139398 186636 152390
rect 186700 151706 186728 152646
rect 186688 151700 186740 151706
rect 186688 151642 186740 151648
rect 186792 147674 186820 160140
rect 186884 158642 186912 160140
rect 186872 158636 186924 158642
rect 186872 158578 186924 158584
rect 186976 158137 187004 160140
rect 186962 158128 187018 158137
rect 186962 158063 187018 158072
rect 186964 152584 187016 152590
rect 186964 152526 187016 152532
rect 186700 147646 186820 147674
rect 186700 143546 186728 147646
rect 186688 143540 186740 143546
rect 186688 143482 186740 143488
rect 186596 139392 186648 139398
rect 186596 139334 186648 139340
rect 186504 132320 186556 132326
rect 186504 132262 186556 132268
rect 186412 126948 186464 126954
rect 186412 126890 186464 126896
rect 186332 16546 186912 16574
rect 184940 3596 184992 3602
rect 184940 3538 184992 3544
rect 186228 3596 186280 3602
rect 186228 3538 186280 3544
rect 184204 3052 184256 3058
rect 184204 2994 184256 3000
rect 184952 480 184980 3538
rect 186136 3052 186188 3058
rect 186136 2994 186188 3000
rect 186148 480 186176 2994
rect 182518 354 182630 480
rect 182192 326 182630 354
rect 182518 -960 182630 326
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 186884 354 186912 16546
rect 186976 3806 187004 152526
rect 187068 152454 187096 160140
rect 187160 158574 187188 160140
rect 187252 158681 187280 160140
rect 187238 158672 187294 158681
rect 187238 158607 187294 158616
rect 187148 158568 187200 158574
rect 187148 158510 187200 158516
rect 187240 157480 187292 157486
rect 187240 157422 187292 157428
rect 187056 152448 187108 152454
rect 187056 152390 187108 152396
rect 187252 149666 187280 157422
rect 187344 152658 187372 160140
rect 187436 157334 187464 160140
rect 187528 158681 187556 160140
rect 187514 158672 187570 158681
rect 187514 158607 187570 158616
rect 187436 157306 187556 157334
rect 187528 155922 187556 157306
rect 187516 155916 187568 155922
rect 187516 155858 187568 155864
rect 187332 152652 187384 152658
rect 187332 152594 187384 152600
rect 187620 152182 187648 160140
rect 187712 152998 187740 160140
rect 187804 153082 187832 160140
rect 187896 153762 187924 160140
rect 187988 154154 188016 160140
rect 188080 158681 188108 160140
rect 188066 158672 188122 158681
rect 188066 158607 188122 158616
rect 187976 154148 188028 154154
rect 187976 154090 188028 154096
rect 187896 153734 188108 153762
rect 187804 153054 188016 153082
rect 187700 152992 187752 152998
rect 187700 152934 187752 152940
rect 187700 152584 187752 152590
rect 187700 152526 187752 152532
rect 187608 152176 187660 152182
rect 187608 152118 187660 152124
rect 187240 149660 187292 149666
rect 187240 149602 187292 149608
rect 187712 142118 187740 152526
rect 187792 152448 187844 152454
rect 187792 152390 187844 152396
rect 187804 143274 187832 152390
rect 187988 148782 188016 153054
rect 188080 150210 188108 153734
rect 188068 150204 188120 150210
rect 188068 150146 188120 150152
rect 187976 148776 188028 148782
rect 187976 148718 188028 148724
rect 188172 147674 188200 160140
rect 188264 158710 188292 160140
rect 188356 159905 188384 160140
rect 188342 159896 188398 159905
rect 188342 159831 188398 159840
rect 188448 159089 188476 160140
rect 188434 159080 188490 159089
rect 188434 159015 188490 159024
rect 188540 158930 188568 160140
rect 188356 158902 188568 158930
rect 188252 158704 188304 158710
rect 188252 158646 188304 158652
rect 188356 158506 188384 158902
rect 188434 158808 188490 158817
rect 188434 158743 188490 158752
rect 188252 158500 188304 158506
rect 188252 158442 188304 158448
rect 188344 158500 188396 158506
rect 188344 158442 188396 158448
rect 188264 157758 188292 158442
rect 188252 157752 188304 157758
rect 188252 157694 188304 157700
rect 188448 152454 188476 158743
rect 188632 158681 188660 160140
rect 188618 158672 188674 158681
rect 188528 158636 188580 158642
rect 188618 158607 188674 158616
rect 188528 158578 188580 158584
rect 188436 152448 188488 152454
rect 188436 152390 188488 152396
rect 188540 151298 188568 158578
rect 188724 152590 188752 160140
rect 188816 154902 188844 160140
rect 188804 154896 188856 154902
rect 188804 154838 188856 154844
rect 188908 153066 188936 160140
rect 189000 157321 189028 160140
rect 188986 157312 189042 157321
rect 188986 157247 189042 157256
rect 189092 153814 189120 160140
rect 189184 158681 189212 160140
rect 189170 158672 189226 158681
rect 189170 158607 189226 158616
rect 189080 153808 189132 153814
rect 189080 153750 189132 153756
rect 189276 153134 189304 160140
rect 189368 158846 189396 160140
rect 189356 158840 189408 158846
rect 189356 158782 189408 158788
rect 189356 158704 189408 158710
rect 189356 158646 189408 158652
rect 189368 156874 189396 158646
rect 189356 156868 189408 156874
rect 189356 156810 189408 156816
rect 189264 153128 189316 153134
rect 189264 153070 189316 153076
rect 188896 153060 188948 153066
rect 188896 153002 188948 153008
rect 189460 152674 189488 160140
rect 189276 152646 189488 152674
rect 188712 152584 188764 152590
rect 188712 152526 188764 152532
rect 189080 152584 189132 152590
rect 189080 152526 189132 152532
rect 188528 151292 188580 151298
rect 188528 151234 188580 151240
rect 187896 147646 188200 147674
rect 187896 147558 187924 147646
rect 187884 147552 187936 147558
rect 187884 147494 187936 147500
rect 187792 143268 187844 143274
rect 187792 143210 187844 143216
rect 187700 142112 187752 142118
rect 187700 142054 187752 142060
rect 189092 125526 189120 152526
rect 189172 152448 189224 152454
rect 189172 152390 189224 152396
rect 189184 136474 189212 152390
rect 189276 141778 189304 152646
rect 189552 152538 189580 160140
rect 189644 159769 189672 160140
rect 189736 159905 189764 160140
rect 189722 159896 189778 159905
rect 189722 159831 189778 159840
rect 189630 159760 189686 159769
rect 189630 159695 189686 159704
rect 189632 158840 189684 158846
rect 189632 158782 189684 158788
rect 189644 157486 189672 158782
rect 189632 157480 189684 157486
rect 189632 157422 189684 157428
rect 189632 153128 189684 153134
rect 189632 153070 189684 153076
rect 189368 152510 189580 152538
rect 189368 144770 189396 152510
rect 189644 148170 189672 153070
rect 189828 152454 189856 160140
rect 189920 158710 189948 160140
rect 189908 158704 189960 158710
rect 190012 158681 190040 160140
rect 189908 158646 189960 158652
rect 189998 158672 190054 158681
rect 189998 158607 190054 158616
rect 189908 158568 189960 158574
rect 189908 158510 189960 158516
rect 189816 152448 189868 152454
rect 189816 152390 189868 152396
rect 189920 151366 189948 158510
rect 189908 151360 189960 151366
rect 189908 151302 189960 151308
rect 189632 148164 189684 148170
rect 189632 148106 189684 148112
rect 190104 147674 190132 160140
rect 190196 159526 190224 160140
rect 190184 159520 190236 159526
rect 190184 159462 190236 159468
rect 190288 158681 190316 160140
rect 190274 158672 190330 158681
rect 190274 158607 190330 158616
rect 190184 158568 190236 158574
rect 190184 158510 190236 158516
rect 190196 158030 190224 158510
rect 190276 158160 190328 158166
rect 190276 158102 190328 158108
rect 190184 158024 190236 158030
rect 190184 157966 190236 157972
rect 190288 157826 190316 158102
rect 190184 157820 190236 157826
rect 190184 157762 190236 157768
rect 190276 157820 190328 157826
rect 190276 157762 190328 157768
rect 190196 150074 190224 157762
rect 190380 152590 190408 160140
rect 190472 158794 190500 160140
rect 190564 158953 190592 160140
rect 190550 158944 190606 158953
rect 190550 158879 190606 158888
rect 190472 158766 190592 158794
rect 190458 158128 190514 158137
rect 190458 158063 190514 158072
rect 190368 152584 190420 152590
rect 190368 152526 190420 152532
rect 190184 150068 190236 150074
rect 190184 150010 190236 150016
rect 189460 147646 190132 147674
rect 189460 145994 189488 147646
rect 189448 145988 189500 145994
rect 189448 145930 189500 145936
rect 189356 144764 189408 144770
rect 189356 144706 189408 144712
rect 189264 141772 189316 141778
rect 189264 141714 189316 141720
rect 190368 141772 190420 141778
rect 190368 141714 190420 141720
rect 189722 141536 189778 141545
rect 189722 141471 189778 141480
rect 189172 136468 189224 136474
rect 189172 136410 189224 136416
rect 189080 125520 189132 125526
rect 189080 125462 189132 125468
rect 187700 68332 187752 68338
rect 187700 68274 187752 68280
rect 187712 16574 187740 68274
rect 189736 16574 189764 141471
rect 190380 105602 190408 141714
rect 190368 105596 190420 105602
rect 190368 105538 190420 105544
rect 187712 16546 188568 16574
rect 189736 16546 189856 16574
rect 186964 3800 187016 3806
rect 186964 3742 187016 3748
rect 188540 480 188568 16546
rect 189724 3868 189776 3874
rect 189724 3810 189776 3816
rect 189736 480 189764 3810
rect 189828 3126 189856 16546
rect 190472 10334 190500 158063
rect 190564 152658 190592 158766
rect 190552 152652 190604 152658
rect 190552 152594 190604 152600
rect 190656 152538 190684 160140
rect 190748 155174 190776 160140
rect 190840 159905 190868 160140
rect 190826 159896 190882 159905
rect 190826 159831 190882 159840
rect 190828 159180 190880 159186
rect 190828 159122 190880 159128
rect 190840 155825 190868 159122
rect 190826 155816 190882 155825
rect 190826 155751 190882 155760
rect 190736 155168 190788 155174
rect 190736 155110 190788 155116
rect 190656 152510 190776 152538
rect 190644 152448 190696 152454
rect 190644 152390 190696 152396
rect 190656 140758 190684 152390
rect 190748 146130 190776 152510
rect 190932 152454 190960 160140
rect 191024 158166 191052 160140
rect 191116 159769 191144 160140
rect 191102 159760 191158 159769
rect 191102 159695 191158 159704
rect 191208 158794 191236 160140
rect 191300 159186 191328 160140
rect 191392 159905 191420 160140
rect 191378 159896 191434 159905
rect 191378 159831 191434 159840
rect 191288 159180 191340 159186
rect 191288 159122 191340 159128
rect 191208 158766 191328 158794
rect 191196 158500 191248 158506
rect 191196 158442 191248 158448
rect 191012 158160 191064 158166
rect 191012 158102 191064 158108
rect 191104 158092 191156 158098
rect 191104 158034 191156 158040
rect 191116 157622 191144 158034
rect 191104 157616 191156 157622
rect 191104 157558 191156 157564
rect 191104 157140 191156 157146
rect 191104 157082 191156 157088
rect 191116 156602 191144 157082
rect 191104 156596 191156 156602
rect 191104 156538 191156 156544
rect 190920 152448 190972 152454
rect 190920 152390 190972 152396
rect 191208 148578 191236 158442
rect 191196 148572 191248 148578
rect 191196 148514 191248 148520
rect 191300 148510 191328 158766
rect 191484 157334 191512 160140
rect 191576 157962 191604 160140
rect 191668 159497 191696 160140
rect 191654 159488 191710 159497
rect 191654 159423 191710 159432
rect 191668 158137 191696 159423
rect 191654 158128 191710 158137
rect 191654 158063 191710 158072
rect 191564 157956 191616 157962
rect 191564 157898 191616 157904
rect 191760 157334 191788 160140
rect 191392 157306 191512 157334
rect 191576 157306 191788 157334
rect 191288 148504 191340 148510
rect 191288 148446 191340 148452
rect 191392 148374 191420 157306
rect 191576 148594 191604 157306
rect 191852 149802 191880 160140
rect 191944 158681 191972 160140
rect 192036 159934 192064 160140
rect 192024 159928 192076 159934
rect 192024 159870 192076 159876
rect 191930 158672 191986 158681
rect 191930 158607 191986 158616
rect 192024 158296 192076 158302
rect 192024 158238 192076 158244
rect 192036 152697 192064 158238
rect 192128 158030 192156 160140
rect 192220 159769 192248 160140
rect 192206 159760 192262 159769
rect 192206 159695 192262 159704
rect 192116 158024 192168 158030
rect 192116 157966 192168 157972
rect 192022 152688 192078 152697
rect 192022 152623 192078 152632
rect 191932 152448 191984 152454
rect 191932 152390 191984 152396
rect 191840 149796 191892 149802
rect 191840 149738 191892 149744
rect 191484 148566 191604 148594
rect 191380 148368 191432 148374
rect 191380 148310 191432 148316
rect 190736 146124 190788 146130
rect 190736 146066 190788 146072
rect 190644 140752 190696 140758
rect 190644 140694 190696 140700
rect 191484 133890 191512 148566
rect 191564 148504 191616 148510
rect 191564 148446 191616 148452
rect 191576 135250 191604 148446
rect 191564 135244 191616 135250
rect 191564 135186 191616 135192
rect 191472 133884 191524 133890
rect 191472 133826 191524 133832
rect 191944 126818 191972 152390
rect 192220 152182 192248 159695
rect 192208 152176 192260 152182
rect 192208 152118 192260 152124
rect 192312 150890 192340 160140
rect 192404 157593 192432 160140
rect 192496 159905 192524 160140
rect 192482 159896 192538 159905
rect 192482 159831 192538 159840
rect 192390 157584 192446 157593
rect 192390 157519 192446 157528
rect 192390 157312 192446 157321
rect 192390 157247 192446 157256
rect 192404 154562 192432 157247
rect 192496 156097 192524 159831
rect 192482 156088 192538 156097
rect 192482 156023 192538 156032
rect 192392 154556 192444 154562
rect 192392 154498 192444 154504
rect 192300 150884 192352 150890
rect 192300 150826 192352 150832
rect 192588 147674 192616 160140
rect 192680 158098 192708 160140
rect 192772 159905 192800 160140
rect 192758 159896 192814 159905
rect 192758 159831 192814 159840
rect 192668 158092 192720 158098
rect 192668 158034 192720 158040
rect 192668 157480 192720 157486
rect 192668 157422 192720 157428
rect 192680 148442 192708 157422
rect 192864 152454 192892 160140
rect 192956 156534 192984 160140
rect 193048 158681 193076 160140
rect 193034 158672 193090 158681
rect 193034 158607 193090 158616
rect 193140 157334 193168 160140
rect 193048 157306 193168 157334
rect 193232 157334 193260 160140
rect 193324 158137 193352 160140
rect 193310 158128 193366 158137
rect 193310 158063 193366 158072
rect 193232 157306 193352 157334
rect 192944 156528 192996 156534
rect 192944 156470 192996 156476
rect 193048 152538 193076 157306
rect 193126 156088 193182 156097
rect 193126 156023 193182 156032
rect 192956 152510 193076 152538
rect 192852 152448 192904 152454
rect 192852 152390 192904 152396
rect 192668 148436 192720 148442
rect 192668 148378 192720 148384
rect 192036 147646 192616 147674
rect 192036 132462 192064 147646
rect 192024 132456 192076 132462
rect 192024 132398 192076 132404
rect 191932 126812 191984 126818
rect 191932 126754 191984 126760
rect 192956 124166 192984 152510
rect 193140 152402 193168 156023
rect 193048 152374 193168 152402
rect 192944 124160 192996 124166
rect 192944 124102 192996 124108
rect 191104 58676 191156 58682
rect 191104 58618 191156 58624
rect 190460 10328 190512 10334
rect 190460 10270 190512 10276
rect 191116 3534 191144 58618
rect 193048 6254 193076 152374
rect 193128 152176 193180 152182
rect 193324 152153 193352 157306
rect 193416 155281 193444 160140
rect 193508 158166 193536 160140
rect 193600 159905 193628 160140
rect 193586 159896 193642 159905
rect 193586 159831 193642 159840
rect 193496 158160 193548 158166
rect 193496 158102 193548 158108
rect 193692 157334 193720 160140
rect 193784 159934 193812 160140
rect 193772 159928 193824 159934
rect 193772 159870 193824 159876
rect 193508 157306 193720 157334
rect 193402 155272 193458 155281
rect 193402 155207 193458 155216
rect 193508 152538 193536 157306
rect 193416 152510 193536 152538
rect 193128 152118 193180 152124
rect 193310 152144 193366 152153
rect 193140 6322 193168 152118
rect 193220 152108 193272 152114
rect 193310 152079 193366 152088
rect 193220 152050 193272 152056
rect 193232 117298 193260 152050
rect 193312 152040 193364 152046
rect 193312 151982 193364 151988
rect 193324 131102 193352 151982
rect 193416 139330 193444 152510
rect 193496 152176 193548 152182
rect 193496 152118 193548 152124
rect 193586 152144 193642 152153
rect 193508 147354 193536 152118
rect 193876 152114 193904 160140
rect 193586 152079 193642 152088
rect 193864 152108 193916 152114
rect 193496 147348 193548 147354
rect 193496 147290 193548 147296
rect 193600 147150 193628 152079
rect 193864 152050 193916 152056
rect 193968 147218 193996 160140
rect 194060 152182 194088 160140
rect 194152 158681 194180 160140
rect 194138 158672 194194 158681
rect 194138 158607 194194 158616
rect 194140 158024 194192 158030
rect 194140 157966 194192 157972
rect 194048 152176 194100 152182
rect 194048 152118 194100 152124
rect 194152 148510 194180 157966
rect 194244 152046 194272 160140
rect 194336 158642 194364 160140
rect 194428 159905 194456 160140
rect 194414 159896 194470 159905
rect 194414 159831 194470 159840
rect 194416 158704 194468 158710
rect 194416 158646 194468 158652
rect 194324 158636 194376 158642
rect 194324 158578 194376 158584
rect 194232 152040 194284 152046
rect 194232 151982 194284 151988
rect 194140 148504 194192 148510
rect 194140 148446 194192 148452
rect 194428 148238 194456 158646
rect 194520 156777 194548 160140
rect 194506 156768 194562 156777
rect 194506 156703 194562 156712
rect 194416 148232 194468 148238
rect 194416 148174 194468 148180
rect 193956 147212 194008 147218
rect 193956 147154 194008 147160
rect 193588 147144 193640 147150
rect 193588 147086 193640 147092
rect 193404 139324 193456 139330
rect 193404 139266 193456 139272
rect 193312 131096 193364 131102
rect 193312 131038 193364 131044
rect 194520 122126 194548 156703
rect 194612 152590 194640 160140
rect 194704 158137 194732 160140
rect 194690 158128 194746 158137
rect 194690 158063 194746 158072
rect 194600 152584 194652 152590
rect 194600 152526 194652 152532
rect 194692 151836 194744 151842
rect 194692 151778 194744 151784
rect 194704 137970 194732 151778
rect 194796 142050 194824 160140
rect 194888 157334 194916 160140
rect 194980 159905 195008 160140
rect 194966 159896 195022 159905
rect 194966 159831 195022 159840
rect 194888 157306 195008 157334
rect 194876 152584 194928 152590
rect 194876 152526 194928 152532
rect 194888 147082 194916 152526
rect 194980 149977 195008 157306
rect 195072 151842 195100 160140
rect 195164 158710 195192 160140
rect 195256 159769 195284 160140
rect 195242 159760 195298 159769
rect 195242 159695 195298 159704
rect 195348 158794 195376 160140
rect 195440 159458 195468 160140
rect 195428 159452 195480 159458
rect 195428 159394 195480 159400
rect 195532 159186 195560 160140
rect 195520 159180 195572 159186
rect 195520 159122 195572 159128
rect 195348 158766 195560 158794
rect 195152 158704 195204 158710
rect 195152 158646 195204 158652
rect 195428 157820 195480 157826
rect 195428 157762 195480 157768
rect 195336 157752 195388 157758
rect 195336 157694 195388 157700
rect 195060 151836 195112 151842
rect 195060 151778 195112 151784
rect 195348 150142 195376 157694
rect 195440 151162 195468 157762
rect 195428 151156 195480 151162
rect 195428 151098 195480 151104
rect 195336 150136 195388 150142
rect 195336 150078 195388 150084
rect 194966 149968 195022 149977
rect 194966 149903 195022 149912
rect 195532 147674 195560 158766
rect 195624 158681 195652 160140
rect 195610 158672 195666 158681
rect 195610 158607 195666 158616
rect 195612 157888 195664 157894
rect 195612 157830 195664 157836
rect 195624 153610 195652 157830
rect 195716 157690 195744 160140
rect 195808 159905 195836 160140
rect 195794 159896 195850 159905
rect 195794 159831 195850 159840
rect 195900 158794 195928 160140
rect 195808 158766 195928 158794
rect 195704 157684 195756 157690
rect 195704 157626 195756 157632
rect 195808 156262 195836 158766
rect 195886 158672 195942 158681
rect 195886 158607 195942 158616
rect 195796 156256 195848 156262
rect 195796 156198 195848 156204
rect 195612 153604 195664 153610
rect 195612 153546 195664 153552
rect 195532 147646 195744 147674
rect 194876 147076 194928 147082
rect 194876 147018 194928 147024
rect 194784 142044 194836 142050
rect 194784 141986 194836 141992
rect 194692 137964 194744 137970
rect 194692 137906 194744 137912
rect 195716 129742 195744 147646
rect 195704 129736 195756 129742
rect 195704 129678 195756 129684
rect 194508 122120 194560 122126
rect 194508 122062 194560 122068
rect 193220 117292 193272 117298
rect 193220 117234 193272 117240
rect 193862 28248 193918 28257
rect 193862 28183 193918 28192
rect 193128 6316 193180 6322
rect 193128 6258 193180 6264
rect 193036 6248 193088 6254
rect 193036 6190 193088 6196
rect 193876 3534 193904 28183
rect 195900 9110 195928 158607
rect 195992 157486 196020 160140
rect 196084 158681 196112 160140
rect 196176 158846 196204 160140
rect 196164 158840 196216 158846
rect 196164 158782 196216 158788
rect 196070 158672 196126 158681
rect 196070 158607 196126 158616
rect 196070 158128 196126 158137
rect 196070 158063 196126 158072
rect 195980 157480 196032 157486
rect 195980 157422 196032 157428
rect 195980 152788 196032 152794
rect 195980 152730 196032 152736
rect 195992 128246 196020 152730
rect 195980 128240 196032 128246
rect 195980 128182 196032 128188
rect 195888 9104 195940 9110
rect 195888 9046 195940 9052
rect 196084 8974 196112 158063
rect 196164 152448 196216 152454
rect 196164 152390 196216 152396
rect 196176 144158 196204 152390
rect 196268 146674 196296 160140
rect 196360 159905 196388 160140
rect 196346 159896 196402 159905
rect 196346 159831 196402 159840
rect 196348 158092 196400 158098
rect 196348 158034 196400 158040
rect 196360 147121 196388 158034
rect 196452 152454 196480 160140
rect 196544 158506 196572 160140
rect 196636 159769 196664 160140
rect 196622 159760 196678 159769
rect 196622 159695 196678 159704
rect 196624 158704 196676 158710
rect 196624 158646 196676 158652
rect 196532 158500 196584 158506
rect 196532 158442 196584 158448
rect 196440 152448 196492 152454
rect 196440 152390 196492 152396
rect 196636 151473 196664 158646
rect 196622 151464 196678 151473
rect 196622 151399 196678 151408
rect 196728 147674 196756 160140
rect 196820 155961 196848 160140
rect 196912 159905 196940 160140
rect 196898 159896 196954 159905
rect 196898 159831 196954 159840
rect 196806 155952 196862 155961
rect 196806 155887 196862 155896
rect 197004 152794 197032 160140
rect 197096 153649 197124 160140
rect 197188 159905 197216 160140
rect 197174 159896 197230 159905
rect 197174 159831 197230 159840
rect 197176 158840 197228 158846
rect 197176 158782 197228 158788
rect 197082 153640 197138 153649
rect 197082 153575 197138 153584
rect 197188 152794 197216 158782
rect 197280 158681 197308 160140
rect 197266 158672 197322 158681
rect 197266 158607 197322 158616
rect 197372 157894 197400 160140
rect 197360 157888 197412 157894
rect 197360 157830 197412 157836
rect 197464 154426 197492 160140
rect 197452 154420 197504 154426
rect 197452 154362 197504 154368
rect 197556 153898 197584 160140
rect 197372 153870 197584 153898
rect 196992 152788 197044 152794
rect 196992 152730 197044 152736
rect 197176 152788 197228 152794
rect 197176 152730 197228 152736
rect 196728 147646 197032 147674
rect 196346 147112 196402 147121
rect 196346 147047 196402 147056
rect 196256 146668 196308 146674
rect 196256 146610 196308 146616
rect 196164 144152 196216 144158
rect 196164 144094 196216 144100
rect 197004 136610 197032 147646
rect 197082 144392 197138 144401
rect 197082 144327 197138 144336
rect 197096 142866 197124 144327
rect 197084 142860 197136 142866
rect 197084 142802 197136 142808
rect 196992 136604 197044 136610
rect 196992 136546 197044 136552
rect 196622 17232 196678 17241
rect 196622 17167 196678 17176
rect 196072 8968 196124 8974
rect 196072 8910 196124 8916
rect 194416 3936 194468 3942
rect 194416 3878 194468 3884
rect 191104 3528 191156 3534
rect 191104 3470 191156 3476
rect 192024 3528 192076 3534
rect 192024 3470 192076 3476
rect 193864 3528 193916 3534
rect 193864 3470 193916 3476
rect 189816 3120 189868 3126
rect 189816 3062 189868 3068
rect 190828 3120 190880 3126
rect 190828 3062 190880 3068
rect 190840 480 190868 3062
rect 192036 480 192064 3470
rect 193220 3460 193272 3466
rect 193220 3402 193272 3408
rect 193232 480 193260 3402
rect 194428 480 194456 3878
rect 196636 3534 196664 17167
rect 197096 9042 197124 142802
rect 197188 17270 197216 152730
rect 197372 150414 197400 153870
rect 197648 153406 197676 160140
rect 197636 153400 197688 153406
rect 197636 153342 197688 153348
rect 197740 152674 197768 160140
rect 197556 152646 197768 152674
rect 197452 152448 197504 152454
rect 197452 152390 197504 152396
rect 197360 150408 197412 150414
rect 197360 150350 197412 150356
rect 197464 133822 197492 152390
rect 197556 139369 197584 152646
rect 197832 152454 197860 160140
rect 197924 159905 197952 160140
rect 197910 159896 197966 159905
rect 197910 159831 197966 159840
rect 197912 159792 197964 159798
rect 198016 159769 198044 160140
rect 197912 159734 197964 159740
rect 198002 159760 198058 159769
rect 197924 159497 197952 159734
rect 198002 159695 198058 159704
rect 197910 159488 197966 159497
rect 197910 159423 197966 159432
rect 197910 158400 197966 158409
rect 197910 158335 197966 158344
rect 197924 158137 197952 158335
rect 198004 158228 198056 158234
rect 198004 158170 198056 158176
rect 197910 158128 197966 158137
rect 197910 158063 197966 158072
rect 197910 155408 197966 155417
rect 197910 155343 197966 155352
rect 197924 155009 197952 155343
rect 198016 155310 198044 158170
rect 198004 155304 198056 155310
rect 198004 155246 198056 155252
rect 197910 155000 197966 155009
rect 197910 154935 197966 154944
rect 197912 154420 197964 154426
rect 197912 154362 197964 154368
rect 197820 152448 197872 152454
rect 197820 152390 197872 152396
rect 197636 152244 197688 152250
rect 197636 152186 197688 152192
rect 197648 140690 197676 152186
rect 197924 150113 197952 154362
rect 198004 153400 198056 153406
rect 198004 153342 198056 153348
rect 197910 150104 197966 150113
rect 197910 150039 197966 150048
rect 198016 145790 198044 153342
rect 198108 147674 198136 160140
rect 198200 157706 198228 160140
rect 198292 158681 198320 160140
rect 198278 158672 198334 158681
rect 198278 158607 198334 158616
rect 198384 158409 198412 160140
rect 198370 158400 198426 158409
rect 198370 158335 198426 158344
rect 198200 157678 198320 157706
rect 198292 157622 198320 157678
rect 198188 157616 198240 157622
rect 198188 157558 198240 157564
rect 198280 157616 198332 157622
rect 198280 157558 198332 157564
rect 198200 151094 198228 157558
rect 198476 156505 198504 160140
rect 198568 159905 198596 160140
rect 198554 159896 198610 159905
rect 198554 159831 198610 159840
rect 198556 159792 198608 159798
rect 198556 159734 198608 159740
rect 198568 158846 198596 159734
rect 198556 158840 198608 158846
rect 198556 158782 198608 158788
rect 198462 156496 198518 156505
rect 198462 156431 198518 156440
rect 198660 152250 198688 160140
rect 198752 157334 198780 160140
rect 198844 159905 198872 160140
rect 198830 159896 198886 159905
rect 198830 159831 198886 159840
rect 198844 157865 198872 159831
rect 198830 157856 198886 157865
rect 198830 157791 198886 157800
rect 198752 157306 198872 157334
rect 198740 152448 198792 152454
rect 198740 152390 198792 152396
rect 198648 152244 198700 152250
rect 198648 152186 198700 152192
rect 198188 151088 198240 151094
rect 198188 151030 198240 151036
rect 198108 147646 198596 147674
rect 198004 145784 198056 145790
rect 198004 145726 198056 145732
rect 197636 140684 197688 140690
rect 197636 140626 197688 140632
rect 197542 139360 197598 139369
rect 197542 139295 197598 139304
rect 197452 133816 197504 133822
rect 197452 133758 197504 133764
rect 198568 126886 198596 147646
rect 198646 139360 198702 139369
rect 198646 139295 198702 139304
rect 198556 126880 198608 126886
rect 198556 126822 198608 126828
rect 197358 116512 197414 116521
rect 197358 116447 197414 116456
rect 197176 17264 197228 17270
rect 197176 17206 197228 17212
rect 197372 16574 197400 116447
rect 198660 73846 198688 139295
rect 198752 125594 198780 152390
rect 198844 145722 198872 157306
rect 198936 148730 198964 160140
rect 199028 148889 199056 160140
rect 199120 159905 199148 160140
rect 199106 159896 199162 159905
rect 199106 159831 199162 159840
rect 199120 158001 199148 159831
rect 199212 158681 199240 160140
rect 199198 158672 199254 158681
rect 199198 158607 199254 158616
rect 199106 157992 199162 158001
rect 199106 157927 199162 157936
rect 199304 157826 199332 160140
rect 199396 159905 199424 160140
rect 199382 159896 199438 159905
rect 199382 159831 199438 159840
rect 199384 159792 199436 159798
rect 199382 159760 199384 159769
rect 199436 159760 199438 159769
rect 199382 159695 199438 159704
rect 199488 158794 199516 160140
rect 199396 158766 199516 158794
rect 199292 157820 199344 157826
rect 199292 157762 199344 157768
rect 199396 152454 199424 158766
rect 199476 157684 199528 157690
rect 199476 157626 199528 157632
rect 199384 152448 199436 152454
rect 199384 152390 199436 152396
rect 199014 148880 199070 148889
rect 199014 148815 199070 148824
rect 199488 148753 199516 157626
rect 199580 151201 199608 160140
rect 199672 159934 199700 160140
rect 199660 159928 199712 159934
rect 199660 159870 199712 159876
rect 199660 158840 199712 158846
rect 199660 158782 199712 158788
rect 199672 154737 199700 158782
rect 199658 154728 199714 154737
rect 199658 154663 199714 154672
rect 199566 151192 199622 151201
rect 199566 151127 199622 151136
rect 199474 148744 199530 148753
rect 198936 148702 199148 148730
rect 198832 145716 198884 145722
rect 198832 145658 198884 145664
rect 199120 144914 199148 148702
rect 199474 148679 199530 148688
rect 198936 144886 199148 144914
rect 198936 132394 198964 144886
rect 199764 142154 199792 160140
rect 199856 158681 199884 160140
rect 199842 158672 199898 158681
rect 199842 158607 199898 158616
rect 199948 158409 199976 160140
rect 200040 158710 200068 160140
rect 200132 159361 200160 160140
rect 200118 159352 200174 159361
rect 200118 159287 200174 159296
rect 200028 158704 200080 158710
rect 200224 158681 200252 160140
rect 200028 158646 200080 158652
rect 200210 158672 200266 158681
rect 200210 158607 200266 158616
rect 199934 158400 199990 158409
rect 199934 158335 199990 158344
rect 200316 158001 200344 160140
rect 200408 158953 200436 160140
rect 200394 158944 200450 158953
rect 200394 158879 200450 158888
rect 200026 157992 200082 158001
rect 200026 157927 200082 157936
rect 200302 157992 200358 158001
rect 200302 157927 200358 157936
rect 199934 157856 199990 157865
rect 199934 157791 199990 157800
rect 199842 154592 199898 154601
rect 199842 154527 199898 154536
rect 199672 142126 199792 142154
rect 198924 132388 198976 132394
rect 198924 132330 198976 132336
rect 199672 129674 199700 142126
rect 199660 129668 199712 129674
rect 199660 129610 199712 129616
rect 198740 125588 198792 125594
rect 198740 125530 198792 125536
rect 198648 73840 198700 73846
rect 198648 73782 198700 73788
rect 197372 16546 197952 16574
rect 197084 9036 197136 9042
rect 197084 8978 197136 8984
rect 195612 3528 195664 3534
rect 195612 3470 195664 3476
rect 196624 3528 196676 3534
rect 196624 3470 196676 3476
rect 195624 480 195652 3470
rect 196808 3392 196860 3398
rect 196808 3334 196860 3340
rect 196820 480 196848 3334
rect 197924 480 197952 16546
rect 199856 6186 199884 154527
rect 199844 6180 199896 6186
rect 199844 6122 199896 6128
rect 199948 3534 199976 157791
rect 199108 3528 199160 3534
rect 199108 3470 199160 3476
rect 199936 3528 199988 3534
rect 199936 3470 199988 3476
rect 199120 480 199148 3470
rect 200040 3466 200068 157927
rect 200212 157888 200264 157894
rect 200212 157830 200264 157836
rect 200120 157820 200172 157826
rect 200120 157762 200172 157768
rect 200132 156194 200160 157762
rect 200224 157690 200252 157830
rect 200212 157684 200264 157690
rect 200212 157626 200264 157632
rect 200500 157334 200528 160140
rect 200224 157306 200528 157334
rect 200120 156188 200172 156194
rect 200120 156130 200172 156136
rect 200120 152448 200172 152454
rect 200120 152390 200172 152396
rect 200132 128314 200160 152390
rect 200224 144129 200252 157306
rect 200302 152552 200358 152561
rect 200302 152487 200358 152496
rect 200316 152289 200344 152487
rect 200592 152454 200620 160140
rect 200684 159934 200712 160140
rect 200672 159928 200724 159934
rect 200672 159870 200724 159876
rect 200672 159180 200724 159186
rect 200672 159122 200724 159128
rect 200684 158846 200712 159122
rect 200672 158840 200724 158846
rect 200672 158782 200724 158788
rect 200672 158024 200724 158030
rect 200672 157966 200724 157972
rect 200684 157321 200712 157966
rect 200670 157312 200726 157321
rect 200670 157247 200726 157256
rect 200580 152448 200632 152454
rect 200580 152390 200632 152396
rect 200302 152280 200358 152289
rect 200302 152215 200358 152224
rect 200776 147674 200804 160140
rect 200868 156913 200896 160140
rect 200960 158681 200988 160140
rect 200946 158672 201002 158681
rect 200946 158607 201002 158616
rect 201052 158409 201080 160140
rect 201038 158400 201094 158409
rect 200948 158364 201000 158370
rect 201038 158335 201094 158344
rect 200948 158306 201000 158312
rect 200960 157554 200988 158306
rect 200948 157548 201000 157554
rect 200948 157490 201000 157496
rect 200854 156904 200910 156913
rect 200854 156839 200910 156848
rect 201038 156904 201094 156913
rect 201038 156839 201094 156848
rect 200856 156800 200908 156806
rect 200856 156742 200908 156748
rect 200868 156330 200896 156742
rect 200856 156324 200908 156330
rect 200856 156266 200908 156272
rect 200948 156188 201000 156194
rect 200948 156130 201000 156136
rect 200856 154488 200908 154494
rect 200856 154430 200908 154436
rect 200868 149938 200896 154430
rect 200856 149932 200908 149938
rect 200856 149874 200908 149880
rect 200868 148102 200896 149874
rect 200856 148096 200908 148102
rect 200856 148038 200908 148044
rect 200960 147674 200988 156130
rect 201052 150249 201080 156839
rect 201144 151609 201172 160140
rect 201236 158030 201264 160140
rect 201328 159905 201356 160140
rect 201314 159896 201370 159905
rect 201314 159831 201370 159840
rect 201316 159316 201368 159322
rect 201316 159258 201368 159264
rect 201328 159186 201356 159258
rect 201316 159180 201368 159186
rect 201316 159122 201368 159128
rect 201420 159089 201448 160140
rect 201406 159080 201462 159089
rect 201406 159015 201462 159024
rect 201512 158817 201540 160140
rect 201498 158808 201554 158817
rect 201498 158743 201554 158752
rect 201316 158568 201368 158574
rect 201316 158510 201368 158516
rect 201224 158024 201276 158030
rect 201224 157966 201276 157972
rect 201328 157706 201356 158510
rect 201406 158400 201462 158409
rect 201406 158335 201462 158344
rect 201236 157678 201356 157706
rect 201130 151600 201186 151609
rect 201130 151535 201186 151544
rect 201236 151026 201264 157678
rect 201314 157448 201370 157457
rect 201314 157383 201370 157392
rect 201224 151020 201276 151026
rect 201224 150962 201276 150968
rect 201038 150240 201094 150249
rect 201038 150175 201094 150184
rect 200316 147646 200804 147674
rect 200868 147646 200988 147674
rect 200316 144294 200344 147646
rect 200868 145586 200896 147646
rect 200856 145580 200908 145586
rect 200856 145522 200908 145528
rect 201132 144628 201184 144634
rect 201132 144570 201184 144576
rect 200304 144288 200356 144294
rect 200304 144230 200356 144236
rect 201144 144242 201172 144570
rect 201224 144560 201276 144566
rect 201224 144502 201276 144508
rect 201236 144401 201264 144502
rect 201222 144392 201278 144401
rect 201222 144327 201278 144336
rect 201224 144288 201276 144294
rect 201144 144236 201224 144242
rect 201144 144230 201276 144236
rect 201144 144214 201264 144230
rect 200210 144120 200266 144129
rect 200210 144055 200266 144064
rect 201130 144120 201186 144129
rect 201130 144055 201186 144064
rect 200120 128308 200172 128314
rect 200120 128250 200172 128256
rect 201144 109750 201172 144055
rect 201132 109744 201184 109750
rect 201132 109686 201184 109692
rect 201236 108322 201264 144214
rect 201224 108316 201276 108322
rect 201224 108258 201276 108264
rect 201328 35222 201356 157383
rect 201420 148986 201448 158335
rect 201500 155780 201552 155786
rect 201500 155722 201552 155728
rect 201512 150346 201540 155722
rect 201500 150340 201552 150346
rect 201500 150282 201552 150288
rect 201408 148980 201460 148986
rect 201408 148922 201460 148928
rect 201408 148096 201460 148102
rect 201408 148038 201460 148044
rect 201316 35216 201368 35222
rect 201316 35158 201368 35164
rect 200304 3664 200356 3670
rect 200304 3606 200356 3612
rect 200028 3460 200080 3466
rect 200028 3402 200080 3408
rect 200316 480 200344 3606
rect 201420 2990 201448 148038
rect 201408 2984 201460 2990
rect 201408 2926 201460 2932
rect 201512 480 201540 150282
rect 201604 124098 201632 160140
rect 201696 154873 201724 160140
rect 201788 158438 201816 160140
rect 201776 158432 201828 158438
rect 201776 158374 201828 158380
rect 201880 156097 201908 160140
rect 201866 156088 201922 156097
rect 201866 156023 201922 156032
rect 201682 154864 201738 154873
rect 201682 154799 201738 154808
rect 201684 152448 201736 152454
rect 201684 152390 201736 152396
rect 201696 146266 201724 152390
rect 201776 152244 201828 152250
rect 201776 152186 201828 152192
rect 201684 146260 201736 146266
rect 201684 146202 201736 146208
rect 201788 146198 201816 152186
rect 201972 147626 202000 160140
rect 202064 154426 202092 160140
rect 202156 158409 202184 160140
rect 202142 158400 202198 158409
rect 202142 158335 202198 158344
rect 202144 155168 202196 155174
rect 202144 155110 202196 155116
rect 202052 154420 202104 154426
rect 202052 154362 202104 154368
rect 202156 147674 202184 155110
rect 202248 153202 202276 160140
rect 202340 159905 202368 160140
rect 202326 159896 202382 159905
rect 202326 159831 202382 159840
rect 202326 159488 202382 159497
rect 202326 159423 202382 159432
rect 202340 159186 202368 159423
rect 202328 159180 202380 159186
rect 202328 159122 202380 159128
rect 202328 158704 202380 158710
rect 202432 158681 202460 160140
rect 202328 158646 202380 158652
rect 202418 158672 202474 158681
rect 202236 153196 202288 153202
rect 202236 153138 202288 153144
rect 202340 148918 202368 158646
rect 202418 158607 202474 158616
rect 202524 152454 202552 160140
rect 202616 155446 202644 160140
rect 202708 158001 202736 160140
rect 202694 157992 202750 158001
rect 202694 157927 202750 157936
rect 202604 155440 202656 155446
rect 202604 155382 202656 155388
rect 202694 154864 202750 154873
rect 202694 154799 202750 154808
rect 202604 153196 202656 153202
rect 202604 153138 202656 153144
rect 202616 152454 202644 153138
rect 202512 152448 202564 152454
rect 202512 152390 202564 152396
rect 202604 152448 202656 152454
rect 202604 152390 202656 152396
rect 202328 148912 202380 148918
rect 202328 148854 202380 148860
rect 202708 147674 202736 154799
rect 202800 152250 202828 160140
rect 202892 159497 202920 160140
rect 202878 159488 202934 159497
rect 202878 159423 202934 159432
rect 202880 158704 202932 158710
rect 202984 158681 203012 160140
rect 202880 158646 202932 158652
rect 202970 158672 203026 158681
rect 202892 155553 202920 158646
rect 202970 158607 203026 158616
rect 203076 155854 203104 160140
rect 203064 155848 203116 155854
rect 203064 155790 203116 155796
rect 202878 155544 202934 155553
rect 202878 155479 202934 155488
rect 203168 154465 203196 160140
rect 203154 154456 203210 154465
rect 203154 154391 203210 154400
rect 202880 153808 202932 153814
rect 202880 153750 202932 153756
rect 202788 152244 202840 152250
rect 202788 152186 202840 152192
rect 202892 149054 202920 153750
rect 202880 149048 202932 149054
rect 202880 148990 202932 148996
rect 203260 147674 203288 160140
rect 203352 158710 203380 160140
rect 203444 159769 203472 160140
rect 203536 159905 203564 160140
rect 203522 159896 203578 159905
rect 203522 159831 203578 159840
rect 203524 159792 203576 159798
rect 203430 159760 203486 159769
rect 203524 159734 203576 159740
rect 203430 159695 203486 159704
rect 203432 159180 203484 159186
rect 203432 159122 203484 159128
rect 203340 158704 203392 158710
rect 203340 158646 203392 158652
rect 203444 154986 203472 159122
rect 203536 158642 203564 159734
rect 203524 158636 203576 158642
rect 203524 158578 203576 158584
rect 203628 155174 203656 160140
rect 203720 158506 203748 160140
rect 203812 159905 203840 160140
rect 203798 159896 203854 159905
rect 203798 159831 203854 159840
rect 203800 159792 203852 159798
rect 203800 159734 203852 159740
rect 203812 159254 203840 159734
rect 203800 159248 203852 159254
rect 203800 159190 203852 159196
rect 203800 158636 203852 158642
rect 203800 158578 203852 158584
rect 203708 158500 203760 158506
rect 203708 158442 203760 158448
rect 203616 155168 203668 155174
rect 203616 155110 203668 155116
rect 203444 154958 203748 154986
rect 203614 154728 203670 154737
rect 203614 154663 203670 154672
rect 202156 147646 202276 147674
rect 202708 147646 202828 147674
rect 201960 147620 202012 147626
rect 201960 147562 202012 147568
rect 202248 146742 202276 147646
rect 202236 146736 202288 146742
rect 202236 146678 202288 146684
rect 201776 146192 201828 146198
rect 201776 146134 201828 146140
rect 202694 144392 202750 144401
rect 202694 144327 202750 144336
rect 202708 144226 202736 144327
rect 202696 144220 202748 144226
rect 202696 144162 202748 144168
rect 201592 124092 201644 124098
rect 201592 124034 201644 124040
rect 201592 105664 201644 105670
rect 201592 105606 201644 105612
rect 201604 16574 201632 105606
rect 202708 101454 202736 144162
rect 202696 101448 202748 101454
rect 202696 101390 202748 101396
rect 201604 16546 202736 16574
rect 202708 480 202736 16546
rect 202800 15910 202828 147646
rect 202892 147646 203288 147674
rect 202892 144906 202920 147646
rect 202880 144900 202932 144906
rect 202880 144842 202932 144848
rect 203628 143410 203656 154663
rect 203720 146810 203748 154958
rect 203812 151745 203840 158578
rect 203798 151736 203854 151745
rect 203798 151671 203854 151680
rect 203708 146804 203760 146810
rect 203708 146746 203760 146752
rect 203904 144702 203932 160140
rect 203996 158681 204024 160140
rect 204088 159769 204116 160140
rect 204074 159760 204130 159769
rect 204074 159695 204130 159704
rect 203982 158672 204038 158681
rect 203982 158607 204038 158616
rect 204088 157334 204116 159695
rect 204180 158642 204208 160140
rect 204168 158636 204220 158642
rect 204168 158578 204220 158584
rect 204272 158574 204300 160140
rect 204364 158681 204392 160140
rect 204350 158672 204406 158681
rect 204350 158607 204406 158616
rect 204260 158568 204312 158574
rect 204260 158510 204312 158516
rect 204258 158400 204314 158409
rect 204258 158335 204314 158344
rect 204168 157752 204220 157758
rect 204168 157694 204220 157700
rect 204180 157350 204208 157694
rect 203996 157306 204116 157334
rect 204168 157344 204220 157350
rect 203892 144696 203944 144702
rect 203892 144638 203944 144644
rect 203706 144392 203762 144401
rect 203706 144327 203762 144336
rect 203720 143993 203748 144327
rect 203706 143984 203762 143993
rect 203706 143919 203762 143928
rect 203616 143404 203668 143410
rect 203616 143346 203668 143352
rect 203996 94518 204024 157306
rect 204168 157286 204220 157292
rect 204166 155544 204222 155553
rect 204166 155479 204222 155488
rect 204076 155168 204128 155174
rect 204076 155110 204128 155116
rect 204088 150385 204116 155110
rect 204074 150376 204130 150385
rect 204074 150311 204130 150320
rect 204076 144900 204128 144906
rect 204076 144842 204128 144848
rect 204088 144294 204116 144842
rect 204076 144288 204128 144294
rect 204076 144230 204128 144236
rect 203984 94512 204036 94518
rect 203984 94454 204036 94460
rect 204088 33794 204116 144230
rect 204180 37942 204208 155479
rect 204168 37936 204220 37942
rect 204168 37878 204220 37884
rect 204076 33788 204128 33794
rect 204076 33730 204128 33736
rect 202788 15904 202840 15910
rect 202788 15846 202840 15852
rect 204272 7614 204300 158335
rect 204456 157434 204484 160140
rect 204548 159254 204576 160140
rect 204640 159905 204668 160140
rect 204626 159896 204682 159905
rect 204626 159831 204682 159840
rect 204536 159248 204588 159254
rect 204536 159190 204588 159196
rect 204456 157406 204576 157434
rect 204548 155281 204576 157406
rect 204534 155272 204590 155281
rect 204534 155207 204590 155216
rect 204732 149025 204760 160140
rect 204824 158642 204852 160140
rect 204916 159089 204944 160140
rect 204902 159080 204958 159089
rect 204902 159015 204958 159024
rect 204812 158636 204864 158642
rect 204812 158578 204864 158584
rect 204718 149016 204774 149025
rect 204718 148951 204774 148960
rect 205008 147674 205036 160140
rect 205100 159338 205128 160140
rect 205192 159905 205220 160140
rect 205178 159896 205234 159905
rect 205178 159831 205234 159840
rect 205100 159310 205220 159338
rect 205088 159180 205140 159186
rect 205088 159122 205140 159128
rect 204364 147646 205036 147674
rect 204364 141982 204392 147646
rect 204352 141976 204404 141982
rect 204352 141918 204404 141924
rect 204718 139360 204774 139369
rect 204718 139295 204774 139304
rect 204732 139210 204760 139295
rect 205100 139262 205128 159122
rect 205192 158409 205220 159310
rect 205178 158400 205234 158409
rect 205178 158335 205234 158344
rect 205180 157888 205232 157894
rect 205180 157830 205232 157836
rect 205192 151337 205220 157830
rect 205284 153134 205312 160140
rect 205376 154329 205404 160140
rect 205468 159769 205496 160140
rect 205454 159760 205510 159769
rect 205454 159695 205510 159704
rect 205468 157334 205496 159695
rect 205560 159186 205588 160140
rect 205652 159769 205680 160140
rect 205638 159760 205694 159769
rect 205638 159695 205694 159704
rect 205548 159180 205600 159186
rect 205548 159122 205600 159128
rect 205468 157306 205588 157334
rect 205454 155272 205510 155281
rect 205454 155207 205510 155216
rect 205362 154320 205418 154329
rect 205362 154255 205418 154264
rect 205272 153128 205324 153134
rect 205272 153070 205324 153076
rect 205178 151328 205234 151337
rect 205178 151263 205234 151272
rect 205088 139256 205140 139262
rect 204994 139224 205050 139233
rect 204732 139182 204994 139210
rect 205088 139198 205140 139204
rect 204994 139159 205050 139168
rect 205468 18630 205496 155207
rect 205560 91798 205588 157306
rect 205744 153270 205772 160140
rect 205836 154494 205864 160140
rect 205928 159866 205956 160140
rect 205916 159860 205968 159866
rect 205916 159802 205968 159808
rect 206020 157334 206048 160140
rect 205928 157306 206048 157334
rect 205824 154488 205876 154494
rect 205824 154430 205876 154436
rect 205732 153264 205784 153270
rect 205732 153206 205784 153212
rect 205640 153196 205692 153202
rect 205928 153184 205956 157306
rect 206008 153264 206060 153270
rect 206008 153206 206060 153212
rect 205640 153138 205692 153144
rect 205836 153156 205956 153184
rect 205652 152538 205680 153138
rect 205652 152510 205772 152538
rect 205640 152040 205692 152046
rect 205640 151982 205692 151988
rect 205652 136542 205680 151982
rect 205744 137902 205772 152510
rect 205836 141710 205864 153156
rect 205916 152312 205968 152318
rect 205916 152254 205968 152260
rect 205824 141704 205876 141710
rect 205824 141646 205876 141652
rect 205836 140826 205864 141646
rect 205928 140894 205956 152254
rect 206020 149122 206048 153206
rect 206008 149116 206060 149122
rect 206008 149058 206060 149064
rect 206112 147490 206140 160140
rect 206204 159089 206232 160140
rect 206296 159905 206324 160140
rect 206282 159896 206338 159905
rect 206282 159831 206338 159840
rect 206190 159080 206246 159089
rect 206190 159015 206246 159024
rect 206192 153264 206244 153270
rect 206192 153206 206244 153212
rect 206204 152318 206232 153206
rect 206296 152402 206324 159831
rect 206388 153202 206416 160140
rect 206480 159934 206508 160140
rect 206468 159928 206520 159934
rect 206572 159905 206600 160140
rect 206468 159870 206520 159876
rect 206558 159896 206614 159905
rect 206558 159831 206614 159840
rect 206376 153196 206428 153202
rect 206376 153138 206428 153144
rect 206572 152538 206600 159831
rect 206664 153270 206692 160140
rect 206756 159934 206784 160140
rect 206744 159928 206796 159934
rect 206848 159905 206876 160140
rect 206744 159870 206796 159876
rect 206834 159896 206890 159905
rect 206834 159831 206890 159840
rect 206744 159180 206796 159186
rect 206744 159122 206796 159128
rect 206756 158710 206784 159122
rect 206744 158704 206796 158710
rect 206744 158646 206796 158652
rect 206652 153264 206704 153270
rect 206652 153206 206704 153212
rect 206572 152510 206784 152538
rect 206296 152374 206692 152402
rect 206192 152312 206244 152318
rect 206192 152254 206244 152260
rect 206560 149116 206612 149122
rect 206560 149058 206612 149064
rect 206572 147665 206600 149058
rect 206558 147656 206614 147665
rect 206558 147591 206614 147600
rect 206100 147484 206152 147490
rect 206100 147426 206152 147432
rect 205916 140888 205968 140894
rect 205916 140830 205968 140836
rect 205824 140820 205876 140826
rect 205824 140762 205876 140768
rect 206468 140820 206520 140826
rect 206468 140762 206520 140768
rect 205732 137896 205784 137902
rect 205732 137838 205784 137844
rect 205640 136536 205692 136542
rect 205640 136478 205692 136484
rect 205548 91792 205600 91798
rect 205548 91734 205600 91740
rect 206480 89010 206508 140762
rect 206572 90370 206600 147591
rect 206560 90364 206612 90370
rect 206560 90306 206612 90312
rect 206468 89004 206520 89010
rect 206468 88946 206520 88952
rect 206664 87650 206692 152374
rect 206652 87644 206704 87650
rect 206652 87586 206704 87592
rect 206756 86290 206784 152510
rect 205640 86284 205692 86290
rect 205640 86226 205692 86232
rect 206744 86284 206796 86290
rect 206744 86226 206796 86232
rect 205456 18624 205508 18630
rect 205456 18566 205508 18572
rect 205652 16574 205680 86226
rect 206848 84862 206876 159831
rect 206940 152046 206968 160140
rect 207032 158681 207060 160140
rect 207018 158672 207074 158681
rect 207018 158607 207074 158616
rect 207020 158160 207072 158166
rect 207124 158137 207152 160140
rect 207216 158794 207244 160140
rect 207308 159905 207336 160140
rect 207294 159896 207350 159905
rect 207294 159831 207350 159840
rect 207400 159769 207428 160140
rect 207386 159760 207442 159769
rect 207386 159695 207442 159704
rect 207216 158766 207336 158794
rect 207204 158704 207256 158710
rect 207204 158646 207256 158652
rect 207020 158102 207072 158108
rect 207110 158128 207166 158137
rect 207032 156602 207060 158102
rect 207110 158063 207166 158072
rect 207112 157956 207164 157962
rect 207112 157898 207164 157904
rect 207020 156596 207072 156602
rect 207020 156538 207072 156544
rect 207124 154902 207152 157898
rect 207216 157350 207244 158646
rect 207308 157729 207336 158766
rect 207400 157865 207428 159695
rect 207492 159186 207520 161094
rect 207480 159180 207532 159186
rect 207480 159122 207532 159128
rect 207584 158522 207612 170303
rect 207676 166274 207704 238546
rect 207860 237114 207888 238726
rect 207848 237108 207900 237114
rect 207848 237050 207900 237056
rect 207756 236020 207808 236026
rect 207756 235962 207808 235968
rect 207768 227186 207796 235962
rect 207860 229022 207888 237050
rect 208044 237046 208072 319359
rect 208216 318980 208268 318986
rect 208216 318922 208268 318928
rect 208124 311432 208176 311438
rect 208124 311374 208176 311380
rect 208032 237040 208084 237046
rect 208032 236982 208084 236988
rect 208044 236026 208072 236982
rect 208032 236020 208084 236026
rect 208032 235962 208084 235968
rect 207848 229016 207900 229022
rect 207848 228958 207900 228964
rect 208136 228954 208164 311374
rect 208228 229090 208256 318922
rect 209596 317076 209648 317082
rect 209596 317018 209648 317024
rect 209044 316940 209096 316946
rect 209044 316882 209096 316888
rect 208308 314696 208360 314702
rect 208308 314638 208360 314644
rect 208216 229084 208268 229090
rect 208216 229026 208268 229032
rect 208124 228948 208176 228954
rect 208124 228890 208176 228896
rect 208228 228886 208256 229026
rect 208216 228880 208268 228886
rect 208216 228822 208268 228828
rect 207756 227180 207808 227186
rect 207756 227122 207808 227128
rect 208320 224369 208348 314638
rect 209056 241534 209084 316882
rect 209504 312792 209556 312798
rect 209504 312734 209556 312740
rect 209412 307080 209464 307086
rect 209412 307022 209464 307028
rect 209228 305176 209280 305182
rect 209228 305118 209280 305124
rect 209044 241528 209096 241534
rect 209044 241470 209096 241476
rect 209056 238754 209084 241470
rect 208964 238726 209084 238754
rect 208964 238241 208992 238726
rect 209044 238536 209096 238542
rect 209044 238478 209096 238484
rect 208950 238232 209006 238241
rect 208950 238167 209006 238176
rect 208860 237788 208912 237794
rect 208860 237730 208912 237736
rect 208400 237244 208452 237250
rect 208400 237186 208452 237192
rect 208412 233918 208440 237186
rect 208766 234560 208822 234569
rect 208766 234495 208822 234504
rect 208492 234456 208544 234462
rect 208492 234398 208544 234404
rect 208400 233912 208452 233918
rect 208400 233854 208452 233860
rect 208504 233753 208532 234398
rect 208490 233744 208546 233753
rect 208490 233679 208546 233688
rect 208780 233617 208808 234495
rect 208766 233608 208822 233617
rect 208766 233543 208822 233552
rect 208306 224360 208362 224369
rect 208306 224295 208362 224304
rect 207754 202192 207810 202201
rect 207754 202127 207810 202136
rect 207768 166433 207796 202127
rect 207846 188320 207902 188329
rect 207846 188255 207902 188264
rect 207754 166424 207810 166433
rect 207754 166359 207810 166368
rect 207676 166246 207796 166274
rect 207662 166152 207718 166161
rect 207662 166087 207718 166096
rect 207676 159866 207704 166087
rect 207664 159860 207716 159866
rect 207664 159802 207716 159808
rect 207768 159730 207796 166246
rect 207756 159724 207808 159730
rect 207756 159666 207808 159672
rect 207756 159180 207808 159186
rect 207756 159122 207808 159128
rect 207584 158494 207704 158522
rect 207480 158296 207532 158302
rect 207676 158273 207704 158494
rect 207480 158238 207532 158244
rect 207662 158264 207718 158273
rect 207386 157856 207442 157865
rect 207386 157791 207442 157800
rect 207294 157720 207350 157729
rect 207294 157655 207350 157664
rect 207296 157480 207348 157486
rect 207296 157422 207348 157428
rect 207204 157344 207256 157350
rect 207204 157286 207256 157292
rect 207204 155780 207256 155786
rect 207204 155722 207256 155728
rect 207112 154896 207164 154902
rect 207112 154838 207164 154844
rect 206928 152040 206980 152046
rect 206928 151982 206980 151988
rect 207216 142154 207244 155722
rect 207308 153610 207336 157422
rect 207492 155825 207520 158238
rect 207572 158228 207624 158234
rect 207662 158199 207718 158208
rect 207572 158170 207624 158176
rect 207478 155816 207534 155825
rect 207478 155751 207534 155760
rect 207584 154562 207612 158170
rect 207768 157978 207796 159122
rect 207860 158098 207888 188255
rect 207938 184240 207994 184249
rect 207938 184175 207994 184184
rect 207952 161226 207980 184175
rect 208766 173632 208822 173641
rect 208766 173567 208822 173576
rect 208030 173496 208086 173505
rect 208030 173431 208086 173440
rect 207940 161220 207992 161226
rect 207940 161162 207992 161168
rect 207940 161084 207992 161090
rect 207940 161026 207992 161032
rect 207952 160138 207980 161026
rect 207940 160132 207992 160138
rect 207940 160074 207992 160080
rect 207848 158092 207900 158098
rect 207848 158034 207900 158040
rect 207940 158092 207992 158098
rect 207940 158034 207992 158040
rect 207768 157950 207888 157978
rect 207756 156732 207808 156738
rect 207756 156674 207808 156680
rect 207768 155786 207796 156674
rect 207756 155780 207808 155786
rect 207756 155722 207808 155728
rect 207572 154556 207624 154562
rect 207572 154498 207624 154504
rect 207296 153604 207348 153610
rect 207296 153546 207348 153552
rect 207860 152658 207888 157950
rect 207952 157418 207980 158034
rect 208044 157894 208072 173431
rect 208122 166424 208178 166433
rect 208122 166359 208178 166368
rect 208032 157888 208084 157894
rect 208032 157830 208084 157836
rect 208136 157826 208164 166359
rect 208400 161424 208452 161430
rect 208214 161392 208270 161401
rect 208400 161366 208452 161372
rect 208214 161327 208270 161336
rect 208228 160313 208256 161327
rect 208308 161220 208360 161226
rect 208308 161162 208360 161168
rect 208214 160304 208270 160313
rect 208214 160239 208270 160248
rect 208214 158128 208270 158137
rect 208320 158098 208348 161162
rect 208412 160954 208440 161366
rect 208400 160948 208452 160954
rect 208400 160890 208452 160896
rect 208398 160712 208454 160721
rect 208398 160647 208454 160656
rect 208412 160177 208440 160647
rect 208398 160168 208454 160177
rect 208398 160103 208454 160112
rect 208780 159934 208808 173567
rect 208768 159928 208820 159934
rect 208768 159870 208820 159876
rect 208584 159656 208636 159662
rect 208584 159598 208636 159604
rect 208214 158063 208270 158072
rect 208308 158092 208360 158098
rect 208124 157820 208176 157826
rect 208124 157762 208176 157768
rect 208122 157720 208178 157729
rect 208122 157655 208178 157664
rect 207940 157412 207992 157418
rect 207940 157354 207992 157360
rect 207848 152652 207900 152658
rect 207848 152594 207900 152600
rect 207032 142126 207244 142154
rect 206928 141432 206980 141438
rect 206928 141374 206980 141380
rect 206940 140894 206968 141374
rect 206928 140888 206980 140894
rect 206928 140830 206980 140836
rect 206836 84856 206888 84862
rect 206836 84798 206888 84804
rect 206940 36582 206968 140830
rect 206928 36576 206980 36582
rect 206928 36518 206980 36524
rect 205652 16546 206232 16574
rect 204260 7608 204312 7614
rect 204260 7550 204312 7556
rect 203892 3800 203944 3806
rect 203892 3742 203944 3748
rect 203904 480 203932 3742
rect 205088 2984 205140 2990
rect 205088 2926 205140 2932
rect 205100 480 205128 2926
rect 206204 480 206232 16546
rect 187302 354 187414 480
rect 186884 326 187414 354
rect 187302 -960 187414 326
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207032 354 207060 142126
rect 208136 134570 208164 157655
rect 208124 134564 208176 134570
rect 208124 134506 208176 134512
rect 208228 83502 208256 158063
rect 208308 158034 208360 158040
rect 208400 158092 208452 158098
rect 208400 158034 208452 158040
rect 208306 157856 208362 157865
rect 208306 157791 208362 157800
rect 208216 83496 208268 83502
rect 208216 83438 208268 83444
rect 208320 80714 208348 157791
rect 208412 155961 208440 158034
rect 208490 157992 208546 158001
rect 208490 157927 208546 157936
rect 208398 155952 208454 155961
rect 208398 155887 208454 155896
rect 208400 153876 208452 153882
rect 208400 153818 208452 153824
rect 208308 80708 208360 80714
rect 208308 80650 208360 80656
rect 208412 16574 208440 153818
rect 208504 153649 208532 157927
rect 208596 157282 208624 159598
rect 208872 159322 208900 237730
rect 208952 202156 209004 202162
rect 208952 202098 209004 202104
rect 208964 160002 208992 202098
rect 208952 159996 209004 160002
rect 208952 159938 209004 159944
rect 209056 159798 209084 238478
rect 209136 238468 209188 238474
rect 209136 238410 209188 238416
rect 209044 159792 209096 159798
rect 209044 159734 209096 159740
rect 209148 159633 209176 238410
rect 209240 237250 209268 305118
rect 209318 304736 209374 304745
rect 209318 304671 209374 304680
rect 209228 237244 209280 237250
rect 209228 237186 209280 237192
rect 209332 234462 209360 304671
rect 209424 234569 209452 307022
rect 209516 236638 209544 312734
rect 209608 240825 209636 317018
rect 209688 315376 209740 315382
rect 209688 315318 209740 315324
rect 209594 240816 209650 240825
rect 209594 240751 209650 240760
rect 209504 236632 209556 236638
rect 209504 236574 209556 236580
rect 209700 235657 209728 315318
rect 210884 312724 210936 312730
rect 210884 312666 210936 312672
rect 210608 307828 210660 307834
rect 210608 307770 210660 307776
rect 210146 307048 210202 307057
rect 210146 306983 210202 306992
rect 209686 235648 209742 235657
rect 209686 235583 209742 235592
rect 209410 234560 209466 234569
rect 209410 234495 209466 234504
rect 209320 234456 209372 234462
rect 210160 234433 210188 306983
rect 210332 305924 210384 305930
rect 210332 305866 210384 305872
rect 210344 239737 210372 305866
rect 210516 295996 210568 296002
rect 210516 295938 210568 295944
rect 210424 241188 210476 241194
rect 210424 241130 210476 241136
rect 210330 239728 210386 239737
rect 210330 239663 210386 239672
rect 210240 238196 210292 238202
rect 210240 238138 210292 238144
rect 209320 234398 209372 234404
rect 210146 234424 210202 234433
rect 210146 234359 210202 234368
rect 209320 207732 209372 207738
rect 209320 207674 209372 207680
rect 209228 175976 209280 175982
rect 209228 175918 209280 175924
rect 209240 173641 209268 175918
rect 209226 173632 209282 173641
rect 209226 173567 209282 173576
rect 209228 161016 209280 161022
rect 209228 160958 209280 160964
rect 209240 160274 209268 160958
rect 209228 160268 209280 160274
rect 209228 160210 209280 160216
rect 209134 159624 209190 159633
rect 209134 159559 209190 159568
rect 208860 159316 208912 159322
rect 208860 159258 208912 159264
rect 209240 159186 209268 160210
rect 209228 159180 209280 159186
rect 209228 159122 209280 159128
rect 209332 158574 209360 207674
rect 209412 207664 209464 207670
rect 209412 207606 209464 207612
rect 209320 158568 209372 158574
rect 209320 158510 209372 158516
rect 209424 158409 209452 207606
rect 209596 206372 209648 206378
rect 209596 206314 209648 206320
rect 209504 206304 209556 206310
rect 209504 206246 209556 206252
rect 209516 158642 209544 206246
rect 209608 160206 209636 206314
rect 209688 205012 209740 205018
rect 209688 204954 209740 204960
rect 209596 160200 209648 160206
rect 209596 160142 209648 160148
rect 209504 158636 209556 158642
rect 209504 158578 209556 158584
rect 209700 158438 209728 204954
rect 210252 159390 210280 238138
rect 210332 180124 210384 180130
rect 210332 180066 210384 180072
rect 210240 159384 210292 159390
rect 210240 159326 210292 159332
rect 209688 158432 209740 158438
rect 209410 158400 209466 158409
rect 209688 158374 209740 158380
rect 209410 158335 209466 158344
rect 209688 158024 209740 158030
rect 209688 157966 209740 157972
rect 208584 157276 208636 157282
rect 208584 157218 208636 157224
rect 209504 156664 209556 156670
rect 209504 156606 209556 156612
rect 208490 153640 208546 153649
rect 208490 153575 208546 153584
rect 209516 147674 209544 156606
rect 209596 153876 209648 153882
rect 209596 153818 209648 153824
rect 209608 152946 209636 153818
rect 209700 153066 209728 157966
rect 210344 157593 210372 180066
rect 210330 157584 210386 157593
rect 210330 157519 210386 157528
rect 210436 157334 210464 241130
rect 210528 214742 210556 295938
rect 210620 238338 210648 307770
rect 210700 292664 210752 292670
rect 210700 292606 210752 292612
rect 210608 238332 210660 238338
rect 210608 238274 210660 238280
rect 210620 237930 210648 238274
rect 210608 237924 210660 237930
rect 210608 237866 210660 237872
rect 210608 234932 210660 234938
rect 210608 234874 210660 234880
rect 210516 214736 210568 214742
rect 210516 214678 210568 214684
rect 210516 200796 210568 200802
rect 210516 200738 210568 200744
rect 210528 158137 210556 200738
rect 210514 158128 210570 158137
rect 210514 158063 210570 158072
rect 210344 157306 210464 157334
rect 210344 155378 210372 157306
rect 210620 155922 210648 234874
rect 210712 213450 210740 292606
rect 210790 239728 210846 239737
rect 210790 239663 210846 239672
rect 210804 239329 210832 239663
rect 210790 239320 210846 239329
rect 210790 239255 210846 239264
rect 210896 235958 210924 312666
rect 210988 236609 211016 320719
rect 217876 320544 217928 320550
rect 217876 320486 217928 320492
rect 215022 319968 215078 319977
rect 215022 319903 215078 319912
rect 213090 319696 213146 319705
rect 213090 319631 213146 319640
rect 211068 319456 211120 319462
rect 211068 319398 211120 319404
rect 210974 236600 211030 236609
rect 210974 236535 211030 236544
rect 210884 235952 210936 235958
rect 210884 235894 210936 235900
rect 210792 234728 210844 234734
rect 210792 234670 210844 234676
rect 210700 213444 210752 213450
rect 210700 213386 210752 213392
rect 210700 199436 210752 199442
rect 210700 199378 210752 199384
rect 210712 158370 210740 199378
rect 210700 158364 210752 158370
rect 210700 158306 210752 158312
rect 210804 156505 210832 234670
rect 210884 228948 210936 228954
rect 210884 228890 210936 228896
rect 210790 156496 210846 156505
rect 210790 156431 210846 156440
rect 210608 155916 210660 155922
rect 210608 155858 210660 155864
rect 210422 155680 210478 155689
rect 210422 155615 210478 155624
rect 210332 155372 210384 155378
rect 210332 155314 210384 155320
rect 209688 153060 209740 153066
rect 209688 153002 209740 153008
rect 209780 153060 209832 153066
rect 209780 153002 209832 153008
rect 209792 152946 209820 153002
rect 209608 152918 209820 152946
rect 209872 152312 209924 152318
rect 209872 152254 209924 152260
rect 209884 152114 209912 152254
rect 209872 152108 209924 152114
rect 209872 152050 209924 152056
rect 209516 147646 209728 147674
rect 208412 16546 208624 16574
rect 208596 480 208624 16546
rect 209700 4146 209728 147646
rect 209884 6914 209912 152050
rect 210344 147674 210372 155314
rect 210436 154873 210464 155615
rect 210422 154864 210478 154873
rect 210422 154799 210478 154808
rect 210896 152318 210924 228890
rect 210988 228818 211016 236535
rect 211080 235414 211108 319398
rect 212264 316668 212316 316674
rect 212264 316610 212316 316616
rect 211988 311228 212040 311234
rect 211988 311170 212040 311176
rect 211618 297392 211674 297401
rect 211618 297327 211674 297336
rect 211068 235408 211120 235414
rect 211068 235350 211120 235356
rect 211080 234682 211108 235350
rect 211080 234654 211200 234682
rect 211068 228880 211120 228886
rect 211068 228822 211120 228828
rect 210976 228812 211028 228818
rect 210976 228754 211028 228760
rect 210884 152312 210936 152318
rect 210884 152254 210936 152260
rect 211080 149870 211108 228822
rect 211068 149864 211120 149870
rect 211068 149806 211120 149812
rect 211080 149410 211108 149806
rect 211172 149569 211200 234654
rect 211632 234054 211660 297327
rect 212000 242078 212028 311170
rect 212172 310480 212224 310486
rect 212172 310422 212224 310428
rect 212078 307456 212134 307465
rect 212078 307391 212134 307400
rect 211988 242072 212040 242078
rect 211988 242014 212040 242020
rect 211710 239184 211766 239193
rect 211710 239119 211766 239128
rect 211620 234048 211672 234054
rect 211620 233990 211672 233996
rect 211724 155009 211752 239119
rect 211988 239012 212040 239018
rect 211988 238954 212040 238960
rect 211804 236972 211856 236978
rect 211804 236914 211856 236920
rect 211816 159526 211844 236914
rect 211896 233912 211948 233918
rect 211896 233854 211948 233860
rect 211804 159520 211856 159526
rect 211804 159462 211856 159468
rect 211804 156324 211856 156330
rect 211804 156266 211856 156272
rect 211816 155990 211844 156266
rect 211804 155984 211856 155990
rect 211804 155926 211856 155932
rect 211710 155000 211766 155009
rect 211710 154935 211766 154944
rect 211158 149560 211214 149569
rect 211158 149495 211214 149504
rect 211080 149382 211200 149410
rect 210344 147646 210464 147674
rect 209792 6886 209912 6914
rect 209688 4140 209740 4146
rect 209688 4082 209740 4088
rect 209792 480 209820 6886
rect 210436 3126 210464 147646
rect 211172 16574 211200 149382
rect 211172 16546 211752 16574
rect 210976 4140 211028 4146
rect 210976 4082 211028 4088
rect 210424 3120 210476 3126
rect 210424 3062 210476 3068
rect 210988 480 211016 4082
rect 207358 354 207470 480
rect 207032 326 207470 354
rect 207358 -960 207470 326
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 211724 354 211752 16546
rect 211816 4010 211844 155926
rect 211908 144673 211936 233854
rect 212000 152250 212028 238954
rect 212092 238377 212120 307391
rect 212078 238368 212134 238377
rect 212078 238303 212134 238312
rect 212184 236473 212212 310422
rect 212276 241058 212304 316610
rect 212354 315344 212410 315353
rect 212354 315279 212410 315288
rect 212264 241052 212316 241058
rect 212264 240994 212316 241000
rect 212276 239018 212304 240994
rect 212264 239012 212316 239018
rect 212264 238954 212316 238960
rect 212368 238134 212396 315279
rect 212448 313336 212500 313342
rect 212448 313278 212500 313284
rect 212356 238128 212408 238134
rect 212356 238070 212408 238076
rect 212368 237862 212396 238070
rect 212356 237856 212408 237862
rect 212356 237798 212408 237804
rect 212170 236464 212226 236473
rect 212170 236399 212226 236408
rect 212184 154057 212212 236399
rect 212460 233918 212488 313278
rect 212908 295928 212960 295934
rect 212908 295870 212960 295876
rect 212448 233912 212500 233918
rect 212448 233854 212500 233860
rect 212448 229968 212500 229974
rect 212448 229910 212500 229916
rect 212264 229900 212316 229906
rect 212264 229842 212316 229848
rect 212276 155990 212304 229842
rect 212264 155984 212316 155990
rect 212264 155926 212316 155932
rect 212460 155038 212488 229910
rect 212920 217462 212948 295870
rect 213000 295792 213052 295798
rect 213000 295734 213052 295740
rect 212908 217456 212960 217462
rect 212908 217398 212960 217404
rect 213012 216102 213040 295734
rect 213104 239766 213132 319631
rect 213828 318096 213880 318102
rect 213828 318038 213880 318044
rect 213552 308508 213604 308514
rect 213552 308450 213604 308456
rect 213276 302320 213328 302326
rect 213276 302262 213328 302268
rect 213184 295860 213236 295866
rect 213184 295802 213236 295808
rect 213092 239760 213144 239766
rect 213092 239702 213144 239708
rect 213104 239601 213132 239702
rect 213090 239592 213146 239601
rect 213090 239527 213146 239536
rect 213092 236904 213144 236910
rect 213092 236846 213144 236852
rect 213000 216096 213052 216102
rect 213000 216038 213052 216044
rect 213104 156777 213132 236846
rect 213196 210594 213224 295802
rect 213288 253910 213316 302262
rect 213276 253904 213328 253910
rect 213276 253846 213328 253852
rect 213564 248414 213592 308450
rect 213736 294568 213788 294574
rect 213736 294510 213788 294516
rect 213380 248386 213592 248414
rect 213380 240446 213408 248386
rect 213368 240440 213420 240446
rect 213368 240382 213420 240388
rect 213458 240408 213514 240417
rect 213276 239012 213328 239018
rect 213276 238954 213328 238960
rect 213184 210588 213236 210594
rect 213184 210530 213236 210536
rect 213090 156768 213146 156777
rect 213090 156703 213146 156712
rect 212448 155032 212500 155038
rect 212448 154974 212500 154980
rect 212460 154630 212488 154974
rect 212448 154624 212500 154630
rect 212448 154566 212500 154572
rect 213184 154624 213236 154630
rect 213184 154566 213236 154572
rect 212170 154048 212226 154057
rect 212170 153983 212226 153992
rect 211988 152244 212040 152250
rect 211988 152186 212040 152192
rect 212538 151056 212594 151065
rect 212538 150991 212594 151000
rect 211894 144664 211950 144673
rect 211894 144599 211950 144608
rect 212552 16574 212580 150991
rect 212552 16546 213132 16574
rect 211804 4004 211856 4010
rect 211804 3946 211856 3952
rect 213104 3482 213132 16546
rect 213196 3942 213224 154566
rect 213288 145450 213316 238954
rect 213380 147393 213408 240382
rect 213458 240343 213514 240352
rect 213472 152425 213500 240343
rect 213644 239352 213696 239358
rect 213644 239294 213696 239300
rect 213552 234796 213604 234802
rect 213552 234738 213604 234744
rect 213458 152416 213514 152425
rect 213458 152351 213514 152360
rect 213564 151706 213592 234738
rect 213656 156670 213684 239294
rect 213748 211954 213776 294510
rect 213840 236706 213868 318038
rect 214840 315512 214892 315518
rect 214840 315454 214892 315460
rect 214748 311296 214800 311302
rect 214748 311238 214800 311244
rect 214472 305720 214524 305726
rect 214472 305662 214524 305668
rect 214484 237182 214512 305662
rect 214656 305652 214708 305658
rect 214656 305594 214708 305600
rect 214564 239828 214616 239834
rect 214564 239770 214616 239776
rect 214472 237176 214524 237182
rect 214472 237118 214524 237124
rect 213828 236700 213880 236706
rect 213828 236642 213880 236648
rect 213840 236570 213868 236642
rect 213828 236564 213880 236570
rect 213828 236506 213880 236512
rect 214484 236230 214512 237118
rect 214472 236224 214524 236230
rect 214472 236166 214524 236172
rect 213736 211948 213788 211954
rect 213736 211890 213788 211896
rect 213644 156664 213696 156670
rect 213644 156606 213696 156612
rect 213918 156632 213974 156641
rect 213918 156567 213974 156576
rect 213552 151700 213604 151706
rect 213552 151642 213604 151648
rect 213366 147384 213422 147393
rect 213366 147319 213422 147328
rect 213276 145444 213328 145450
rect 213276 145386 213328 145392
rect 213932 16574 213960 156567
rect 214576 153950 214604 239770
rect 214668 237153 214696 305594
rect 214760 239222 214788 311238
rect 214852 240378 214880 315454
rect 214932 315444 214984 315450
rect 214932 315386 214984 315392
rect 214944 240922 214972 315386
rect 214932 240916 214984 240922
rect 214932 240858 214984 240864
rect 214840 240372 214892 240378
rect 214840 240314 214892 240320
rect 214748 239216 214800 239222
rect 214748 239158 214800 239164
rect 214654 237144 214710 237153
rect 214654 237079 214710 237088
rect 214564 153944 214616 153950
rect 214564 153886 214616 153892
rect 214380 151768 214432 151774
rect 214380 151710 214432 151716
rect 214392 150482 214420 151710
rect 214380 150476 214432 150482
rect 214380 150418 214432 150424
rect 213932 16546 214512 16574
rect 213184 3936 213236 3942
rect 213184 3878 213236 3884
rect 213104 3454 213408 3482
rect 213380 480 213408 3454
rect 214484 480 214512 16546
rect 214576 3874 214604 153886
rect 214668 150346 214696 237079
rect 214852 235385 214880 240314
rect 214838 235376 214894 235385
rect 214838 235311 214894 235320
rect 214748 234592 214800 234598
rect 214748 234534 214800 234540
rect 214760 234122 214788 234534
rect 214748 234116 214800 234122
rect 214748 234058 214800 234064
rect 214748 230444 214800 230450
rect 214748 230386 214800 230392
rect 214656 150340 214708 150346
rect 214656 150282 214708 150288
rect 214760 147257 214788 230386
rect 214944 228750 214972 240858
rect 215036 239562 215064 319903
rect 216312 319592 216364 319598
rect 216312 319534 216364 319540
rect 215116 316804 215168 316810
rect 215116 316746 215168 316752
rect 215024 239556 215076 239562
rect 215024 239498 215076 239504
rect 215128 236881 215156 316746
rect 216220 314016 216272 314022
rect 216220 313958 216272 313964
rect 215208 313404 215260 313410
rect 215208 313346 215260 313352
rect 215114 236872 215170 236881
rect 215114 236807 215170 236816
rect 215024 236224 215076 236230
rect 215024 236166 215076 236172
rect 214932 228744 214984 228750
rect 214932 228686 214984 228692
rect 215036 153785 215064 236166
rect 215022 153776 215078 153785
rect 215022 153711 215078 153720
rect 215128 152726 215156 236807
rect 215220 234598 215248 313346
rect 216126 307320 216182 307329
rect 216126 307255 216182 307264
rect 216036 299668 216088 299674
rect 216036 299610 216088 299616
rect 215944 291848 215996 291854
rect 215944 291790 215996 291796
rect 215956 246362 215984 291790
rect 215944 246356 215996 246362
rect 215944 246298 215996 246304
rect 215760 241460 215812 241466
rect 215760 241402 215812 241408
rect 215772 239154 215800 241402
rect 216048 239426 216076 299610
rect 216036 239420 216088 239426
rect 216036 239362 216088 239368
rect 215760 239148 215812 239154
rect 215760 239090 215812 239096
rect 215208 234592 215260 234598
rect 215208 234534 215260 234540
rect 215208 230036 215260 230042
rect 215208 229978 215260 229984
rect 215116 152720 215168 152726
rect 215116 152662 215168 152668
rect 215220 151774 215248 229978
rect 215772 155582 215800 239090
rect 215944 238876 215996 238882
rect 215944 238818 215996 238824
rect 215852 237312 215904 237318
rect 215852 237254 215904 237260
rect 215760 155576 215812 155582
rect 215760 155518 215812 155524
rect 215208 151768 215260 151774
rect 215208 151710 215260 151716
rect 215864 148617 215892 237254
rect 215956 155786 215984 238818
rect 216140 237017 216168 307255
rect 216232 241346 216260 313958
rect 216324 241466 216352 319534
rect 217692 316056 217744 316062
rect 217692 315998 217744 316004
rect 216404 315308 216456 315314
rect 216404 315250 216456 315256
rect 216312 241460 216364 241466
rect 216312 241402 216364 241408
rect 216232 241318 216352 241346
rect 216324 239494 216352 241318
rect 216312 239488 216364 239494
rect 216312 239430 216364 239436
rect 216126 237008 216182 237017
rect 216126 236943 216182 236952
rect 216036 235476 216088 235482
rect 216036 235418 216088 235424
rect 215944 155780 215996 155786
rect 215944 155722 215996 155728
rect 215944 150476 215996 150482
rect 215944 150418 215996 150424
rect 215850 148608 215906 148617
rect 215850 148543 215906 148552
rect 215864 147801 215892 148543
rect 215298 147792 215354 147801
rect 215298 147727 215354 147736
rect 215850 147792 215906 147801
rect 215850 147727 215906 147736
rect 214746 147248 214802 147257
rect 214746 147183 214802 147192
rect 214564 3868 214616 3874
rect 214564 3810 214616 3816
rect 212142 354 212254 480
rect 211724 326 212254 354
rect 212142 -960 212254 326
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215312 354 215340 147727
rect 215956 3670 215984 150418
rect 216048 144362 216076 235418
rect 216140 230450 216168 236943
rect 216312 235068 216364 235074
rect 216312 235010 216364 235016
rect 216220 235000 216272 235006
rect 216220 234942 216272 234948
rect 216128 230444 216180 230450
rect 216128 230386 216180 230392
rect 216232 149666 216260 234942
rect 216324 155242 216352 235010
rect 216416 233918 216444 315250
rect 217600 307148 217652 307154
rect 217600 307090 217652 307096
rect 217416 305856 217468 305862
rect 217416 305798 217468 305804
rect 216496 294024 216548 294030
rect 216496 293966 216548 293972
rect 216404 233912 216456 233918
rect 216404 233854 216456 233860
rect 216416 232762 216444 233854
rect 216404 232756 216456 232762
rect 216404 232698 216456 232704
rect 216508 213382 216536 293966
rect 216588 292732 216640 292738
rect 216588 292674 216640 292680
rect 216496 213376 216548 213382
rect 216496 213318 216548 213324
rect 216600 212158 216628 292674
rect 217232 291712 217284 291718
rect 217232 291654 217284 291660
rect 217244 247722 217272 291654
rect 217324 291304 217376 291310
rect 217324 291246 217376 291252
rect 217232 247716 217284 247722
rect 217232 247658 217284 247664
rect 217336 244934 217364 291246
rect 217324 244928 217376 244934
rect 217324 244870 217376 244876
rect 217428 241233 217456 305798
rect 217508 305788 217560 305794
rect 217508 305730 217560 305736
rect 217414 241224 217470 241233
rect 217414 241159 217470 241168
rect 217428 239426 217456 241159
rect 217416 239420 217468 239426
rect 217416 239362 217468 239368
rect 217520 238785 217548 305730
rect 217612 241262 217640 307090
rect 217600 241256 217652 241262
rect 217600 241198 217652 241204
rect 217612 239834 217640 241198
rect 217704 241194 217732 315998
rect 217782 315480 217838 315489
rect 217782 315415 217838 315424
rect 217692 241188 217744 241194
rect 217692 241130 217744 241136
rect 217600 239828 217652 239834
rect 217600 239770 217652 239776
rect 217600 239420 217652 239426
rect 217600 239362 217652 239368
rect 217506 238776 217562 238785
rect 217506 238711 217562 238720
rect 217414 237280 217470 237289
rect 217414 237215 217470 237224
rect 217428 236881 217456 237215
rect 217414 236872 217470 236881
rect 217414 236807 217470 236816
rect 217324 235952 217376 235958
rect 217324 235894 217376 235900
rect 217232 234932 217284 234938
rect 217232 234874 217284 234880
rect 217244 234734 217272 234874
rect 217232 234728 217284 234734
rect 217232 234670 217284 234676
rect 216588 212152 216640 212158
rect 216588 212094 216640 212100
rect 216312 155236 216364 155242
rect 216312 155178 216364 155184
rect 217336 154086 217364 235894
rect 217324 154080 217376 154086
rect 217324 154022 217376 154028
rect 217324 153196 217376 153202
rect 217324 153138 217376 153144
rect 217336 152522 217364 153138
rect 217324 152516 217376 152522
rect 217324 152458 217376 152464
rect 216220 149660 216272 149666
rect 216220 149602 216272 149608
rect 216036 144356 216088 144362
rect 216036 144298 216088 144304
rect 216678 140040 216734 140049
rect 216678 139975 216734 139984
rect 216692 16574 216720 139975
rect 216692 16546 216904 16574
rect 215944 3664 215996 3670
rect 215944 3606 215996 3612
rect 216876 480 216904 16546
rect 217336 3806 217364 152458
rect 217428 141409 217456 236807
rect 217520 149734 217548 238711
rect 217612 152833 217640 239362
rect 217796 237289 217824 315415
rect 217888 239358 217916 320486
rect 217876 239352 217928 239358
rect 217876 239294 217928 239300
rect 217980 237998 218008 320991
rect 218612 291984 218664 291990
rect 218612 291926 218664 291932
rect 218520 291916 218572 291922
rect 218520 291858 218572 291864
rect 218058 291816 218114 291825
rect 218058 291751 218114 291760
rect 218072 289338 218100 291751
rect 218060 289332 218112 289338
rect 218060 289274 218112 289280
rect 217968 237992 218020 237998
rect 217968 237934 218020 237940
rect 217782 237280 217838 237289
rect 217782 237215 217838 237224
rect 217692 236020 217744 236026
rect 217692 235962 217744 235968
rect 217704 157049 217732 235962
rect 217784 228744 217836 228750
rect 217784 228686 217836 228692
rect 217690 157040 217746 157049
rect 217690 156975 217746 156984
rect 217796 153202 217824 228686
rect 218532 201385 218560 291858
rect 218624 271182 218652 291926
rect 218612 271176 218664 271182
rect 218612 271118 218664 271124
rect 218612 240848 218664 240854
rect 218612 240790 218664 240796
rect 218624 240310 218652 240790
rect 218612 240304 218664 240310
rect 218612 240246 218664 240252
rect 218716 240174 218744 321710
rect 219072 316872 219124 316878
rect 219072 316814 219124 316820
rect 218978 307184 219034 307193
rect 218978 307119 219034 307128
rect 218796 298308 218848 298314
rect 218796 298250 218848 298256
rect 218704 240168 218756 240174
rect 218704 240110 218756 240116
rect 218716 239970 218744 240110
rect 218704 239964 218756 239970
rect 218704 239906 218756 239912
rect 218612 239488 218664 239494
rect 218612 239430 218664 239436
rect 218704 239488 218756 239494
rect 218704 239430 218756 239436
rect 218624 237289 218652 239430
rect 218610 237280 218666 237289
rect 218610 237215 218666 237224
rect 218716 233714 218744 239430
rect 218704 233708 218756 233714
rect 218704 233650 218756 233656
rect 218716 232393 218744 233650
rect 218702 232384 218758 232393
rect 218702 232319 218758 232328
rect 218704 229764 218756 229770
rect 218704 229706 218756 229712
rect 218058 201376 218114 201385
rect 218058 201311 218114 201320
rect 218518 201376 218574 201385
rect 218518 201311 218574 201320
rect 218072 200705 218100 201311
rect 218058 200696 218114 200705
rect 218058 200631 218114 200640
rect 217784 153196 217836 153202
rect 217784 153138 217836 153144
rect 217598 152824 217654 152833
rect 217598 152759 217654 152768
rect 217508 149728 217560 149734
rect 217508 149670 217560 149676
rect 218060 145512 218112 145518
rect 218060 145454 218112 145460
rect 218072 144906 218100 145454
rect 218060 144900 218112 144906
rect 218060 144842 218112 144848
rect 218072 142154 218100 144842
rect 218072 142126 218192 142154
rect 217414 141400 217470 141409
rect 217414 141335 217470 141344
rect 218164 16574 218192 142126
rect 218716 141574 218744 229706
rect 218808 210458 218836 298250
rect 218888 292392 218940 292398
rect 218888 292334 218940 292340
rect 218900 269822 218928 292334
rect 218888 269816 218940 269822
rect 218888 269758 218940 269764
rect 218886 240000 218942 240009
rect 218886 239935 218942 239944
rect 218900 239562 218928 239935
rect 218888 239556 218940 239562
rect 218888 239498 218940 239504
rect 218992 239290 219020 307119
rect 219084 247034 219112 316814
rect 219164 312588 219216 312594
rect 219164 312530 219216 312536
rect 219176 248414 219204 312530
rect 219268 292602 219296 374614
rect 219348 374060 219400 374066
rect 219348 374002 219400 374008
rect 219256 292596 219308 292602
rect 219256 292538 219308 292544
rect 219268 286346 219296 292538
rect 219360 291825 219388 374002
rect 220096 373930 220124 699654
rect 234632 461650 234660 703582
rect 235000 703474 235028 703582
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 250444 700324 250496 700330
rect 250444 700266 250496 700272
rect 234620 461644 234672 461650
rect 234620 461586 234672 461592
rect 220176 403640 220228 403646
rect 220176 403582 220228 403588
rect 220188 403034 220216 403582
rect 220176 403028 220228 403034
rect 220176 402970 220228 402976
rect 220084 373924 220136 373930
rect 220084 373866 220136 373872
rect 220188 291990 220216 402970
rect 244924 379840 244976 379846
rect 244924 379782 244976 379788
rect 242164 376916 242216 376922
rect 242164 376858 242216 376864
rect 232504 375624 232556 375630
rect 232504 375566 232556 375572
rect 220728 373312 220780 373318
rect 220728 373254 220780 373260
rect 220636 371884 220688 371890
rect 220636 371826 220688 371832
rect 220544 320272 220596 320278
rect 220544 320214 220596 320220
rect 220452 313948 220504 313954
rect 220452 313890 220504 313896
rect 220268 302932 220320 302938
rect 220268 302874 220320 302880
rect 220176 291984 220228 291990
rect 220176 291926 220228 291932
rect 219346 291816 219402 291825
rect 219346 291751 219402 291760
rect 219900 291780 219952 291786
rect 219900 291722 219952 291728
rect 219808 291372 219860 291378
rect 219808 291314 219860 291320
rect 219716 289808 219768 289814
rect 219716 289750 219768 289756
rect 219256 286340 219308 286346
rect 219256 286282 219308 286288
rect 219176 248386 219388 248414
rect 219084 247006 219204 247034
rect 219176 240514 219204 247006
rect 219164 240508 219216 240514
rect 219164 240450 219216 240456
rect 219072 239556 219124 239562
rect 219072 239498 219124 239504
rect 218980 239284 219032 239290
rect 218980 239226 219032 239232
rect 218992 238746 219020 239226
rect 218980 238740 219032 238746
rect 218980 238682 219032 238688
rect 218888 237992 218940 237998
rect 218888 237934 218940 237940
rect 218900 236774 218928 237934
rect 218888 236768 218940 236774
rect 218888 236710 218940 236716
rect 218980 236768 219032 236774
rect 218980 236710 219032 236716
rect 218888 235340 218940 235346
rect 218888 235282 218940 235288
rect 218796 210452 218848 210458
rect 218796 210394 218848 210400
rect 218900 149598 218928 235282
rect 218992 153066 219020 236710
rect 219084 155650 219112 239498
rect 219176 235958 219204 240450
rect 219360 239494 219388 248386
rect 219348 239488 219400 239494
rect 219348 239430 219400 239436
rect 219440 238740 219492 238746
rect 219440 238682 219492 238688
rect 219164 235952 219216 235958
rect 219164 235894 219216 235900
rect 219256 235272 219308 235278
rect 219256 235214 219308 235220
rect 219268 159458 219296 235214
rect 219256 159452 219308 159458
rect 219256 159394 219308 159400
rect 219072 155644 219124 155650
rect 219072 155586 219124 155592
rect 218980 153060 219032 153066
rect 218980 153002 219032 153008
rect 219452 150006 219480 238682
rect 219728 238338 219756 289750
rect 219820 273970 219848 291314
rect 219808 273964 219860 273970
rect 219808 273906 219860 273912
rect 219912 272542 219940 291722
rect 219990 291680 220046 291689
rect 219990 291615 220046 291624
rect 219900 272536 219952 272542
rect 219900 272478 219952 272484
rect 220004 242282 220032 291615
rect 220084 291508 220136 291514
rect 220084 291450 220136 291456
rect 219992 242276 220044 242282
rect 219992 242218 220044 242224
rect 220096 239698 220124 291450
rect 219992 239692 220044 239698
rect 219992 239634 220044 239640
rect 220084 239692 220136 239698
rect 220084 239634 220136 239640
rect 220004 239601 220032 239634
rect 219990 239592 220046 239601
rect 219990 239527 220046 239536
rect 219898 239048 219954 239057
rect 219898 238983 219954 238992
rect 219716 238332 219768 238338
rect 219716 238274 219768 238280
rect 219912 238270 219940 238983
rect 219900 238264 219952 238270
rect 219900 238206 219952 238212
rect 220280 237318 220308 302874
rect 220360 290216 220412 290222
rect 220360 290158 220412 290164
rect 220268 237312 220320 237318
rect 220268 237254 220320 237260
rect 220176 236700 220228 236706
rect 220176 236642 220228 236648
rect 220082 228304 220138 228313
rect 220082 228239 220138 228248
rect 219440 150000 219492 150006
rect 219440 149942 219492 149948
rect 218888 149592 218940 149598
rect 218888 149534 218940 149540
rect 218704 141568 218756 141574
rect 218704 141510 218756 141516
rect 220096 141273 220124 228239
rect 220188 152561 220216 236642
rect 220372 212498 220400 290158
rect 220464 236201 220492 313890
rect 220556 240650 220584 320214
rect 220648 290766 220676 371826
rect 220636 290760 220688 290766
rect 220636 290702 220688 290708
rect 220740 290698 220768 373254
rect 222106 372872 222162 372881
rect 222106 372807 222162 372816
rect 222014 312488 222070 312497
rect 222014 312423 222070 312432
rect 221924 308440 221976 308446
rect 221924 308382 221976 308388
rect 221740 299464 221792 299470
rect 221740 299406 221792 299412
rect 221464 292120 221516 292126
rect 221464 292062 221516 292068
rect 220820 292052 220872 292058
rect 220820 291994 220872 292000
rect 220728 290692 220780 290698
rect 220728 290634 220780 290640
rect 220740 290465 220768 290634
rect 220726 290456 220782 290465
rect 220726 290391 220782 290400
rect 220832 280838 220860 291994
rect 221280 291644 221332 291650
rect 221280 291586 221332 291592
rect 220912 291440 220964 291446
rect 220912 291382 220964 291388
rect 220924 284986 220952 291382
rect 221292 287054 221320 291586
rect 221372 291576 221424 291582
rect 221372 291518 221424 291524
rect 221016 287026 221320 287054
rect 220912 284980 220964 284986
rect 220912 284922 220964 284928
rect 221016 283642 221044 287026
rect 220924 283626 221044 283642
rect 220912 283620 221044 283626
rect 220964 283614 221044 283620
rect 220912 283562 220964 283568
rect 221384 282282 221412 291518
rect 220924 282254 221412 282282
rect 220924 282198 220952 282254
rect 220912 282192 220964 282198
rect 220912 282134 220964 282140
rect 220820 280832 220872 280838
rect 220820 280774 220872 280780
rect 221476 279562 221504 292062
rect 221752 291854 221780 299406
rect 221740 291848 221792 291854
rect 221740 291790 221792 291796
rect 221556 290352 221608 290358
rect 221556 290294 221608 290300
rect 220924 279534 221504 279562
rect 220924 279478 220952 279534
rect 220912 279472 220964 279478
rect 220912 279414 220964 279420
rect 221096 242072 221148 242078
rect 221096 242014 221148 242020
rect 221188 242072 221240 242078
rect 221188 242014 221240 242020
rect 220544 240644 220596 240650
rect 220544 240586 220596 240592
rect 220556 238796 220584 240586
rect 221108 240378 221136 242014
rect 221200 241913 221228 242014
rect 221186 241904 221242 241913
rect 221186 241839 221242 241848
rect 221096 240372 221148 240378
rect 221096 240314 221148 240320
rect 221096 239828 221148 239834
rect 221096 239770 221148 239776
rect 220636 239556 220688 239562
rect 220636 239498 220688 239504
rect 220728 239556 220780 239562
rect 220728 239498 220780 239504
rect 220648 238921 220676 239498
rect 220634 238912 220690 238921
rect 220634 238847 220690 238856
rect 220556 238768 220676 238796
rect 220544 238332 220596 238338
rect 220544 238274 220596 238280
rect 220556 238134 220584 238274
rect 220544 238128 220596 238134
rect 220544 238070 220596 238076
rect 220450 236192 220506 236201
rect 220450 236127 220506 236136
rect 220464 232801 220492 236127
rect 220450 232792 220506 232801
rect 220450 232727 220506 232736
rect 220360 212492 220412 212498
rect 220360 212434 220412 212440
rect 220556 156534 220584 238070
rect 220544 156528 220596 156534
rect 220544 156470 220596 156476
rect 220648 155514 220676 238768
rect 220636 155508 220688 155514
rect 220636 155450 220688 155456
rect 220740 153746 220768 239498
rect 220912 239488 220964 239494
rect 220912 239430 220964 239436
rect 220924 239329 220952 239430
rect 220910 239320 220966 239329
rect 220910 239255 220966 239264
rect 221108 239222 221136 239770
rect 221096 239216 221148 239222
rect 221096 239158 221148 239164
rect 221200 239086 221228 241839
rect 221462 240952 221518 240961
rect 221462 240887 221518 240896
rect 221372 240236 221424 240242
rect 221372 240178 221424 240184
rect 221280 240100 221332 240106
rect 221280 240042 221332 240048
rect 221188 239080 221240 239086
rect 221188 239022 221240 239028
rect 221292 238814 221320 240042
rect 221280 238808 221332 238814
rect 221280 238750 221332 238756
rect 221384 238542 221412 240178
rect 221476 240038 221504 240887
rect 221464 240032 221516 240038
rect 221464 239974 221516 239980
rect 221462 239456 221518 239465
rect 221462 239391 221518 239400
rect 221476 238814 221504 239391
rect 221464 238808 221516 238814
rect 221464 238750 221516 238756
rect 221372 238536 221424 238542
rect 221372 238478 221424 238484
rect 221004 235612 221056 235618
rect 221004 235554 221056 235560
rect 221016 235414 221044 235554
rect 221004 235408 221056 235414
rect 221004 235350 221056 235356
rect 221462 233744 221518 233753
rect 221462 233679 221518 233688
rect 220728 153740 220780 153746
rect 220728 153682 220780 153688
rect 220174 152552 220230 152561
rect 220174 152487 220230 152496
rect 220728 150000 220780 150006
rect 220728 149942 220780 149948
rect 220740 149734 220768 149942
rect 220728 149728 220780 149734
rect 220728 149670 220780 149676
rect 221476 144498 221504 233679
rect 221568 212226 221596 290294
rect 221648 290284 221700 290290
rect 221648 290226 221700 290232
rect 221660 212294 221688 290226
rect 221740 289944 221792 289950
rect 221740 289886 221792 289892
rect 221648 212288 221700 212294
rect 221648 212230 221700 212236
rect 221556 212220 221608 212226
rect 221556 212162 221608 212168
rect 221752 212022 221780 289886
rect 221830 246392 221886 246401
rect 221830 246327 221886 246336
rect 221844 235958 221872 246327
rect 221936 244338 221964 308382
rect 222028 246401 222056 312423
rect 222120 291922 222148 372807
rect 229744 371952 229796 371958
rect 229744 371894 229796 371900
rect 224866 370152 224922 370161
rect 224866 370087 224922 370096
rect 224222 370016 224278 370025
rect 224222 369951 224278 369960
rect 222200 310004 222252 310010
rect 222200 309946 222252 309952
rect 222108 291916 222160 291922
rect 222108 291858 222160 291864
rect 222212 269114 222240 309946
rect 222476 294704 222528 294710
rect 222476 294646 222528 294652
rect 222120 269086 222240 269114
rect 222014 246392 222070 246401
rect 222014 246327 222070 246336
rect 221936 244310 222056 244338
rect 222028 244202 222056 244310
rect 221936 244174 222056 244202
rect 221832 235952 221884 235958
rect 221832 235894 221884 235900
rect 221936 232694 221964 244174
rect 222120 240394 222148 269086
rect 222488 242078 222516 294646
rect 224236 293078 224264 369951
rect 224316 319048 224368 319054
rect 224316 318990 224368 318996
rect 224224 293072 224276 293078
rect 224224 293014 224276 293020
rect 224328 290306 224356 318990
rect 224880 294642 224908 370087
rect 228362 369336 228418 369345
rect 228362 369271 228418 369280
rect 225602 369200 225658 369209
rect 225602 369135 225658 369144
rect 224868 294636 224920 294642
rect 224868 294578 224920 294584
rect 224880 293978 224908 294578
rect 225616 294438 225644 369135
rect 226984 358828 227036 358834
rect 226984 358770 227036 358776
rect 225694 321192 225750 321201
rect 225694 321127 225750 321136
rect 225604 294432 225656 294438
rect 225604 294374 225656 294380
rect 225616 294098 225644 294374
rect 225604 294092 225656 294098
rect 225604 294034 225656 294040
rect 224880 293950 225000 293978
rect 224684 293072 224736 293078
rect 224684 293014 224736 293020
rect 224408 291916 224460 291922
rect 224408 291858 224460 291864
rect 224144 290278 224356 290306
rect 224144 289898 224172 290278
rect 224222 290184 224278 290193
rect 224420 290170 224448 291858
rect 224222 290119 224278 290128
rect 224328 290142 224448 290170
rect 224236 289921 224264 290119
rect 223592 289870 224172 289898
rect 224222 289912 224278 289921
rect 223592 289814 223620 289870
rect 224328 289884 224356 290142
rect 224696 289884 224724 293014
rect 224972 289898 225000 293950
rect 225708 293350 225736 321127
rect 225786 317520 225842 317529
rect 225786 317455 225842 317464
rect 225800 295361 225828 317455
rect 226996 296714 227024 358770
rect 227076 351212 227128 351218
rect 227076 351154 227128 351160
rect 226904 296686 227024 296714
rect 227088 296714 227116 351154
rect 227166 318608 227222 318617
rect 227166 318543 227222 318552
rect 227180 301617 227208 318543
rect 228376 306374 228404 369271
rect 228456 322244 228508 322250
rect 228456 322186 228508 322192
rect 228284 306346 228404 306374
rect 227166 301608 227222 301617
rect 227166 301543 227222 301552
rect 227088 296686 227208 296714
rect 225786 295352 225842 295361
rect 225786 295287 225842 295296
rect 226904 294166 226932 296686
rect 226892 294160 226944 294166
rect 226892 294102 226944 294108
rect 225788 294092 225840 294098
rect 225788 294034 225840 294040
rect 225696 293344 225748 293350
rect 225696 293286 225748 293292
rect 225708 289898 225736 293286
rect 224972 289870 225078 289898
rect 225446 289870 225736 289898
rect 225800 289884 225828 294034
rect 226340 293956 226392 293962
rect 226340 293898 226392 293904
rect 226352 293282 226380 293898
rect 226340 293276 226392 293282
rect 226340 293218 226392 293224
rect 226154 291272 226210 291281
rect 226154 291207 226210 291216
rect 226168 289884 226196 291207
rect 226352 289898 226380 293218
rect 226352 289870 226550 289898
rect 226904 289884 226932 294102
rect 227180 291310 227208 296686
rect 228284 294846 228312 306346
rect 228468 296714 228496 322186
rect 228376 296686 228496 296714
rect 228272 294840 228324 294846
rect 228272 294782 228324 294788
rect 227718 291816 227774 291825
rect 227718 291751 227774 291760
rect 227732 291310 227760 291751
rect 227168 291304 227220 291310
rect 227168 291246 227220 291252
rect 227720 291304 227772 291310
rect 227720 291246 227772 291252
rect 227180 289898 227208 291246
rect 227812 291236 227864 291242
rect 227812 291178 227864 291184
rect 227824 290766 227852 291178
rect 227812 290760 227864 290766
rect 227812 290702 227864 290708
rect 227626 290456 227682 290465
rect 227626 290391 227682 290400
rect 227180 289870 227286 289898
rect 227640 289884 227668 290391
rect 228284 289898 228312 294782
rect 228376 291417 228404 296686
rect 229100 294772 229152 294778
rect 229100 294714 229152 294720
rect 228732 292596 228784 292602
rect 228732 292538 228784 292544
rect 228362 291408 228418 291417
rect 228362 291343 228418 291352
rect 228022 289870 228312 289898
rect 228376 289884 228404 291343
rect 228744 289884 228772 292538
rect 229112 289884 229140 294714
rect 229756 293962 229784 371894
rect 231768 370660 231820 370666
rect 231768 370602 231820 370608
rect 229836 368688 229888 368694
rect 229836 368630 229888 368636
rect 229926 368656 229982 368665
rect 229848 294778 229876 368630
rect 229926 368591 229982 368600
rect 231124 368620 231176 368626
rect 229836 294772 229888 294778
rect 229836 294714 229888 294720
rect 229940 294370 229968 368591
rect 231124 368562 231176 368568
rect 230018 323640 230074 323649
rect 230018 323575 230074 323584
rect 229928 294364 229980 294370
rect 229928 294306 229980 294312
rect 229744 293956 229796 293962
rect 229744 293898 229796 293904
rect 230032 291718 230060 323575
rect 230480 297492 230532 297498
rect 230480 297434 230532 297440
rect 230492 296070 230520 297434
rect 230480 296064 230532 296070
rect 230480 296006 230532 296012
rect 230204 294364 230256 294370
rect 230204 294306 230256 294312
rect 229468 291712 229520 291718
rect 229468 291654 229520 291660
rect 230020 291712 230072 291718
rect 230020 291654 230072 291660
rect 229480 289884 229508 291654
rect 229836 291236 229888 291242
rect 229836 291178 229888 291184
rect 229848 289884 229876 291178
rect 230216 289884 230244 294306
rect 230492 289898 230520 296006
rect 230940 295384 230992 295390
rect 230940 295326 230992 295332
rect 230952 290834 230980 295326
rect 231136 294506 231164 368562
rect 231780 296714 231808 370602
rect 232516 296714 232544 375566
rect 236644 375556 236696 375562
rect 236644 375498 236696 375504
rect 233884 373244 233936 373250
rect 233884 373186 233936 373192
rect 233148 370728 233200 370734
rect 233148 370670 233200 370676
rect 233160 298790 233188 370670
rect 233330 318472 233386 318481
rect 233330 318407 233386 318416
rect 233344 315625 233372 318407
rect 233330 315616 233386 315625
rect 233330 315551 233386 315560
rect 233148 298784 233200 298790
rect 233148 298726 233200 298732
rect 231688 296686 231808 296714
rect 232424 296686 232544 296714
rect 231688 295390 231716 296686
rect 232424 295594 232452 296686
rect 232412 295588 232464 295594
rect 232412 295530 232464 295536
rect 231676 295384 231728 295390
rect 231676 295326 231728 295332
rect 232044 294568 232096 294574
rect 232044 294510 232096 294516
rect 231124 294500 231176 294506
rect 231124 294442 231176 294448
rect 230940 290828 230992 290834
rect 230940 290770 230992 290776
rect 230492 289870 230598 289898
rect 230952 289884 230980 290770
rect 231136 289898 231164 294442
rect 231582 289912 231638 289921
rect 231136 289870 231334 289898
rect 224222 289847 224278 289856
rect 231638 289870 231702 289898
rect 232056 289884 232084 294510
rect 232424 289884 232452 295530
rect 233160 294574 233188 298726
rect 233896 295662 233924 373186
rect 235264 370388 235316 370394
rect 235264 370330 235316 370336
rect 233976 369164 234028 369170
rect 233976 369106 234028 369112
rect 233884 295656 233936 295662
rect 233884 295598 233936 295604
rect 233896 295390 233924 295598
rect 233988 295526 234016 369106
rect 234068 324964 234120 324970
rect 234068 324906 234120 324912
rect 234080 297294 234108 324906
rect 235276 306374 235304 370330
rect 235356 327752 235408 327758
rect 235356 327694 235408 327700
rect 235184 306346 235304 306374
rect 234068 297288 234120 297294
rect 234068 297230 234120 297236
rect 233976 295520 234028 295526
rect 233976 295462 234028 295468
rect 233884 295384 233936 295390
rect 233884 295326 233936 295332
rect 233148 294568 233200 294574
rect 233148 294510 233200 294516
rect 233988 293842 234016 295462
rect 233804 293814 234016 293842
rect 233148 293140 233200 293146
rect 233148 293082 233200 293088
rect 232780 292868 232832 292874
rect 232780 292810 232832 292816
rect 232792 291718 232820 292810
rect 232780 291712 232832 291718
rect 232780 291654 232832 291660
rect 232792 289884 232820 291654
rect 233160 291106 233188 293082
rect 233148 291100 233200 291106
rect 233148 291042 233200 291048
rect 233160 289884 233188 291042
rect 233804 289898 233832 293814
rect 234080 289898 234108 297230
rect 235184 296002 235212 306346
rect 235368 296954 235396 327694
rect 236656 297090 236684 375498
rect 238668 375488 238720 375494
rect 238668 375430 238720 375436
rect 238024 370048 238076 370054
rect 238024 369990 238076 369996
rect 236644 297084 236696 297090
rect 236644 297026 236696 297032
rect 235356 296948 235408 296954
rect 235356 296890 235408 296896
rect 235368 296714 235396 296890
rect 235276 296686 235396 296714
rect 236656 296714 236684 297026
rect 238036 296714 238064 369990
rect 238574 316024 238630 316033
rect 238574 315959 238630 315968
rect 238588 306513 238616 315959
rect 238574 306504 238630 306513
rect 238574 306439 238630 306448
rect 238680 306374 238708 375430
rect 238852 374128 238904 374134
rect 238852 374070 238904 374076
rect 238760 318164 238812 318170
rect 238760 318106 238812 318112
rect 238772 314129 238800 318106
rect 238758 314120 238814 314129
rect 238758 314055 238814 314064
rect 236656 296686 237052 296714
rect 235172 295996 235224 296002
rect 235172 295938 235224 295944
rect 234528 295384 234580 295390
rect 234528 295326 234580 295332
rect 234540 292482 234568 295326
rect 235184 292534 235212 295938
rect 235172 292528 235224 292534
rect 234540 292454 234660 292482
rect 235172 292470 235224 292476
rect 234252 291304 234304 291310
rect 234252 291246 234304 291252
rect 234158 290184 234214 290193
rect 234158 290119 234214 290128
rect 234172 289921 234200 290119
rect 233542 289870 233832 289898
rect 233910 289870 234108 289898
rect 234158 289912 234214 289921
rect 231582 289847 231638 289856
rect 234264 289884 234292 291246
rect 234632 289884 234660 292454
rect 235276 289898 235304 296686
rect 236828 296132 236880 296138
rect 236828 296074 236880 296080
rect 236840 295730 236868 296074
rect 236828 295724 236880 295730
rect 236828 295666 236880 295672
rect 235724 294772 235776 294778
rect 235724 294714 235776 294720
rect 235356 293276 235408 293282
rect 235356 293218 235408 293224
rect 235368 292738 235396 293218
rect 235356 292732 235408 292738
rect 235356 292674 235408 292680
rect 235014 289870 235304 289898
rect 235368 289884 235396 292674
rect 235736 289898 235764 294714
rect 236092 293344 236144 293350
rect 236092 293286 236144 293292
rect 236104 292806 236132 293286
rect 236092 292800 236144 292806
rect 236092 292742 236144 292748
rect 236460 292800 236512 292806
rect 236460 292742 236512 292748
rect 236092 292528 236144 292534
rect 236092 292470 236144 292476
rect 235552 289884 235764 289898
rect 236104 289884 236132 292470
rect 236472 289884 236500 292742
rect 236840 289884 236868 295666
rect 237024 289898 237052 296686
rect 237944 296686 238064 296714
rect 238588 306346 238708 306374
rect 237472 294636 237524 294642
rect 237472 294578 237524 294584
rect 237380 293412 237432 293418
rect 237380 293354 237432 293360
rect 237392 292942 237420 293354
rect 237484 293214 237512 294578
rect 237944 294234 237972 296686
rect 237932 294228 237984 294234
rect 237932 294170 237984 294176
rect 237472 293208 237524 293214
rect 237472 293150 237524 293156
rect 237380 292936 237432 292942
rect 237380 292878 237432 292884
rect 237392 292618 237420 292878
rect 237392 292590 237604 292618
rect 237472 292528 237524 292534
rect 237472 292470 237524 292476
rect 237380 292120 237432 292126
rect 237380 292062 237432 292068
rect 237392 291922 237420 292062
rect 237484 292058 237512 292470
rect 237472 292052 237524 292058
rect 237472 291994 237524 292000
rect 237380 291916 237432 291922
rect 237380 291858 237432 291864
rect 235552 289870 235750 289884
rect 237024 289870 237222 289898
rect 237576 289884 237604 292590
rect 237944 289884 237972 294170
rect 238484 293208 238536 293214
rect 238484 293150 238536 293156
rect 238300 291916 238352 291922
rect 238300 291858 238352 291864
rect 238312 289884 238340 291858
rect 238496 289898 238524 293150
rect 238588 292534 238616 306346
rect 238666 306232 238722 306241
rect 238666 306167 238722 306176
rect 238680 296857 238708 306167
rect 238666 296848 238722 296857
rect 238666 296783 238722 296792
rect 238666 296712 238722 296721
rect 238666 296647 238722 296656
rect 238576 292528 238628 292534
rect 238576 292470 238628 292476
rect 238680 290193 238708 296647
rect 238666 290184 238722 290193
rect 238666 290119 238722 290128
rect 238864 289898 238892 374070
rect 240140 368552 240192 368558
rect 240140 368494 240192 368500
rect 240152 306374 240180 368494
rect 240152 306346 241100 306374
rect 240140 296064 240192 296070
rect 240140 296006 240192 296012
rect 239772 293004 239824 293010
rect 239772 292946 239824 292952
rect 239404 292528 239456 292534
rect 239404 292470 239456 292476
rect 238496 289870 238694 289898
rect 238864 289882 239062 289898
rect 239416 289884 239444 292470
rect 239784 291174 239812 292946
rect 239772 291168 239824 291174
rect 239772 291110 239824 291116
rect 239784 289884 239812 291110
rect 240152 289884 240180 296006
rect 240874 292632 240930 292641
rect 240874 292567 240930 292576
rect 240888 292466 240916 292567
rect 240876 292460 240928 292466
rect 240876 292402 240928 292408
rect 240508 292256 240560 292262
rect 240508 292198 240560 292204
rect 240416 289944 240468 289950
rect 240520 289898 240548 292198
rect 240468 289892 240548 289898
rect 240416 289886 240548 289892
rect 240428 289884 240548 289886
rect 240888 289884 240916 292402
rect 241072 289898 241100 306346
rect 242176 296714 242204 376858
rect 242254 371376 242310 371385
rect 242254 371311 242310 371320
rect 242268 297498 242296 371311
rect 243542 360904 243598 360913
rect 243542 360839 243598 360848
rect 242532 318300 242584 318306
rect 242532 318242 242584 318248
rect 242544 316985 242572 318242
rect 242530 316976 242586 316985
rect 242530 316911 242586 316920
rect 243556 306374 243584 360839
rect 243556 306346 243676 306374
rect 242256 297492 242308 297498
rect 242256 297434 242308 297440
rect 241900 296686 242204 296714
rect 241900 291650 241928 296686
rect 243084 295860 243136 295866
rect 243084 295802 243136 295808
rect 242808 294840 242860 294846
rect 242808 294782 242860 294788
rect 242716 294296 242768 294302
rect 242716 294238 242768 294244
rect 241980 294024 242032 294030
rect 241980 293966 242032 293972
rect 241888 291644 241940 291650
rect 241888 291586 241940 291592
rect 241900 289898 241928 291586
rect 238852 289876 239062 289882
rect 234158 289847 234214 289856
rect 223580 289808 223632 289814
rect 223580 289750 223632 289756
rect 235552 289406 235580 289870
rect 238904 289870 239062 289876
rect 240428 289870 240534 289884
rect 241072 289870 241270 289898
rect 241638 289870 241928 289898
rect 241992 289884 242020 293966
rect 242256 292528 242308 292534
rect 242728 292505 242756 294238
rect 242820 294030 242848 294782
rect 242808 294024 242860 294030
rect 242808 293966 242860 293972
rect 242256 292470 242308 292476
rect 242714 292496 242770 292505
rect 238852 289818 238904 289824
rect 238864 289787 238892 289818
rect 241072 289785 241100 289870
rect 241058 289776 241114 289785
rect 241058 289711 241114 289720
rect 242268 289490 242296 292470
rect 242714 292431 242770 292440
rect 242728 289884 242756 292431
rect 243096 289884 243124 295802
rect 243648 291582 243676 306346
rect 244556 298104 244608 298110
rect 244556 298046 244608 298052
rect 244568 296818 244596 298046
rect 244556 296812 244608 296818
rect 244556 296754 244608 296760
rect 244188 292052 244240 292058
rect 244188 291994 244240 292000
rect 243636 291576 243688 291582
rect 243636 291518 243688 291524
rect 243452 290692 243504 290698
rect 243452 290634 243504 290640
rect 243464 290426 243492 290634
rect 243452 290420 243504 290426
rect 243452 290362 243504 290368
rect 243464 289884 243492 290362
rect 243648 289898 243676 291518
rect 244200 289898 244228 291994
rect 244280 291304 244332 291310
rect 244280 291246 244332 291252
rect 244292 290193 244320 291246
rect 244278 290184 244334 290193
rect 244278 290119 244334 290128
rect 243648 289870 243846 289898
rect 244016 289884 244228 289898
rect 244568 289884 244596 296754
rect 244936 291514 244964 379782
rect 249064 379772 249116 379778
rect 249064 379714 249116 379720
rect 245016 376780 245068 376786
rect 245016 376722 245068 376728
rect 245028 297226 245056 376722
rect 245108 374196 245160 374202
rect 245108 374138 245160 374144
rect 245016 297220 245068 297226
rect 245016 297162 245068 297168
rect 244924 291508 244976 291514
rect 244924 291450 244976 291456
rect 244936 289884 244964 291450
rect 245028 291242 245056 297162
rect 245120 296138 245148 374138
rect 245752 370592 245804 370598
rect 245752 370534 245804 370540
rect 245200 370184 245252 370190
rect 245200 370126 245252 370132
rect 245212 298110 245240 370126
rect 245660 367804 245712 367810
rect 245660 367746 245712 367752
rect 245672 367062 245700 367746
rect 245660 367056 245712 367062
rect 245660 366998 245712 367004
rect 245764 354674 245792 370534
rect 248418 368928 248474 368937
rect 248418 368863 248474 368872
rect 246304 367056 246356 367062
rect 246304 366998 246356 367004
rect 245672 354646 245792 354674
rect 245672 306374 245700 354646
rect 245672 306346 245792 306374
rect 245200 298104 245252 298110
rect 245200 298046 245252 298052
rect 245108 296132 245160 296138
rect 245108 296074 245160 296080
rect 245764 292574 245792 306346
rect 245672 292546 245792 292574
rect 245292 292188 245344 292194
rect 245292 292130 245344 292136
rect 245016 291236 245068 291242
rect 245016 291178 245068 291184
rect 244016 289870 244214 289884
rect 242268 289474 242664 289490
rect 242268 289468 242676 289474
rect 242268 289462 242624 289468
rect 242624 289410 242676 289416
rect 244016 289406 244044 289870
rect 244832 289808 244884 289814
rect 244830 289776 244832 289785
rect 244884 289776 244886 289785
rect 244830 289711 244886 289720
rect 245304 289626 245332 292130
rect 245672 289626 245700 292546
rect 246316 291310 246344 366998
rect 247040 365084 247092 365090
rect 247040 365026 247092 365032
rect 246394 353968 246450 353977
rect 246394 353903 246450 353912
rect 246408 291446 246436 353903
rect 246672 292324 246724 292330
rect 246672 292266 246724 292272
rect 246396 291440 246448 291446
rect 246396 291382 246448 291388
rect 246304 291304 246356 291310
rect 246304 291246 246356 291252
rect 246408 290170 246436 291382
rect 246316 290142 246436 290170
rect 246316 289898 246344 290142
rect 246684 289898 246712 292266
rect 246764 291304 246816 291310
rect 246764 291246 246816 291252
rect 246948 291304 247000 291310
rect 246948 291246 247000 291252
rect 246054 289870 246344 289898
rect 246422 289884 246712 289898
rect 246776 289884 246804 291246
rect 246960 290737 246988 291246
rect 246946 290728 247002 290737
rect 246946 290663 247002 290672
rect 246408 289870 246712 289884
rect 246212 289808 246264 289814
rect 246408 289762 246436 289870
rect 246264 289756 246436 289762
rect 246212 289750 246436 289756
rect 246224 289748 246436 289750
rect 246224 289734 246422 289748
rect 245304 289612 245516 289626
rect 245318 289598 245516 289612
rect 245488 289513 245516 289598
rect 245580 289612 245700 289626
rect 245580 289598 245686 289612
rect 245474 289504 245530 289513
rect 245474 289439 245530 289448
rect 245580 289406 245608 289598
rect 247052 289513 247080 365026
rect 247684 365016 247736 365022
rect 247684 364958 247736 364964
rect 247696 291689 247724 364958
rect 247774 358048 247830 358057
rect 247774 357983 247830 357992
rect 247682 291680 247738 291689
rect 247682 291615 247738 291624
rect 247408 291372 247460 291378
rect 247408 291314 247460 291320
rect 247420 291122 247448 291314
rect 247696 291281 247724 291615
rect 247682 291272 247738 291281
rect 247682 291207 247738 291216
rect 247788 291122 247816 357983
rect 248432 306374 248460 368863
rect 248432 306346 248828 306374
rect 248604 295792 248656 295798
rect 248604 295734 248656 295740
rect 248234 291272 248290 291281
rect 247868 291236 247920 291242
rect 248234 291207 248290 291216
rect 247868 291178 247920 291184
rect 247420 291094 247816 291122
rect 247420 289898 247448 291094
rect 247158 289870 247448 289898
rect 247880 289884 247908 291178
rect 248248 289884 248276 291207
rect 248616 289884 248644 295734
rect 248800 289626 248828 306346
rect 249076 291786 249104 379714
rect 250456 368393 250484 700266
rect 267660 697610 267688 703520
rect 283852 702434 283880 703520
rect 282932 702406 283880 702434
rect 266360 697604 266412 697610
rect 266360 697546 266412 697552
rect 267648 697604 267700 697610
rect 267648 697546 267700 697552
rect 266372 450838 266400 697546
rect 276020 465724 276072 465730
rect 276020 465666 276072 465672
rect 276032 465118 276060 465666
rect 276020 465112 276072 465118
rect 276020 465054 276072 465060
rect 277308 465112 277360 465118
rect 277308 465054 277360 465060
rect 273260 464364 273312 464370
rect 273260 464306 273312 464312
rect 273272 463758 273300 464306
rect 273260 463752 273312 463758
rect 273260 463694 273312 463700
rect 274548 463752 274600 463758
rect 274548 463694 274600 463700
rect 266360 450832 266412 450838
rect 266360 450774 266412 450780
rect 271328 450832 271380 450838
rect 271328 450774 271380 450780
rect 255964 403640 256016 403646
rect 255964 403582 256016 403588
rect 253848 380996 253900 381002
rect 253848 380938 253900 380944
rect 253202 370424 253258 370433
rect 253202 370359 253258 370368
rect 251822 369064 251878 369073
rect 251822 368999 251878 369008
rect 250442 368384 250498 368393
rect 250442 368319 250498 368328
rect 250456 364334 250484 368319
rect 250456 364306 250576 364334
rect 249156 363656 249208 363662
rect 249156 363598 249208 363604
rect 250442 363624 250498 363633
rect 249168 295798 249196 363598
rect 250442 363559 250498 363568
rect 249800 317688 249852 317694
rect 249800 317630 249852 317636
rect 249812 312769 249840 317630
rect 249798 312760 249854 312769
rect 249798 312695 249854 312704
rect 250076 298104 250128 298110
rect 250076 298046 250128 298052
rect 250088 296886 250116 298046
rect 250076 296880 250128 296886
rect 250076 296822 250128 296828
rect 249156 295792 249208 295798
rect 249156 295734 249208 295740
rect 249706 291952 249762 291961
rect 249706 291887 249762 291896
rect 249064 291780 249116 291786
rect 249064 291722 249116 291728
rect 249076 290170 249104 291722
rect 249720 291310 249748 291887
rect 249708 291304 249760 291310
rect 249708 291246 249760 291252
rect 249076 290142 249196 290170
rect 249168 289898 249196 290142
rect 249168 289870 249366 289898
rect 249720 289884 249748 291246
rect 250088 289884 250116 296822
rect 250456 291553 250484 363559
rect 250548 298110 250576 364306
rect 250536 298104 250588 298110
rect 250536 298046 250588 298052
rect 251180 295452 251232 295458
rect 251180 295394 251232 295400
rect 251192 292233 251220 295394
rect 251178 292224 251234 292233
rect 251178 292159 251234 292168
rect 250442 291544 250498 291553
rect 250442 291479 250498 291488
rect 250456 289884 250484 291479
rect 250810 291136 250866 291145
rect 250810 291071 250866 291080
rect 250626 290048 250682 290057
rect 250626 289983 250682 289992
rect 250640 289898 250668 289983
rect 250824 289898 250852 291071
rect 250640 289884 250852 289898
rect 251192 289884 251220 292159
rect 251546 292088 251602 292097
rect 251546 292023 251602 292032
rect 251560 289884 251588 292023
rect 251836 290601 251864 368999
rect 251914 362264 251970 362273
rect 251914 362199 251970 362208
rect 251928 292097 251956 362199
rect 253216 298246 253244 370359
rect 253388 360868 253440 360874
rect 253388 360810 253440 360816
rect 253296 356720 253348 356726
rect 253296 356662 253348 356668
rect 253204 298240 253256 298246
rect 253204 298182 253256 298188
rect 253112 293480 253164 293486
rect 253112 293422 253164 293428
rect 252650 292360 252706 292369
rect 252650 292295 252706 292304
rect 251914 292088 251970 292097
rect 251914 292023 251970 292032
rect 251916 291780 251968 291786
rect 251916 291722 251968 291728
rect 251822 290592 251878 290601
rect 251822 290527 251878 290536
rect 251928 289921 251956 291722
rect 252098 290592 252154 290601
rect 252098 290527 252154 290536
rect 251914 289912 251970 289921
rect 250640 289870 250838 289884
rect 252112 289898 252140 290527
rect 252112 289870 252310 289898
rect 252664 289884 252692 292295
rect 252836 292120 252888 292126
rect 252836 292062 252888 292068
rect 252848 290494 252876 292062
rect 253124 291582 253152 293422
rect 253112 291576 253164 291582
rect 253112 291518 253164 291524
rect 252836 290488 252888 290494
rect 252836 290430 252888 290436
rect 252848 289898 252876 290430
rect 253216 289898 253244 298182
rect 253308 292369 253336 356662
rect 253400 298178 253428 360810
rect 253860 300778 253888 380938
rect 254124 378344 254176 378350
rect 254124 378286 254176 378292
rect 253860 300750 254072 300778
rect 254044 300150 254072 300750
rect 254032 300144 254084 300150
rect 254032 300086 254084 300092
rect 253388 298172 253440 298178
rect 253388 298114 253440 298120
rect 253400 296714 253428 298114
rect 253400 296686 253612 296714
rect 253294 292360 253350 292369
rect 253294 292295 253350 292304
rect 253584 289898 253612 296686
rect 254044 293078 254072 300086
rect 254032 293072 254084 293078
rect 254032 293014 254084 293020
rect 254136 290358 254164 378286
rect 255504 376848 255556 376854
rect 255504 376790 255556 376796
rect 255412 345704 255464 345710
rect 255412 345646 255464 345652
rect 255424 345098 255452 345646
rect 255412 345092 255464 345098
rect 255412 345034 255464 345040
rect 255424 301374 255452 345034
rect 255412 301368 255464 301374
rect 255412 301310 255464 301316
rect 255424 301034 255452 301310
rect 255412 301028 255464 301034
rect 255412 300970 255464 300976
rect 255412 300824 255464 300830
rect 255412 300766 255464 300772
rect 255424 299538 255452 300766
rect 255412 299532 255464 299538
rect 255412 299474 255464 299480
rect 254308 293072 254360 293078
rect 254308 293014 254360 293020
rect 254124 290352 254176 290358
rect 254124 290294 254176 290300
rect 252848 289870 253046 289898
rect 253216 289870 253414 289898
rect 253584 289870 253782 289898
rect 254136 289884 254164 290294
rect 254320 289898 254348 293014
rect 254860 291984 254912 291990
rect 254860 291926 254912 291932
rect 254320 289870 254518 289898
rect 254872 289884 254900 291926
rect 255044 291644 255096 291650
rect 255044 291586 255096 291592
rect 255056 290562 255084 291586
rect 255044 290556 255096 290562
rect 255044 290498 255096 290504
rect 255056 289898 255084 290498
rect 255424 289898 255452 299474
rect 255516 290086 255544 376790
rect 255976 300830 256004 403582
rect 266174 402112 266230 402121
rect 266174 402047 266230 402056
rect 262128 399628 262180 399634
rect 262128 399570 262180 399576
rect 256884 397520 256936 397526
rect 256884 397462 256936 397468
rect 256792 359508 256844 359514
rect 256792 359450 256844 359456
rect 256056 355360 256108 355366
rect 256056 355302 256108 355308
rect 255964 300824 256016 300830
rect 255964 300766 256016 300772
rect 256068 296714 256096 355302
rect 256148 301368 256200 301374
rect 256148 301310 256200 301316
rect 255976 296686 256096 296714
rect 255976 292398 256004 296686
rect 255964 292392 256016 292398
rect 255964 292334 256016 292340
rect 255504 290080 255556 290086
rect 255504 290022 255556 290028
rect 255056 289870 255254 289898
rect 255424 289870 255622 289898
rect 255976 289884 256004 292334
rect 256160 291310 256188 301310
rect 256700 299464 256752 299470
rect 256700 299406 256752 299412
rect 256712 291514 256740 299406
rect 256700 291508 256752 291514
rect 256700 291450 256752 291456
rect 256148 291304 256200 291310
rect 256148 291246 256200 291252
rect 256804 290290 256832 359450
rect 256896 297022 256924 397462
rect 260746 396808 260802 396817
rect 260746 396743 260802 396752
rect 260654 390008 260710 390017
rect 260654 389943 260710 389952
rect 259274 388376 259330 388385
rect 259274 388311 259330 388320
rect 259184 384328 259236 384334
rect 259184 384270 259236 384276
rect 258724 383716 258776 383722
rect 258724 383658 258776 383664
rect 257344 382288 257396 382294
rect 257344 382230 257396 382236
rect 257068 371272 257120 371278
rect 257068 371214 257120 371220
rect 257080 306374 257108 371214
rect 257080 306346 257292 306374
rect 256884 297016 256936 297022
rect 256884 296958 256936 296964
rect 256792 290284 256844 290290
rect 256792 290226 256844 290232
rect 256148 290080 256200 290086
rect 256148 290022 256200 290028
rect 256160 289898 256188 290022
rect 256896 289898 256924 296958
rect 257068 290284 257120 290290
rect 257068 290226 257120 290232
rect 256160 289870 256358 289898
rect 256726 289870 256924 289898
rect 257080 289884 257108 290226
rect 257264 290154 257292 306346
rect 257356 299470 257384 382230
rect 258264 319116 258316 319122
rect 258264 319058 258316 319064
rect 258276 306374 258304 319058
rect 258276 306346 258396 306374
rect 257344 299464 257396 299470
rect 257344 299406 257396 299412
rect 258172 291848 258224 291854
rect 258172 291790 258224 291796
rect 257804 291304 257856 291310
rect 257804 291246 257856 291252
rect 257252 290148 257304 290154
rect 257252 290090 257304 290096
rect 257436 290148 257488 290154
rect 257436 290090 257488 290096
rect 257448 289884 257476 290090
rect 257816 289884 257844 291246
rect 258184 289884 258212 291790
rect 258368 289898 258396 306346
rect 258736 291582 258764 383658
rect 258816 370524 258868 370530
rect 258816 370466 258868 370472
rect 258828 319122 258856 370466
rect 258816 319116 258868 319122
rect 258816 319058 258868 319064
rect 259196 318073 259224 384270
rect 259182 318064 259238 318073
rect 259182 317999 259238 318008
rect 259196 317966 259224 317999
rect 259184 317960 259236 317966
rect 259184 317902 259236 317908
rect 259288 311846 259316 388311
rect 260104 382356 260156 382362
rect 260104 382298 260156 382304
rect 259368 379568 259420 379574
rect 259368 379510 259420 379516
rect 259276 311840 259328 311846
rect 259276 311782 259328 311788
rect 258724 291576 258776 291582
rect 258724 291518 258776 291524
rect 258736 289898 258764 291518
rect 259276 291508 259328 291514
rect 259276 291450 259328 291456
rect 258368 289870 258566 289898
rect 258736 289870 258934 289898
rect 259288 289884 259316 291450
rect 259380 291242 259408 379510
rect 259736 378276 259788 378282
rect 259736 378218 259788 378224
rect 259552 302320 259604 302326
rect 259552 302262 259604 302268
rect 259564 293078 259592 302262
rect 259748 296714 259776 378218
rect 260116 299674 260144 382298
rect 260668 317014 260696 389943
rect 260656 317008 260708 317014
rect 260656 316950 260708 316956
rect 260196 309868 260248 309874
rect 260196 309810 260248 309816
rect 260208 302326 260236 309810
rect 260760 307630 260788 396743
rect 262034 389872 262090 389881
rect 262034 389807 262090 389816
rect 261944 388612 261996 388618
rect 261944 388554 261996 388560
rect 261484 383784 261536 383790
rect 261484 383726 261536 383732
rect 261300 375420 261352 375426
rect 261300 375362 261352 375368
rect 260748 307624 260800 307630
rect 260748 307566 260800 307572
rect 260760 306921 260788 307566
rect 260746 306912 260802 306921
rect 260746 306847 260802 306856
rect 261312 306374 261340 375362
rect 261312 306346 261432 306374
rect 260196 302320 260248 302326
rect 260196 302262 260248 302268
rect 259828 299668 259880 299674
rect 259828 299610 259880 299616
rect 260104 299668 260156 299674
rect 260104 299610 260156 299616
rect 259656 296686 259776 296714
rect 259552 293072 259604 293078
rect 259552 293014 259604 293020
rect 259368 291236 259420 291242
rect 259368 291178 259420 291184
rect 259380 290630 259408 291178
rect 259368 290624 259420 290630
rect 259368 290566 259420 290572
rect 259656 290222 259684 296686
rect 259644 290216 259696 290222
rect 259644 290158 259696 290164
rect 259656 289884 259684 290158
rect 259840 289898 259868 299610
rect 260196 293072 260248 293078
rect 260196 293014 260248 293020
rect 260208 289898 260236 293014
rect 261404 291394 261432 306346
rect 261496 300966 261524 383726
rect 261852 380180 261904 380186
rect 261852 380122 261904 380128
rect 261864 310298 261892 380122
rect 261956 310457 261984 388554
rect 261942 310448 261998 310457
rect 261942 310383 261998 310392
rect 261864 310270 261984 310298
rect 261956 307766 261984 310270
rect 261944 307760 261996 307766
rect 261944 307702 261996 307708
rect 261956 307222 261984 307702
rect 261944 307216 261996 307222
rect 261944 307158 261996 307164
rect 262048 301458 262076 389807
rect 262140 301578 262168 399570
rect 266082 391232 266138 391241
rect 266082 391167 266138 391176
rect 265992 389836 266044 389842
rect 265992 389778 266044 389784
rect 263416 388476 263468 388482
rect 263416 388418 263468 388424
rect 263324 387388 263376 387394
rect 263324 387330 263376 387336
rect 262956 385144 263008 385150
rect 262956 385086 263008 385092
rect 262864 380928 262916 380934
rect 262864 380870 262916 380876
rect 262496 302252 262548 302258
rect 262496 302194 262548 302200
rect 262128 301572 262180 301578
rect 262128 301514 262180 301520
rect 262048 301430 262168 301458
rect 261484 300960 261536 300966
rect 261484 300902 261536 300908
rect 261496 292534 261524 300902
rect 262140 300830 262168 301430
rect 262128 300824 262180 300830
rect 262128 300766 262180 300772
rect 262140 300218 262168 300766
rect 262128 300212 262180 300218
rect 262128 300154 262180 300160
rect 262508 293078 262536 302194
rect 262876 297158 262904 380870
rect 262968 302258 262996 385086
rect 263232 383036 263284 383042
rect 263232 382978 263284 382984
rect 263244 313274 263272 382978
rect 263336 315654 263364 387330
rect 263324 315648 263376 315654
rect 263324 315590 263376 315596
rect 263336 314265 263364 315590
rect 263322 314256 263378 314265
rect 263322 314191 263378 314200
rect 263232 313268 263284 313274
rect 263232 313210 263284 313216
rect 263244 312798 263272 313210
rect 263232 312792 263284 312798
rect 263232 312734 263284 312740
rect 263428 311778 263456 388418
rect 264888 387116 264940 387122
rect 264888 387058 264940 387064
rect 264336 385076 264388 385082
rect 264336 385018 264388 385024
rect 263508 378208 263560 378214
rect 263508 378150 263560 378156
rect 263048 311772 263100 311778
rect 263048 311714 263100 311720
rect 263416 311772 263468 311778
rect 263416 311714 263468 311720
rect 263060 311370 263088 311714
rect 263048 311364 263100 311370
rect 263048 311306 263100 311312
rect 262956 302252 263008 302258
rect 262956 302194 263008 302200
rect 263520 297634 263548 378150
rect 264244 376984 264296 376990
rect 264244 376926 264296 376932
rect 263876 305312 263928 305318
rect 263876 305254 263928 305260
rect 263888 305046 263916 305254
rect 263876 305040 263928 305046
rect 263876 304982 263928 304988
rect 263692 301368 263744 301374
rect 263692 301310 263744 301316
rect 263704 300898 263732 301310
rect 263692 300892 263744 300898
rect 263692 300834 263744 300840
rect 263508 297628 263560 297634
rect 263508 297570 263560 297576
rect 263520 297430 263548 297570
rect 263508 297424 263560 297430
rect 263508 297366 263560 297372
rect 262864 297152 262916 297158
rect 262864 297094 262916 297100
rect 262496 293072 262548 293078
rect 262496 293014 262548 293020
rect 261484 292528 261536 292534
rect 261484 292470 261536 292476
rect 262220 292528 262272 292534
rect 262220 292470 262272 292476
rect 261404 291366 261708 291394
rect 261116 291304 261168 291310
rect 261116 291246 261168 291252
rect 260748 291236 260800 291242
rect 260748 291178 260800 291184
rect 259840 289870 260038 289898
rect 260208 289870 260406 289898
rect 260760 289884 260788 291178
rect 261128 289884 261156 291246
rect 261484 291236 261536 291242
rect 261484 291178 261536 291184
rect 261496 289884 261524 291178
rect 261680 290018 261708 291366
rect 261668 290012 261720 290018
rect 261668 289954 261720 289960
rect 261680 289898 261708 289954
rect 261680 289870 261878 289898
rect 262232 289884 262260 292470
rect 262588 291372 262640 291378
rect 262588 291314 262640 291320
rect 262600 289884 262628 291314
rect 262876 289898 262904 297094
rect 263704 293078 263732 300834
rect 263140 293072 263192 293078
rect 263140 293014 263192 293020
rect 263692 293072 263744 293078
rect 263692 293014 263744 293020
rect 263152 289898 263180 293014
rect 263888 293010 263916 304982
rect 264060 297628 264112 297634
rect 264060 297570 264112 297576
rect 263876 293004 263928 293010
rect 263876 292946 263928 292952
rect 263692 291440 263744 291446
rect 263692 291382 263744 291388
rect 262876 289870 262982 289898
rect 263152 289870 263350 289898
rect 263704 289884 263732 291382
rect 264072 289884 264100 297570
rect 264256 296714 264284 376926
rect 264348 301374 264376 385018
rect 264704 379704 264756 379710
rect 264704 379646 264756 379652
rect 264428 379636 264480 379642
rect 264428 379578 264480 379584
rect 264336 301368 264388 301374
rect 264336 301310 264388 301316
rect 264440 298314 264468 379578
rect 264520 375760 264572 375766
rect 264520 375702 264572 375708
rect 264428 298308 264480 298314
rect 264428 298250 264480 298256
rect 264164 296686 264284 296714
rect 264164 291786 264192 296686
rect 264244 293072 264296 293078
rect 264244 293014 264296 293020
rect 264152 291780 264204 291786
rect 264152 291722 264204 291728
rect 264256 289898 264284 293014
rect 264440 292534 264468 298250
rect 264532 296070 264560 375702
rect 264612 370320 264664 370326
rect 264612 370262 264664 370268
rect 264520 296064 264572 296070
rect 264520 296006 264572 296012
rect 264624 293162 264652 370262
rect 264716 305318 264744 379646
rect 264900 310185 264928 387058
rect 265900 385892 265952 385898
rect 265900 385834 265952 385840
rect 265624 383852 265676 383858
rect 265624 383794 265676 383800
rect 264886 310176 264942 310185
rect 264886 310111 264942 310120
rect 264704 305312 264756 305318
rect 264704 305254 264756 305260
rect 264980 302184 265032 302190
rect 264980 302126 265032 302132
rect 264992 301510 265020 302126
rect 264980 301504 265032 301510
rect 264980 301446 265032 301452
rect 265636 300762 265664 383794
rect 265912 317218 265940 385834
rect 265900 317212 265952 317218
rect 265900 317154 265952 317160
rect 265912 312730 265940 317154
rect 265900 312724 265952 312730
rect 265900 312666 265952 312672
rect 266004 310078 266032 389778
rect 265992 310072 266044 310078
rect 265992 310014 266044 310020
rect 265716 309936 265768 309942
rect 265716 309878 265768 309884
rect 265728 305114 265756 309878
rect 266096 306338 266124 391167
rect 266188 307601 266216 402047
rect 269026 400616 269082 400625
rect 269026 400551 269082 400560
rect 266266 396672 266322 396681
rect 266266 396607 266322 396616
rect 266174 307592 266230 307601
rect 266174 307527 266230 307536
rect 266084 306332 266136 306338
rect 266084 306274 266136 306280
rect 266096 305930 266124 306274
rect 266084 305924 266136 305930
rect 266084 305866 266136 305872
rect 265716 305108 265768 305114
rect 265716 305050 265768 305056
rect 265072 300756 265124 300762
rect 265072 300698 265124 300704
rect 265624 300756 265676 300762
rect 265624 300698 265676 300704
rect 265084 299606 265112 300698
rect 265072 299600 265124 299606
rect 265072 299542 265124 299548
rect 264532 293134 264652 293162
rect 264428 292528 264480 292534
rect 264428 292470 264480 292476
rect 264532 292262 264560 293134
rect 264612 293004 264664 293010
rect 264612 292946 264664 292952
rect 264520 292256 264572 292262
rect 264520 292198 264572 292204
rect 264624 289898 264652 292946
rect 264980 292528 265032 292534
rect 264980 292470 265032 292476
rect 264992 289898 265020 292470
rect 265084 290170 265112 299542
rect 265084 290142 265388 290170
rect 265360 289898 265388 290142
rect 265728 289898 265756 305050
rect 266280 302190 266308 396607
rect 267002 395448 267058 395457
rect 267002 395383 267058 395392
rect 268476 395412 268528 395418
rect 266358 317384 266414 317393
rect 266358 317319 266414 317328
rect 266372 317082 266400 317319
rect 266360 317076 266412 317082
rect 266360 317018 266412 317024
rect 267016 305182 267044 395383
rect 268476 395354 268528 395360
rect 267372 393984 267424 393990
rect 267372 393926 267424 393932
rect 267096 375692 267148 375698
rect 267096 375634 267148 375640
rect 267004 305176 267056 305182
rect 267004 305118 267056 305124
rect 266268 302184 266320 302190
rect 266268 302126 266320 302132
rect 267108 291145 267136 375634
rect 267188 374740 267240 374746
rect 267188 374682 267240 374688
rect 267200 292330 267228 374682
rect 267280 374604 267332 374610
rect 267280 374546 267332 374552
rect 267292 294778 267320 374546
rect 267384 314702 267412 393926
rect 267556 393372 267608 393378
rect 267556 393314 267608 393320
rect 267568 317393 267596 393314
rect 267648 388544 267700 388550
rect 267648 388486 267700 388492
rect 267554 317384 267610 317393
rect 267554 317319 267610 317328
rect 267372 314696 267424 314702
rect 267372 314638 267424 314644
rect 267384 313585 267412 314638
rect 267370 313576 267426 313585
rect 267370 313511 267426 313520
rect 267660 311370 267688 388486
rect 268384 374808 268436 374814
rect 268384 374750 268436 374756
rect 267648 311364 267700 311370
rect 267648 311306 267700 311312
rect 267554 302832 267610 302841
rect 267554 302767 267610 302776
rect 267280 294772 267332 294778
rect 267280 294714 267332 294720
rect 267188 292324 267240 292330
rect 267188 292266 267240 292272
rect 267094 291136 267150 291145
rect 267094 291071 267150 291080
rect 264256 289870 264454 289898
rect 264624 289870 264822 289898
rect 264992 289870 265190 289898
rect 265360 289870 265558 289898
rect 265728 289870 265926 289898
rect 251914 289847 251970 289856
rect 248970 289640 249026 289649
rect 248800 289598 248970 289626
rect 248970 289575 249026 289584
rect 247038 289504 247094 289513
rect 247038 289439 247094 289448
rect 235540 289400 235592 289406
rect 235540 289342 235592 289348
rect 244004 289400 244056 289406
rect 244004 289342 244056 289348
rect 245568 289400 245620 289406
rect 245568 289342 245620 289348
rect 247498 289368 247554 289377
rect 247498 289303 247554 289312
rect 267568 247034 267596 302767
rect 268396 291106 268424 374750
rect 268488 325694 268516 395354
rect 268844 394120 268896 394126
rect 268658 394088 268714 394097
rect 268844 394062 268896 394068
rect 268658 394023 268714 394032
rect 268752 394052 268804 394058
rect 268488 325666 268608 325694
rect 268580 321774 268608 325666
rect 268568 321768 268620 321774
rect 268568 321710 268620 321716
rect 268580 317898 268608 321710
rect 268568 317892 268620 317898
rect 268568 317834 268620 317840
rect 268672 315790 268700 394023
rect 268752 393994 268804 394000
rect 268660 315784 268712 315790
rect 268660 315726 268712 315732
rect 268764 315722 268792 393994
rect 268752 315716 268804 315722
rect 268752 315658 268804 315664
rect 268764 315382 268792 315658
rect 268752 315376 268804 315382
rect 268752 315318 268804 315324
rect 268856 314537 268884 394062
rect 268936 392080 268988 392086
rect 268936 392022 268988 392028
rect 268842 314528 268898 314537
rect 268842 314463 268898 314472
rect 268948 304178 268976 392022
rect 269040 304881 269068 400551
rect 270314 398032 270370 398041
rect 270314 397967 270370 397976
rect 270132 396772 270184 396778
rect 270132 396714 270184 396720
rect 269856 392624 269908 392630
rect 269856 392566 269908 392572
rect 269670 387152 269726 387161
rect 269670 387087 269726 387096
rect 269578 385656 269634 385665
rect 269578 385591 269634 385600
rect 269304 318708 269356 318714
rect 269304 318650 269356 318656
rect 269026 304872 269082 304881
rect 269026 304807 269082 304816
rect 269040 304337 269068 304807
rect 269026 304328 269082 304337
rect 269026 304263 269082 304272
rect 268948 304150 269068 304178
rect 269040 303618 269068 304150
rect 269028 303612 269080 303618
rect 269028 303554 269080 303560
rect 269040 303006 269068 303554
rect 269028 303000 269080 303006
rect 269028 302942 269080 302948
rect 268384 291100 268436 291106
rect 268384 291042 268436 291048
rect 269028 287700 269080 287706
rect 269028 287642 269080 287648
rect 268396 285122 268976 285138
rect 268396 285116 268988 285122
rect 268396 285110 268936 285116
rect 267646 260128 267702 260137
rect 267646 260063 267702 260072
rect 267476 247006 267596 247034
rect 222476 242072 222528 242078
rect 222476 242014 222528 242020
rect 267476 240922 267504 247006
rect 267554 241904 267610 241913
rect 267554 241839 267610 241848
rect 267568 241398 267596 241839
rect 267556 241392 267608 241398
rect 267556 241334 267608 241340
rect 267556 241188 267608 241194
rect 267556 241130 267608 241136
rect 267568 240990 267596 241130
rect 267556 240984 267608 240990
rect 267556 240926 267608 240932
rect 267464 240916 267516 240922
rect 267464 240858 267516 240864
rect 222198 240680 222254 240689
rect 222198 240615 222254 240624
rect 222212 240514 222240 240615
rect 222200 240508 222252 240514
rect 222200 240450 222252 240456
rect 222028 240366 222148 240394
rect 222290 240408 222346 240417
rect 222200 240372 222252 240378
rect 222028 239358 222056 240366
rect 222290 240343 222292 240352
rect 222200 240314 222252 240320
rect 222344 240343 222346 240352
rect 222292 240314 222344 240320
rect 222106 240272 222162 240281
rect 222106 240207 222162 240216
rect 222016 239352 222068 239358
rect 222016 239294 222068 239300
rect 222028 238105 222056 239294
rect 222014 238096 222070 238105
rect 222014 238031 222070 238040
rect 222016 235952 222068 235958
rect 222016 235894 222068 235900
rect 222028 235550 222056 235894
rect 222016 235544 222068 235550
rect 222016 235486 222068 235492
rect 222028 233073 222056 235486
rect 222014 233064 222070 233073
rect 222014 232999 222070 233008
rect 221924 232688 221976 232694
rect 221924 232630 221976 232636
rect 221936 232393 221964 232630
rect 221922 232384 221978 232393
rect 221922 232319 221978 232328
rect 221832 230172 221884 230178
rect 221832 230114 221884 230120
rect 221740 212016 221792 212022
rect 221740 211958 221792 211964
rect 221844 155310 221872 230114
rect 222120 229498 222148 240207
rect 222212 240174 222240 240314
rect 267398 240230 267596 240258
rect 222200 240168 222252 240174
rect 222200 240110 222252 240116
rect 222534 239952 222562 240108
rect 222396 239924 222562 239952
rect 222292 239896 222344 239902
rect 222198 239864 222254 239873
rect 222292 239838 222344 239844
rect 222198 239799 222254 239808
rect 222108 229492 222160 229498
rect 222108 229434 222160 229440
rect 222016 225820 222068 225826
rect 222016 225762 222068 225768
rect 221832 155304 221884 155310
rect 221832 155246 221884 155252
rect 222028 144498 222056 225762
rect 221464 144492 221516 144498
rect 221464 144434 221516 144440
rect 222016 144492 222068 144498
rect 222016 144434 222068 144440
rect 222120 142934 222148 229434
rect 222212 218793 222240 239799
rect 222304 239714 222332 239838
rect 222396 239816 222424 239924
rect 222626 239816 222654 240108
rect 222718 239834 222746 240108
rect 222810 239902 222838 240108
rect 222902 239902 222930 240108
rect 222798 239896 222850 239902
rect 222890 239896 222942 239902
rect 222798 239838 222850 239844
rect 222888 239864 222890 239873
rect 222942 239864 222944 239873
rect 222396 239788 222516 239816
rect 222382 239728 222438 239737
rect 222304 239686 222382 239714
rect 222382 239663 222438 239672
rect 222292 239624 222344 239630
rect 222292 239566 222344 239572
rect 222198 218784 222254 218793
rect 222198 218719 222254 218728
rect 222304 180130 222332 239566
rect 222396 238678 222424 239663
rect 222384 238672 222436 238678
rect 222384 238614 222436 238620
rect 222488 237046 222516 239788
rect 222580 239788 222654 239816
rect 222706 239828 222758 239834
rect 222580 237114 222608 239788
rect 222888 239799 222944 239808
rect 222706 239770 222758 239776
rect 222994 239714 223022 240108
rect 223086 239970 223114 240108
rect 223074 239964 223126 239970
rect 223074 239906 223126 239912
rect 223178 239902 223206 240108
rect 223166 239896 223218 239902
rect 223166 239838 223218 239844
rect 223270 239816 223298 240108
rect 223362 239970 223390 240108
rect 223350 239964 223402 239970
rect 223350 239906 223402 239912
rect 223454 239902 223482 240108
rect 223442 239896 223494 239902
rect 223546 239873 223574 240108
rect 223638 239902 223666 240108
rect 223730 239970 223758 240108
rect 223718 239964 223770 239970
rect 223718 239906 223770 239912
rect 223626 239896 223678 239902
rect 223442 239838 223494 239844
rect 223532 239864 223588 239873
rect 223270 239788 223344 239816
rect 223822 239850 223850 240108
rect 223914 239970 223942 240108
rect 223902 239964 223954 239970
rect 223902 239906 223954 239912
rect 224006 239873 224034 240108
rect 224098 239970 224126 240108
rect 224190 239970 224218 240108
rect 224086 239964 224138 239970
rect 224086 239906 224138 239912
rect 224178 239964 224230 239970
rect 224178 239906 224230 239912
rect 224282 239902 224310 240108
rect 224270 239896 224322 239902
rect 223626 239838 223678 239844
rect 223532 239799 223588 239808
rect 223776 239822 223850 239850
rect 223992 239864 224048 239873
rect 223316 239748 223344 239788
rect 223672 239760 223724 239766
rect 223316 239720 223436 239748
rect 222752 239692 222804 239698
rect 222856 239686 223022 239714
rect 223120 239692 223172 239698
rect 222856 239680 222884 239686
rect 222804 239652 222884 239680
rect 222752 239634 222804 239640
rect 223120 239634 223172 239640
rect 222752 239556 222804 239562
rect 222752 239498 222804 239504
rect 222764 238338 222792 239498
rect 223132 239086 223160 239634
rect 223212 239624 223264 239630
rect 223212 239566 223264 239572
rect 223120 239080 223172 239086
rect 223120 239022 223172 239028
rect 223118 238912 223174 238921
rect 223118 238847 223174 238856
rect 223132 238678 223160 238847
rect 223120 238672 223172 238678
rect 223120 238614 223172 238620
rect 222752 238332 222804 238338
rect 222752 238274 222804 238280
rect 222936 238264 222988 238270
rect 222936 238206 222988 238212
rect 222568 237108 222620 237114
rect 222568 237050 222620 237056
rect 222476 237040 222528 237046
rect 222476 236982 222528 236988
rect 222844 237040 222896 237046
rect 222844 236982 222896 236988
rect 222292 180124 222344 180130
rect 222292 180066 222344 180072
rect 222200 144492 222252 144498
rect 222200 144434 222252 144440
rect 222108 142928 222160 142934
rect 222108 142870 222160 142876
rect 220082 141264 220138 141273
rect 220082 141199 220138 141208
rect 220084 137284 220136 137290
rect 220084 137226 220136 137232
rect 220096 136406 220124 137226
rect 219440 136400 219492 136406
rect 219440 136342 219492 136348
rect 220084 136400 220136 136406
rect 220084 136342 220136 136348
rect 219452 16574 219480 136342
rect 222212 16574 222240 144434
rect 222856 140350 222884 236982
rect 222948 143206 222976 238206
rect 223224 237998 223252 239566
rect 223408 239358 223436 239720
rect 223672 239702 223724 239708
rect 223488 239624 223540 239630
rect 223488 239566 223540 239572
rect 223580 239624 223632 239630
rect 223580 239566 223632 239572
rect 223500 239465 223528 239566
rect 223486 239456 223542 239465
rect 223486 239391 223542 239400
rect 223396 239352 223448 239358
rect 223396 239294 223448 239300
rect 223396 239216 223448 239222
rect 223396 239158 223448 239164
rect 223488 239216 223540 239222
rect 223488 239158 223540 239164
rect 223212 237992 223264 237998
rect 223212 237934 223264 237940
rect 223304 229152 223356 229158
rect 223304 229094 223356 229100
rect 223212 227248 223264 227254
rect 223212 227190 223264 227196
rect 223120 227180 223172 227186
rect 223120 227122 223172 227128
rect 223026 224360 223082 224369
rect 223026 224295 223082 224304
rect 222936 143200 222988 143206
rect 222936 143142 222988 143148
rect 222844 140344 222896 140350
rect 222844 140286 222896 140292
rect 223040 138553 223068 224295
rect 223132 141642 223160 227122
rect 223224 149802 223252 227190
rect 223316 154018 223344 229094
rect 223408 224954 223436 239158
rect 223500 238241 223528 239158
rect 223486 238232 223542 238241
rect 223486 238167 223542 238176
rect 223592 232665 223620 239566
rect 223684 238513 223712 239702
rect 223776 238950 223804 239822
rect 223992 239799 224048 239808
rect 224130 239864 224186 239873
rect 224374 239873 224402 240108
rect 224270 239838 224322 239844
rect 224360 239864 224416 239873
rect 224130 239799 224132 239808
rect 224184 239799 224186 239808
rect 224360 239799 224416 239808
rect 224466 239816 224494 240108
rect 224558 239970 224586 240108
rect 224546 239964 224598 239970
rect 224546 239906 224598 239912
rect 224650 239816 224678 240108
rect 224132 239770 224184 239776
rect 223948 239760 224000 239766
rect 223854 239728 223910 239737
rect 223948 239702 224000 239708
rect 224224 239760 224276 239766
rect 224374 239748 224402 239799
rect 224466 239788 224540 239816
rect 224374 239720 224448 239748
rect 224224 239702 224276 239708
rect 223854 239663 223856 239672
rect 223908 239663 223910 239672
rect 223856 239634 223908 239640
rect 223856 239556 223908 239562
rect 223856 239498 223908 239504
rect 223868 239222 223896 239498
rect 223856 239216 223908 239222
rect 223856 239158 223908 239164
rect 223764 238944 223816 238950
rect 223762 238912 223764 238921
rect 223856 238944 223908 238950
rect 223816 238912 223818 238921
rect 223856 238886 223908 238892
rect 223762 238847 223818 238856
rect 223776 238821 223804 238847
rect 223868 238814 223896 238886
rect 223856 238808 223908 238814
rect 223856 238750 223908 238756
rect 223670 238504 223726 238513
rect 223670 238439 223726 238448
rect 223670 238232 223726 238241
rect 223670 238167 223726 238176
rect 223578 232656 223634 232665
rect 223578 232591 223634 232600
rect 223580 229832 223632 229838
rect 223580 229774 223632 229780
rect 223408 224926 223528 224954
rect 223500 215966 223528 224926
rect 223488 215960 223540 215966
rect 223488 215902 223540 215908
rect 223592 213926 223620 229774
rect 223580 213920 223632 213926
rect 223580 213862 223632 213868
rect 223684 162217 223712 238167
rect 223960 236502 223988 239702
rect 224040 239692 224092 239698
rect 224040 239634 224092 239640
rect 223948 236496 224000 236502
rect 223948 236438 224000 236444
rect 223764 236428 223816 236434
rect 223764 236370 223816 236376
rect 223776 235890 223804 236370
rect 223764 235884 223816 235890
rect 223764 235826 223816 235832
rect 223776 229702 223804 235826
rect 223856 235748 223908 235754
rect 223856 235690 223908 235696
rect 223764 229696 223816 229702
rect 223764 229638 223816 229644
rect 223764 229560 223816 229566
rect 223764 229502 223816 229508
rect 223776 219337 223804 229502
rect 223868 220726 223896 235690
rect 224052 233234 224080 239634
rect 224052 233206 224172 233234
rect 224144 229786 224172 233206
rect 223960 229758 224172 229786
rect 223960 220794 223988 229758
rect 224040 229696 224092 229702
rect 224040 229638 224092 229644
rect 223948 220788 224000 220794
rect 223948 220730 224000 220736
rect 223856 220720 223908 220726
rect 223856 220662 223908 220668
rect 223762 219328 223818 219337
rect 223762 219263 223818 219272
rect 223670 162208 223726 162217
rect 223670 162143 223726 162152
rect 224052 159225 224080 229638
rect 224236 229566 224264 239702
rect 224316 239624 224368 239630
rect 224316 239566 224368 239572
rect 224328 238406 224356 239566
rect 224316 238400 224368 238406
rect 224316 238342 224368 238348
rect 224316 236496 224368 236502
rect 224316 236438 224368 236444
rect 224224 229560 224276 229566
rect 224224 229502 224276 229508
rect 224328 226273 224356 236438
rect 224420 231854 224448 239720
rect 224512 235754 224540 239788
rect 224604 239788 224678 239816
rect 224742 239816 224770 240108
rect 224834 239970 224862 240108
rect 224822 239964 224874 239970
rect 224822 239906 224874 239912
rect 224926 239873 224954 240108
rect 224912 239864 224968 239873
rect 224742 239788 224816 239816
rect 224912 239799 224968 239808
rect 224604 237697 224632 239788
rect 224684 239692 224736 239698
rect 224684 239634 224736 239640
rect 224590 237688 224646 237697
rect 224590 237623 224646 237632
rect 224500 235748 224552 235754
rect 224500 235690 224552 235696
rect 224420 231826 224540 231854
rect 224512 229537 224540 231826
rect 224498 229528 224554 229537
rect 224498 229463 224554 229472
rect 224498 229392 224554 229401
rect 224498 229327 224554 229336
rect 224408 226976 224460 226982
rect 224408 226918 224460 226924
rect 224314 226264 224370 226273
rect 224314 226199 224370 226208
rect 224222 224496 224278 224505
rect 224222 224431 224278 224440
rect 224038 159216 224094 159225
rect 224038 159151 224094 159160
rect 223304 154012 223356 154018
rect 223304 153954 223356 153960
rect 223212 149796 223264 149802
rect 223212 149738 223264 149744
rect 224236 142769 224264 224431
rect 224316 220788 224368 220794
rect 224316 220730 224368 220736
rect 224328 220658 224356 220730
rect 224316 220652 224368 220658
rect 224316 220594 224368 220600
rect 224328 143342 224356 220594
rect 224420 170377 224448 226918
rect 224512 222194 224540 229327
rect 224604 226982 224632 237623
rect 224696 236570 224724 239634
rect 224684 236564 224736 236570
rect 224684 236506 224736 236512
rect 224788 233234 224816 239788
rect 225018 239748 225046 240108
rect 225110 239873 225138 240108
rect 225096 239864 225152 239873
rect 225096 239799 225152 239808
rect 225202 239748 225230 240108
rect 225294 239970 225322 240108
rect 225282 239964 225334 239970
rect 225282 239906 225334 239912
rect 225386 239816 225414 240108
rect 225478 239970 225506 240108
rect 225570 239970 225598 240108
rect 225466 239964 225518 239970
rect 225466 239906 225518 239912
rect 225558 239964 225610 239970
rect 225558 239906 225610 239912
rect 225662 239850 225690 240108
rect 225754 239970 225782 240108
rect 225846 239970 225874 240108
rect 225742 239964 225794 239970
rect 225742 239906 225794 239912
rect 225834 239964 225886 239970
rect 225834 239906 225886 239912
rect 225616 239822 225690 239850
rect 225786 239864 225842 239873
rect 225386 239788 225460 239816
rect 225018 239720 225092 239748
rect 224868 239692 224920 239698
rect 224868 239634 224920 239640
rect 224880 238542 224908 239634
rect 225064 239562 225092 239720
rect 225156 239720 225368 239748
rect 225052 239556 225104 239562
rect 225052 239498 225104 239504
rect 225156 239442 225184 239720
rect 225236 239624 225288 239630
rect 225236 239566 225288 239572
rect 225064 239414 225184 239442
rect 224960 239216 225012 239222
rect 224960 239158 225012 239164
rect 224868 238536 224920 238542
rect 224868 238478 224920 238484
rect 224868 236564 224920 236570
rect 224868 236506 224920 236512
rect 224696 233206 224816 233234
rect 224592 226976 224644 226982
rect 224592 226918 224644 226924
rect 224512 222166 224632 222194
rect 224500 220720 224552 220726
rect 224500 220662 224552 220668
rect 224512 220522 224540 220662
rect 224500 220516 224552 220522
rect 224500 220458 224552 220464
rect 224406 170368 224462 170377
rect 224406 170303 224462 170312
rect 224512 160954 224540 220458
rect 224604 200802 224632 222166
rect 224696 216646 224724 233206
rect 224880 229838 224908 236506
rect 224868 229832 224920 229838
rect 224868 229774 224920 229780
rect 224972 217977 225000 239158
rect 225064 224233 225092 239414
rect 225050 224224 225106 224233
rect 225050 224159 225106 224168
rect 225248 223574 225276 239566
rect 225340 239465 225368 239720
rect 225326 239456 225382 239465
rect 225326 239391 225382 239400
rect 225432 237640 225460 239788
rect 225512 239556 225564 239562
rect 225512 239498 225564 239504
rect 225524 239329 225552 239498
rect 225510 239320 225566 239329
rect 225510 239255 225566 239264
rect 225616 237998 225644 239822
rect 225938 239850 225966 240108
rect 226030 239970 226058 240108
rect 226018 239964 226070 239970
rect 226018 239906 226070 239912
rect 225786 239799 225842 239808
rect 225892 239822 225966 239850
rect 225800 239630 225828 239799
rect 225788 239624 225840 239630
rect 225694 239592 225750 239601
rect 225788 239566 225840 239572
rect 225694 239527 225696 239536
rect 225748 239527 225750 239536
rect 225696 239498 225748 239504
rect 225708 239222 225736 239498
rect 225696 239216 225748 239222
rect 225696 239158 225748 239164
rect 225604 237992 225656 237998
rect 225604 237934 225656 237940
rect 225432 237612 225552 237640
rect 225420 237516 225472 237522
rect 225420 237458 225472 237464
rect 225432 237386 225460 237458
rect 225420 237380 225472 237386
rect 225420 237322 225472 237328
rect 225418 225992 225474 226001
rect 225418 225927 225474 225936
rect 225156 223546 225276 223574
rect 224958 217968 225014 217977
rect 224958 217903 225014 217912
rect 224684 216640 224736 216646
rect 224684 216582 224736 216588
rect 224592 200796 224644 200802
rect 224592 200738 224644 200744
rect 225156 199442 225184 223546
rect 225144 199436 225196 199442
rect 225144 199378 225196 199384
rect 224500 160948 224552 160954
rect 224500 160890 224552 160896
rect 225432 146946 225460 225927
rect 225524 218006 225552 237612
rect 225616 231305 225644 237934
rect 225694 237552 225750 237561
rect 225694 237487 225750 237496
rect 225602 231296 225658 231305
rect 225602 231231 225658 231240
rect 225512 218000 225564 218006
rect 225512 217942 225564 217948
rect 225604 155508 225656 155514
rect 225604 155450 225656 155456
rect 225420 146940 225472 146946
rect 225420 146882 225472 146888
rect 224316 143336 224368 143342
rect 224316 143278 224368 143284
rect 224222 142760 224278 142769
rect 224222 142695 224278 142704
rect 223120 141636 223172 141642
rect 223120 141578 223172 141584
rect 223026 138544 223082 138553
rect 223026 138479 223082 138488
rect 223580 135924 223632 135930
rect 223580 135866 223632 135872
rect 218164 16546 219296 16574
rect 219452 16546 220032 16574
rect 222212 16546 222792 16574
rect 217324 3800 217376 3806
rect 217324 3742 217376 3748
rect 218060 3120 218112 3126
rect 218060 3062 218112 3068
rect 218072 480 218100 3062
rect 219268 480 219296 16546
rect 215638 354 215750 480
rect 215312 326 215750 354
rect 215638 -960 215750 326
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220004 354 220032 16546
rect 221556 4004 221608 4010
rect 221556 3946 221608 3952
rect 221568 480 221596 3946
rect 222764 480 222792 16546
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 220422 -960 220534 326
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223592 354 223620 135866
rect 225144 3936 225196 3942
rect 225144 3878 225196 3884
rect 225156 480 225184 3878
rect 225616 3058 225644 155450
rect 225708 140418 225736 237487
rect 225892 236337 225920 239822
rect 226122 239816 226150 240108
rect 226076 239788 226150 239816
rect 226214 239816 226242 240108
rect 226306 239970 226334 240108
rect 226294 239964 226346 239970
rect 226294 239906 226346 239912
rect 226398 239850 226426 240108
rect 226490 239902 226518 240108
rect 226352 239822 226426 239850
rect 226478 239896 226530 239902
rect 226582 239873 226610 240108
rect 226674 239902 226702 240108
rect 226662 239896 226714 239902
rect 226478 239838 226530 239844
rect 226568 239864 226624 239873
rect 226214 239788 226288 239816
rect 226076 239748 226104 239788
rect 226030 239720 226104 239748
rect 226030 239680 226058 239720
rect 226260 239680 226288 239788
rect 226030 239652 226104 239680
rect 225972 239148 226024 239154
rect 225972 239090 226024 239096
rect 225984 238678 226012 239090
rect 225972 238672 226024 238678
rect 225972 238614 226024 238620
rect 226076 236502 226104 239652
rect 226168 239652 226288 239680
rect 226064 236496 226116 236502
rect 226064 236438 226116 236444
rect 225878 236328 225934 236337
rect 225878 236263 225934 236272
rect 226168 235906 226196 239652
rect 226352 239612 226380 239822
rect 226662 239838 226714 239844
rect 226568 239799 226624 239808
rect 226432 239760 226484 239766
rect 226432 239702 226484 239708
rect 226570 239760 226622 239766
rect 226766 239748 226794 240108
rect 226858 239970 226886 240108
rect 226846 239964 226898 239970
rect 226846 239906 226898 239912
rect 226950 239748 226978 240108
rect 226622 239720 226702 239748
rect 226766 239720 226840 239748
rect 226570 239702 226622 239708
rect 226260 239584 226380 239612
rect 226260 237250 226288 239584
rect 226444 239544 226472 239702
rect 226674 239612 226702 239720
rect 226352 239516 226472 239544
rect 226522 239592 226578 239601
rect 226522 239527 226578 239536
rect 226628 239584 226702 239612
rect 226248 237244 226300 237250
rect 226248 237186 226300 237192
rect 226352 236434 226380 239516
rect 226432 239420 226484 239426
rect 226432 239362 226484 239368
rect 226444 238746 226472 239362
rect 226432 238740 226484 238746
rect 226432 238682 226484 238688
rect 226536 237250 226564 239527
rect 226628 239057 226656 239584
rect 226614 239048 226670 239057
rect 226614 238983 226670 238992
rect 226614 238232 226670 238241
rect 226614 238167 226670 238176
rect 226628 237794 226656 238167
rect 226616 237788 226668 237794
rect 226616 237730 226668 237736
rect 226708 237788 226760 237794
rect 226708 237730 226760 237736
rect 226616 237584 226668 237590
rect 226616 237526 226668 237532
rect 226524 237244 226576 237250
rect 226524 237186 226576 237192
rect 226340 236428 226392 236434
rect 226340 236370 226392 236376
rect 226432 236156 226484 236162
rect 226432 236098 226484 236104
rect 226076 235878 226196 235906
rect 226076 229022 226104 235878
rect 226156 235748 226208 235754
rect 226156 235690 226208 235696
rect 226064 229016 226116 229022
rect 226064 228958 226116 228964
rect 226168 224954 226196 235690
rect 225892 224926 226196 224954
rect 225786 224224 225842 224233
rect 225786 224159 225842 224168
rect 225800 142633 225828 224159
rect 225892 220250 225920 224926
rect 226248 224256 226300 224262
rect 226248 224198 226300 224204
rect 225880 220244 225932 220250
rect 225880 220186 225932 220192
rect 225786 142624 225842 142633
rect 225786 142559 225842 142568
rect 225892 140593 225920 220186
rect 225878 140584 225934 140593
rect 225878 140519 225934 140528
rect 225696 140412 225748 140418
rect 225696 140354 225748 140360
rect 226260 139126 226288 224198
rect 226444 220454 226472 236098
rect 226522 235920 226578 235929
rect 226522 235855 226578 235864
rect 226536 235754 226564 235855
rect 226524 235748 226576 235754
rect 226524 235690 226576 235696
rect 226524 233300 226576 233306
rect 226524 233242 226576 233248
rect 226432 220448 226484 220454
rect 226432 220390 226484 220396
rect 226536 220318 226564 233242
rect 226628 229090 226656 237526
rect 226616 229084 226668 229090
rect 226616 229026 226668 229032
rect 226524 220312 226576 220318
rect 226524 220254 226576 220260
rect 226720 217326 226748 237730
rect 226812 237368 226840 239720
rect 226904 239720 226978 239748
rect 227042 239737 227070 240108
rect 227028 239728 227084 239737
rect 226904 237590 226932 239720
rect 227028 239663 227084 239672
rect 227134 239680 227162 240108
rect 227226 239748 227254 240108
rect 227318 239850 227346 240108
rect 227410 239970 227438 240108
rect 227398 239964 227450 239970
rect 227398 239906 227450 239912
rect 227318 239822 227392 239850
rect 227226 239720 227300 239748
rect 227134 239652 227208 239680
rect 226984 239624 227036 239630
rect 226984 239566 227036 239572
rect 226996 239465 227024 239566
rect 227076 239488 227128 239494
rect 226982 239456 227038 239465
rect 227076 239430 227128 239436
rect 226982 239391 227038 239400
rect 226982 239048 227038 239057
rect 226982 238983 227038 238992
rect 226996 238542 227024 238983
rect 226984 238536 227036 238542
rect 226984 238478 227036 238484
rect 227088 237794 227116 239430
rect 227076 237788 227128 237794
rect 227076 237730 227128 237736
rect 226892 237584 226944 237590
rect 226892 237526 226944 237532
rect 226812 237340 226932 237368
rect 226800 237244 226852 237250
rect 226800 237186 226852 237192
rect 226812 217841 226840 237186
rect 226904 230489 226932 237340
rect 226984 237176 227036 237182
rect 226984 237118 227036 237124
rect 226890 230480 226946 230489
rect 226890 230415 226946 230424
rect 226798 217832 226854 217841
rect 226798 217767 226854 217776
rect 226708 217320 226760 217326
rect 226708 217262 226760 217268
rect 226996 145654 227024 237118
rect 227076 235136 227128 235142
rect 227076 235078 227128 235084
rect 226984 145648 227036 145654
rect 226984 145590 227036 145596
rect 227088 144906 227116 235078
rect 227180 231849 227208 239652
rect 227272 237833 227300 239720
rect 227258 237824 227314 237833
rect 227258 237759 227314 237768
rect 227364 233306 227392 239822
rect 227502 239816 227530 240108
rect 227594 239970 227622 240108
rect 227582 239964 227634 239970
rect 227582 239906 227634 239912
rect 227686 239873 227714 240108
rect 227672 239864 227728 239873
rect 227502 239788 227576 239816
rect 227672 239799 227728 239808
rect 227442 239728 227498 239737
rect 227442 239663 227444 239672
rect 227496 239663 227498 239672
rect 227444 239634 227496 239640
rect 227444 239488 227496 239494
rect 227442 239456 227444 239465
rect 227496 239456 227498 239465
rect 227442 239391 227498 239400
rect 227444 237788 227496 237794
rect 227444 237730 227496 237736
rect 227456 235074 227484 237730
rect 227444 235068 227496 235074
rect 227444 235010 227496 235016
rect 227352 233300 227404 233306
rect 227352 233242 227404 233248
rect 227166 231840 227222 231849
rect 227166 231775 227222 231784
rect 227168 229628 227220 229634
rect 227168 229570 227220 229576
rect 227180 148238 227208 229570
rect 227352 223644 227404 223650
rect 227352 223586 227404 223592
rect 227260 220312 227312 220318
rect 227260 220254 227312 220260
rect 227168 148232 227220 148238
rect 227168 148174 227220 148180
rect 227076 144900 227128 144906
rect 227076 144842 227128 144848
rect 227272 140486 227300 220254
rect 227364 148306 227392 223586
rect 227444 220788 227496 220794
rect 227444 220730 227496 220736
rect 227456 220454 227484 220730
rect 227444 220448 227496 220454
rect 227444 220390 227496 220396
rect 227456 160818 227484 220390
rect 227548 215286 227576 239788
rect 227778 239748 227806 240108
rect 227870 239816 227898 240108
rect 227962 239970 227990 240108
rect 228054 239970 228082 240108
rect 227950 239964 228002 239970
rect 227950 239906 228002 239912
rect 228042 239964 228094 239970
rect 228042 239906 228094 239912
rect 228146 239873 228174 240108
rect 228238 239970 228266 240108
rect 228226 239964 228278 239970
rect 228226 239906 228278 239912
rect 228132 239864 228188 239873
rect 227870 239788 227944 239816
rect 228330 239816 228358 240108
rect 228422 239970 228450 240108
rect 228514 239970 228542 240108
rect 228410 239964 228462 239970
rect 228410 239906 228462 239912
rect 228502 239964 228554 239970
rect 228502 239906 228554 239912
rect 228606 239902 228634 240108
rect 228698 239902 228726 240108
rect 228790 239902 228818 240108
rect 228594 239896 228646 239902
rect 228132 239799 228188 239808
rect 227732 239720 227806 239748
rect 227628 239624 227680 239630
rect 227628 239566 227680 239572
rect 227640 236162 227668 239566
rect 227732 238950 227760 239720
rect 227916 239680 227944 239788
rect 228284 239788 228358 239816
rect 228454 239864 228510 239873
rect 228594 239838 228646 239844
rect 228686 239896 228738 239902
rect 228686 239838 228738 239844
rect 228778 239896 228830 239902
rect 228778 239838 228830 239844
rect 228454 239799 228510 239808
rect 227824 239652 227944 239680
rect 227994 239728 228050 239737
rect 227994 239663 228050 239672
rect 228088 239692 228140 239698
rect 227720 238944 227772 238950
rect 227720 238886 227772 238892
rect 227824 236638 227852 239652
rect 227904 239420 227956 239426
rect 227904 239362 227956 239368
rect 227916 239222 227944 239362
rect 227904 239216 227956 239222
rect 227904 239158 227956 239164
rect 228008 238950 228036 239663
rect 228140 239652 228220 239680
rect 228088 239634 228140 239640
rect 228088 239488 228140 239494
rect 228088 239430 228140 239436
rect 228100 239086 228128 239430
rect 228192 239329 228220 239652
rect 228178 239320 228234 239329
rect 228178 239255 228234 239264
rect 228180 239216 228232 239222
rect 228180 239158 228232 239164
rect 228088 239080 228140 239086
rect 228088 239022 228140 239028
rect 227996 238944 228048 238950
rect 227996 238886 228048 238892
rect 227994 238776 228050 238785
rect 227994 238711 228050 238720
rect 227904 238332 227956 238338
rect 227904 238274 227956 238280
rect 227812 236632 227864 236638
rect 227812 236574 227864 236580
rect 227628 236156 227680 236162
rect 227628 236098 227680 236104
rect 227720 227860 227772 227866
rect 227720 227802 227772 227808
rect 227536 215280 227588 215286
rect 227536 215222 227588 215228
rect 227732 211993 227760 227802
rect 227916 217569 227944 238274
rect 228008 238184 228036 238711
rect 228100 238338 228128 239022
rect 228088 238332 228140 238338
rect 228088 238274 228140 238280
rect 228008 238156 228128 238184
rect 227996 236632 228048 236638
rect 227996 236574 228048 236580
rect 227902 217560 227958 217569
rect 227902 217495 227958 217504
rect 227718 211984 227774 211993
rect 227718 211919 227774 211928
rect 227444 160812 227496 160818
rect 227444 160754 227496 160760
rect 227352 148300 227404 148306
rect 227352 148242 227404 148248
rect 227260 140480 227312 140486
rect 227260 140422 227312 140428
rect 228008 139194 228036 236574
rect 228100 161809 228128 238156
rect 228192 234394 228220 239158
rect 228180 234388 228232 234394
rect 228180 234330 228232 234336
rect 228284 231928 228312 239788
rect 228362 239728 228418 239737
rect 228362 239663 228418 239672
rect 228376 239562 228404 239663
rect 228364 239556 228416 239562
rect 228364 239498 228416 239504
rect 228376 232529 228404 239498
rect 228468 235793 228496 239799
rect 228640 239760 228692 239766
rect 228640 239702 228692 239708
rect 228548 239624 228600 239630
rect 228652 239601 228680 239702
rect 228882 239680 228910 240108
rect 228974 239816 229002 240108
rect 229066 239970 229094 240108
rect 229158 239970 229186 240108
rect 229054 239964 229106 239970
rect 229054 239906 229106 239912
rect 229146 239964 229198 239970
rect 229146 239906 229198 239912
rect 229250 239873 229278 240108
rect 229236 239864 229292 239873
rect 228974 239788 229048 239816
rect 229236 239799 229292 239808
rect 229342 239816 229370 240108
rect 229434 239970 229462 240108
rect 229526 239970 229554 240108
rect 229618 239970 229646 240108
rect 229422 239964 229474 239970
rect 229422 239906 229474 239912
rect 229514 239964 229566 239970
rect 229514 239906 229566 239912
rect 229606 239964 229658 239970
rect 229606 239906 229658 239912
rect 229710 239850 229738 240108
rect 229802 239873 229830 240108
rect 229894 239902 229922 240108
rect 229986 239970 230014 240108
rect 229974 239964 230026 239970
rect 229974 239906 230026 239912
rect 229882 239896 229934 239902
rect 229468 239828 229520 239834
rect 229342 239788 229416 239816
rect 228882 239652 228956 239680
rect 228548 239566 228600 239572
rect 228638 239592 228694 239601
rect 228454 235784 228510 235793
rect 228454 235719 228510 235728
rect 228560 232778 228588 239566
rect 228638 239527 228694 239536
rect 228640 239488 228692 239494
rect 228640 239430 228692 239436
rect 228822 239456 228878 239465
rect 228468 232750 228588 232778
rect 228362 232520 228418 232529
rect 228362 232455 228418 232464
rect 228192 231900 228312 231928
rect 228192 228993 228220 231900
rect 228468 231854 228496 232750
rect 228548 232620 228600 232626
rect 228548 232562 228600 232568
rect 228284 231826 228496 231854
rect 228178 228984 228234 228993
rect 228178 228919 228234 228928
rect 228284 218822 228312 231826
rect 228456 227384 228508 227390
rect 228456 227326 228508 227332
rect 228272 218816 228324 218822
rect 228272 218758 228324 218764
rect 228086 161800 228142 161809
rect 228086 161735 228142 161744
rect 228364 153740 228416 153746
rect 228364 153682 228416 153688
rect 227996 139188 228048 139194
rect 227996 139130 228048 139136
rect 226248 139120 226300 139126
rect 226248 139062 226300 139068
rect 226260 138122 226288 139062
rect 226260 138094 226380 138122
rect 225604 3052 225656 3058
rect 225604 2994 225656 3000
rect 226352 480 226380 138094
rect 226430 121000 226486 121009
rect 226430 120935 226486 120944
rect 226444 16574 226472 120935
rect 226444 16546 227576 16574
rect 227548 480 227576 16546
rect 228376 3942 228404 153682
rect 228468 142905 228496 227326
rect 228560 154290 228588 232562
rect 228652 227866 228680 239430
rect 228732 239420 228784 239426
rect 228822 239391 228878 239400
rect 228732 239362 228784 239368
rect 228744 231810 228772 239362
rect 228836 239086 228864 239391
rect 228824 239080 228876 239086
rect 228824 239022 228876 239028
rect 228928 238456 228956 239652
rect 229020 239426 229048 239788
rect 229100 239760 229152 239766
rect 229100 239702 229152 239708
rect 229282 239728 229338 239737
rect 229112 239426 229140 239702
rect 229192 239692 229244 239698
rect 229282 239663 229284 239672
rect 229192 239634 229244 239640
rect 229336 239663 229338 239672
rect 229284 239634 229336 239640
rect 229008 239420 229060 239426
rect 229008 239362 229060 239368
rect 229100 239420 229152 239426
rect 229100 239362 229152 239368
rect 228928 238428 229048 238456
rect 228916 238332 228968 238338
rect 228916 238274 228968 238280
rect 228732 231804 228784 231810
rect 228732 231746 228784 231752
rect 228732 229696 228784 229702
rect 228732 229638 228784 229644
rect 228640 227860 228692 227866
rect 228640 227802 228692 227808
rect 228640 221536 228692 221542
rect 228640 221478 228692 221484
rect 228548 154284 228600 154290
rect 228548 154226 228600 154232
rect 228652 144294 228680 221478
rect 228744 152590 228772 229638
rect 228928 229094 228956 238274
rect 229020 233238 229048 238428
rect 229112 237182 229140 239362
rect 229204 238785 229232 239634
rect 229282 239592 229338 239601
rect 229282 239527 229284 239536
rect 229336 239527 229338 239536
rect 229284 239498 229336 239504
rect 229190 238776 229246 238785
rect 229190 238711 229246 238720
rect 229296 238474 229324 239498
rect 229284 238468 229336 238474
rect 229284 238410 229336 238416
rect 229388 238377 229416 239788
rect 229468 239770 229520 239776
rect 229664 239822 229738 239850
rect 229788 239864 229844 239873
rect 229480 239737 229508 239770
rect 229466 239728 229522 239737
rect 229466 239663 229522 239672
rect 229664 239630 229692 239822
rect 230078 239850 230106 240108
rect 229882 239838 229934 239844
rect 229788 239799 229844 239808
rect 230032 239822 230106 239850
rect 229744 239760 229796 239766
rect 229744 239702 229796 239708
rect 229652 239624 229704 239630
rect 229558 239592 229614 239601
rect 229652 239566 229704 239572
rect 229558 239527 229614 239536
rect 229468 239012 229520 239018
rect 229468 238954 229520 238960
rect 229374 238368 229430 238377
rect 229374 238303 229430 238312
rect 229376 237448 229428 237454
rect 229376 237390 229428 237396
rect 229284 237380 229336 237386
rect 229284 237322 229336 237328
rect 229100 237176 229152 237182
rect 229100 237118 229152 237124
rect 229100 236632 229152 236638
rect 229100 236574 229152 236580
rect 229008 233232 229060 233238
rect 229008 233174 229060 233180
rect 229112 231854 229140 236574
rect 229112 231826 229232 231854
rect 228928 229066 229048 229094
rect 228916 219360 228968 219366
rect 228916 219302 228968 219308
rect 228928 218822 228956 219302
rect 228916 218816 228968 218822
rect 228916 218758 228968 218764
rect 229020 203590 229048 229066
rect 229204 219434 229232 231826
rect 229296 220318 229324 237322
rect 229388 222970 229416 237390
rect 229376 222964 229428 222970
rect 229376 222906 229428 222912
rect 229284 220312 229336 220318
rect 229284 220254 229336 220260
rect 229296 220114 229324 220254
rect 229284 220108 229336 220114
rect 229284 220050 229336 220056
rect 229192 219428 229244 219434
rect 229192 219370 229244 219376
rect 229008 203584 229060 203590
rect 229008 203526 229060 203532
rect 229020 200114 229048 203526
rect 228836 200086 229048 200114
rect 228732 152584 228784 152590
rect 228732 152526 228784 152532
rect 228836 149054 228864 200086
rect 229100 151020 229152 151026
rect 229100 150962 229152 150968
rect 228824 149048 228876 149054
rect 228824 148990 228876 148996
rect 228640 144288 228692 144294
rect 228640 144230 228692 144236
rect 228454 142896 228510 142905
rect 228454 142831 228510 142840
rect 229112 16574 229140 150962
rect 229480 140622 229508 238954
rect 229572 161294 229600 239527
rect 229664 237810 229692 239566
rect 229756 238377 229784 239702
rect 229836 239692 229888 239698
rect 229836 239634 229888 239640
rect 229928 239692 229980 239698
rect 229928 239634 229980 239640
rect 229848 239086 229876 239634
rect 229836 239080 229888 239086
rect 229836 239022 229888 239028
rect 229742 238368 229798 238377
rect 229742 238303 229798 238312
rect 229756 237969 229784 238303
rect 229742 237960 229798 237969
rect 229742 237895 229798 237904
rect 229664 237782 229784 237810
rect 229650 237280 229706 237289
rect 229650 237215 229706 237224
rect 229664 236201 229692 237215
rect 229650 236192 229706 236201
rect 229650 236127 229706 236136
rect 229650 236056 229706 236065
rect 229650 235991 229706 236000
rect 229664 217433 229692 235991
rect 229756 233234 229784 237782
rect 229848 236450 229876 239022
rect 229940 236609 229968 239634
rect 230032 239465 230060 239822
rect 230170 239680 230198 240108
rect 230262 239970 230290 240108
rect 230250 239964 230302 239970
rect 230250 239906 230302 239912
rect 230354 239873 230382 240108
rect 230340 239864 230396 239873
rect 230446 239850 230474 240108
rect 230538 239970 230566 240108
rect 230526 239964 230578 239970
rect 230526 239906 230578 239912
rect 230446 239822 230520 239850
rect 230340 239799 230396 239808
rect 230388 239760 230440 239766
rect 230124 239652 230198 239680
rect 230294 239728 230350 239737
rect 230388 239702 230440 239708
rect 230294 239663 230350 239672
rect 230018 239456 230074 239465
rect 230018 239391 230074 239400
rect 230032 237046 230060 239391
rect 230124 237454 230152 239652
rect 230308 239630 230336 239663
rect 230296 239624 230348 239630
rect 230296 239566 230348 239572
rect 230204 239556 230256 239562
rect 230204 239498 230256 239504
rect 230112 237448 230164 237454
rect 230112 237390 230164 237396
rect 230216 237386 230244 239498
rect 230296 239488 230348 239494
rect 230294 239456 230296 239465
rect 230348 239456 230350 239465
rect 230294 239391 230350 239400
rect 230400 238270 230428 239702
rect 230388 238264 230440 238270
rect 230388 238206 230440 238212
rect 230492 237538 230520 239822
rect 230630 239748 230658 240108
rect 230400 237510 230520 237538
rect 230584 239720 230658 239748
rect 230204 237380 230256 237386
rect 230204 237322 230256 237328
rect 230020 237040 230072 237046
rect 230020 236982 230072 236988
rect 229926 236600 229982 236609
rect 229926 236535 229982 236544
rect 229848 236422 229968 236450
rect 229940 233234 229968 236422
rect 230400 234614 230428 237510
rect 230478 235784 230534 235793
rect 230478 235719 230534 235728
rect 230492 235550 230520 235719
rect 230480 235544 230532 235550
rect 230480 235486 230532 235492
rect 230216 234586 230428 234614
rect 229756 233206 229876 233234
rect 229940 233206 230060 233234
rect 229848 231854 229876 233206
rect 229848 231826 229968 231854
rect 229742 227352 229798 227361
rect 229742 227287 229798 227296
rect 229650 217424 229706 217433
rect 229650 217359 229706 217368
rect 229560 161288 229612 161294
rect 229560 161230 229612 161236
rect 229468 140616 229520 140622
rect 229468 140558 229520 140564
rect 229756 138825 229784 227287
rect 229940 225690 229968 231826
rect 230032 229094 230060 233206
rect 230032 229066 230152 229094
rect 229928 225684 229980 225690
rect 229928 225626 229980 225632
rect 229836 224052 229888 224058
rect 229836 223994 229888 224000
rect 229848 151026 229876 223994
rect 230020 222964 230072 222970
rect 230020 222906 230072 222912
rect 229928 219428 229980 219434
rect 229928 219370 229980 219376
rect 229940 219094 229968 219370
rect 229928 219088 229980 219094
rect 229928 219030 229980 219036
rect 229940 158982 229968 219030
rect 230032 188329 230060 222906
rect 230018 188320 230074 188329
rect 230018 188255 230074 188264
rect 230124 160750 230152 229066
rect 230216 220833 230244 234586
rect 230584 224954 230612 239720
rect 230722 239714 230750 240108
rect 230814 239902 230842 240108
rect 230906 239902 230934 240108
rect 230998 239902 231026 240108
rect 231090 239902 231118 240108
rect 230802 239896 230854 239902
rect 230800 239864 230802 239873
rect 230894 239896 230946 239902
rect 230854 239864 230856 239873
rect 230894 239838 230946 239844
rect 230986 239896 231038 239902
rect 230986 239838 231038 239844
rect 231078 239896 231130 239902
rect 231182 239873 231210 240108
rect 231274 239970 231302 240108
rect 231262 239964 231314 239970
rect 231262 239906 231314 239912
rect 231078 239838 231130 239844
rect 231168 239864 231224 239873
rect 230800 239799 230856 239808
rect 231366 239850 231394 240108
rect 231458 239970 231486 240108
rect 231550 239970 231578 240108
rect 231446 239964 231498 239970
rect 231446 239906 231498 239912
rect 231538 239964 231590 239970
rect 231538 239906 231590 239912
rect 231366 239822 231440 239850
rect 231168 239799 231224 239808
rect 231412 239816 231440 239822
rect 231642 239816 231670 240108
rect 231734 239970 231762 240108
rect 231722 239964 231774 239970
rect 231722 239906 231774 239912
rect 231826 239816 231854 240108
rect 231918 239873 231946 240108
rect 232010 239970 232038 240108
rect 232102 239970 232130 240108
rect 231998 239964 232050 239970
rect 231998 239906 232050 239912
rect 232090 239964 232142 239970
rect 232090 239906 232142 239912
rect 231412 239788 231532 239816
rect 230848 239760 230900 239766
rect 230722 239686 230796 239714
rect 231216 239760 231268 239766
rect 231122 239728 231178 239737
rect 230900 239708 230980 239714
rect 230848 239702 230980 239708
rect 230860 239686 230980 239702
rect 230664 239556 230716 239562
rect 230664 239498 230716 239504
rect 230676 238134 230704 239498
rect 230664 238128 230716 238134
rect 230664 238070 230716 238076
rect 230768 237386 230796 239686
rect 230848 239624 230900 239630
rect 230848 239566 230900 239572
rect 230860 238474 230888 239566
rect 230848 238468 230900 238474
rect 230848 238410 230900 238416
rect 230756 237380 230808 237386
rect 230756 237322 230808 237328
rect 230756 236564 230808 236570
rect 230756 236506 230808 236512
rect 230492 224926 230612 224954
rect 230202 220824 230258 220833
rect 230202 220759 230258 220768
rect 230492 220425 230520 224926
rect 230768 221610 230796 236506
rect 230860 231169 230888 238410
rect 230952 236570 230980 239686
rect 231504 239737 231532 239788
rect 231596 239788 231670 239816
rect 231780 239788 231854 239816
rect 231904 239864 231960 239873
rect 232194 239850 232222 240108
rect 232286 239970 232314 240108
rect 232378 239970 232406 240108
rect 232274 239964 232326 239970
rect 232274 239906 232326 239912
rect 232366 239964 232418 239970
rect 232366 239906 232418 239912
rect 231904 239799 231960 239808
rect 232044 239828 232096 239834
rect 231216 239702 231268 239708
rect 231490 239728 231546 239737
rect 231122 239663 231178 239672
rect 231136 239630 231164 239663
rect 231124 239624 231176 239630
rect 231044 239584 231124 239612
rect 230940 236564 230992 236570
rect 230940 236506 230992 236512
rect 230846 231160 230902 231169
rect 230846 231095 230902 231104
rect 230756 221604 230808 221610
rect 230756 221546 230808 221552
rect 230478 220416 230534 220425
rect 230478 220351 230534 220360
rect 230492 217705 230520 220351
rect 230572 219360 230624 219366
rect 230572 219302 230624 219308
rect 230478 217696 230534 217705
rect 230478 217631 230534 217640
rect 230584 217297 230612 219302
rect 230570 217288 230626 217297
rect 230570 217223 230626 217232
rect 231044 217161 231072 239584
rect 231124 239566 231176 239572
rect 231124 238944 231176 238950
rect 231124 238886 231176 238892
rect 231136 238785 231164 238886
rect 231122 238776 231178 238785
rect 231122 238711 231178 238720
rect 231122 238232 231178 238241
rect 231122 238167 231178 238176
rect 231136 231577 231164 238167
rect 231228 236638 231256 239702
rect 231308 239692 231360 239698
rect 231490 239663 231546 239672
rect 231308 239634 231360 239640
rect 231320 238134 231348 239634
rect 231492 239624 231544 239630
rect 231492 239566 231544 239572
rect 231504 238660 231532 239566
rect 231596 238950 231624 239788
rect 231780 239714 231808 239788
rect 232194 239822 232268 239850
rect 232044 239770 232096 239776
rect 231688 239686 231808 239714
rect 231584 238944 231636 238950
rect 231584 238886 231636 238892
rect 231412 238632 231532 238660
rect 231412 238218 231440 238632
rect 231412 238202 231624 238218
rect 231412 238196 231636 238202
rect 231412 238190 231584 238196
rect 231308 238128 231360 238134
rect 231308 238070 231360 238076
rect 231216 236632 231268 236638
rect 231216 236574 231268 236580
rect 231412 231854 231440 238190
rect 231584 238138 231636 238144
rect 231492 238128 231544 238134
rect 231492 238070 231544 238076
rect 231320 231826 231440 231854
rect 231504 231854 231532 238070
rect 231688 237590 231716 239686
rect 231768 239624 231820 239630
rect 231766 239592 231768 239601
rect 231820 239592 231822 239601
rect 231766 239527 231822 239536
rect 231950 239592 232006 239601
rect 231950 239527 232006 239536
rect 231780 238270 231808 239527
rect 231860 239488 231912 239494
rect 231860 239430 231912 239436
rect 231768 238264 231820 238270
rect 231768 238206 231820 238212
rect 231676 237584 231728 237590
rect 231676 237526 231728 237532
rect 231504 231826 231624 231854
rect 231122 231568 231178 231577
rect 231122 231503 231178 231512
rect 231320 229094 231348 231826
rect 231320 229066 231440 229094
rect 231124 227588 231176 227594
rect 231124 227530 231176 227536
rect 231030 217152 231086 217161
rect 231030 217087 231086 217096
rect 230112 160744 230164 160750
rect 230112 160686 230164 160692
rect 229928 158976 229980 158982
rect 229928 158918 229980 158924
rect 229836 151020 229888 151026
rect 229836 150962 229888 150968
rect 231136 143138 231164 227530
rect 231306 221368 231362 221377
rect 231306 221303 231362 221312
rect 231214 218784 231270 218793
rect 231214 218719 231270 218728
rect 231124 143132 231176 143138
rect 231124 143074 231176 143080
rect 231228 138961 231256 218719
rect 231320 145761 231348 221303
rect 231412 173505 231440 229066
rect 231492 221604 231544 221610
rect 231492 221546 231544 221552
rect 231398 173496 231454 173505
rect 231398 173431 231454 173440
rect 231504 158778 231532 221546
rect 231596 184249 231624 231826
rect 231688 215937 231716 237526
rect 231768 237380 231820 237386
rect 231768 237322 231820 237328
rect 231780 219366 231808 237322
rect 231872 232626 231900 239430
rect 231860 232620 231912 232626
rect 231860 232562 231912 232568
rect 231768 219360 231820 219366
rect 231768 219302 231820 219308
rect 231674 215928 231730 215937
rect 231674 215863 231730 215872
rect 231964 213625 231992 239527
rect 232056 238785 232084 239770
rect 232136 239760 232188 239766
rect 232136 239702 232188 239708
rect 232042 238776 232098 238785
rect 232042 238711 232098 238720
rect 232056 231854 232084 238711
rect 232148 238610 232176 239702
rect 232136 238604 232188 238610
rect 232136 238546 232188 238552
rect 232148 237658 232176 238546
rect 232136 237652 232188 237658
rect 232136 237594 232188 237600
rect 232240 237425 232268 239822
rect 232320 239828 232372 239834
rect 232470 239816 232498 240108
rect 232320 239770 232372 239776
rect 232424 239788 232498 239816
rect 232332 239737 232360 239770
rect 232318 239728 232374 239737
rect 232318 239663 232374 239672
rect 232424 238814 232452 239788
rect 232562 239714 232590 240108
rect 232654 239816 232682 240108
rect 232746 239970 232774 240108
rect 232838 239970 232866 240108
rect 232734 239964 232786 239970
rect 232734 239906 232786 239912
rect 232826 239964 232878 239970
rect 232826 239906 232878 239912
rect 232930 239850 232958 240108
rect 232884 239822 232958 239850
rect 233022 239850 233050 240108
rect 233114 239970 233142 240108
rect 233102 239964 233154 239970
rect 233102 239906 233154 239912
rect 233206 239873 233234 240108
rect 233192 239864 233248 239873
rect 233022 239822 233096 239850
rect 232654 239788 232728 239816
rect 232516 239686 232590 239714
rect 232320 238808 232372 238814
rect 232320 238750 232372 238756
rect 232412 238808 232464 238814
rect 232412 238750 232464 238756
rect 232332 238610 232360 238750
rect 232320 238604 232372 238610
rect 232320 238546 232372 238552
rect 232226 237416 232282 237425
rect 232226 237351 232282 237360
rect 232056 231826 232176 231854
rect 232044 231464 232096 231470
rect 232044 231406 232096 231412
rect 232056 225758 232084 231406
rect 232148 229094 232176 231826
rect 232424 231470 232452 238750
rect 232412 231464 232464 231470
rect 232412 231406 232464 231412
rect 232148 229066 232452 229094
rect 232044 225752 232096 225758
rect 232044 225694 232096 225700
rect 232424 215121 232452 229066
rect 232516 224738 232544 239686
rect 232596 239624 232648 239630
rect 232596 239566 232648 239572
rect 232608 238406 232636 239566
rect 232596 238400 232648 238406
rect 232596 238342 232648 238348
rect 232700 234614 232728 239788
rect 232884 239601 232912 239822
rect 233068 239714 233096 239822
rect 233192 239799 233248 239808
rect 233298 239816 233326 240108
rect 233390 239970 233418 240108
rect 233482 239970 233510 240108
rect 233378 239964 233430 239970
rect 233378 239906 233430 239912
rect 233470 239964 233522 239970
rect 233470 239906 233522 239912
rect 233422 239864 233478 239873
rect 233206 239748 233234 239799
rect 233298 239788 233372 239816
rect 233422 239799 233424 239808
rect 232976 239686 233096 239714
rect 233160 239720 233234 239748
rect 232870 239592 232926 239601
rect 232870 239527 232926 239536
rect 232780 239352 232832 239358
rect 232780 239294 232832 239300
rect 232792 238649 232820 239294
rect 232778 238640 232834 238649
rect 232778 238575 232834 238584
rect 232870 235784 232926 235793
rect 232870 235719 232926 235728
rect 232884 235550 232912 235719
rect 232872 235544 232924 235550
rect 232872 235486 232924 235492
rect 232608 234586 232728 234614
rect 232608 229094 232636 234586
rect 232976 234002 233004 239686
rect 233056 239624 233108 239630
rect 233056 239566 233108 239572
rect 233068 235618 233096 239566
rect 233056 235612 233108 235618
rect 233056 235554 233108 235560
rect 233054 235376 233110 235385
rect 233054 235311 233110 235320
rect 232792 233974 233004 234002
rect 232792 230450 232820 233974
rect 232872 233776 232924 233782
rect 232872 233718 232924 233724
rect 232780 230444 232832 230450
rect 232780 230386 232832 230392
rect 232608 229066 232820 229094
rect 232504 224732 232556 224738
rect 232504 224674 232556 224680
rect 232410 215112 232466 215121
rect 232410 215047 232466 215056
rect 231950 213616 232006 213625
rect 231950 213551 232006 213560
rect 231582 184240 231638 184249
rect 231582 184175 231638 184184
rect 232516 159050 232544 224674
rect 232688 224664 232740 224670
rect 232688 224606 232740 224612
rect 232596 221944 232648 221950
rect 232596 221886 232648 221892
rect 232504 159044 232556 159050
rect 232504 158986 232556 158992
rect 231492 158772 231544 158778
rect 231492 158714 231544 158720
rect 232504 149728 232556 149734
rect 232504 149670 232556 149676
rect 231306 145752 231362 145761
rect 231306 145687 231362 145696
rect 231214 138952 231270 138961
rect 231214 138887 231270 138896
rect 229742 138816 229798 138825
rect 229742 138751 229798 138760
rect 230478 124808 230534 124817
rect 230478 124743 230534 124752
rect 230492 16574 230520 124743
rect 229112 16546 229416 16574
rect 230492 16546 231072 16574
rect 228364 3936 228416 3942
rect 228364 3878 228416 3884
rect 228732 3052 228784 3058
rect 228732 2994 228784 3000
rect 228744 480 228772 2994
rect 223918 354 224030 480
rect 223592 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229388 354 229416 16546
rect 231044 480 231072 16546
rect 232516 4146 232544 149670
rect 232608 138689 232636 221886
rect 232700 149841 232728 224606
rect 232792 222970 232820 229066
rect 232780 222964 232832 222970
rect 232780 222906 232832 222912
rect 232792 213353 232820 222906
rect 232778 213344 232834 213353
rect 232778 213279 232834 213288
rect 232884 159118 232912 233718
rect 233068 229094 233096 235311
rect 233160 233782 233188 239720
rect 233240 239624 233292 239630
rect 233344 239601 233372 239788
rect 233476 239799 233478 239808
rect 233424 239770 233476 239776
rect 233574 239748 233602 240108
rect 233666 239970 233694 240108
rect 233758 239970 233786 240108
rect 233654 239964 233706 239970
rect 233654 239906 233706 239912
rect 233746 239964 233798 239970
rect 233746 239906 233798 239912
rect 233700 239828 233752 239834
rect 233700 239770 233752 239776
rect 233422 239728 233478 239737
rect 233422 239663 233478 239672
rect 233528 239720 233602 239748
rect 233712 239737 233740 239770
rect 233698 239728 233754 239737
rect 233240 239566 233292 239572
rect 233330 239592 233386 239601
rect 233252 239465 233280 239566
rect 233436 239562 233464 239663
rect 233330 239527 233386 239536
rect 233424 239556 233476 239562
rect 233424 239498 233476 239504
rect 233238 239456 233294 239465
rect 233238 239391 233294 239400
rect 233424 239420 233476 239426
rect 233252 239034 233280 239391
rect 233424 239362 233476 239368
rect 233436 239222 233464 239362
rect 233424 239216 233476 239222
rect 233424 239158 233476 239164
rect 233252 239006 233372 239034
rect 233238 238776 233294 238785
rect 233238 238711 233294 238720
rect 233148 233776 233200 233782
rect 233148 233718 233200 233724
rect 233252 229945 233280 238711
rect 233238 229936 233294 229945
rect 233238 229871 233294 229880
rect 233068 229066 233188 229094
rect 232872 159112 232924 159118
rect 232872 159054 232924 159060
rect 233160 154222 233188 229066
rect 233148 154216 233200 154222
rect 233148 154158 233200 154164
rect 233240 151088 233292 151094
rect 233240 151030 233292 151036
rect 233252 150482 233280 151030
rect 233240 150476 233292 150482
rect 233240 150418 233292 150424
rect 232686 149832 232742 149841
rect 232686 149767 232742 149776
rect 232594 138680 232650 138689
rect 232594 138615 232650 138624
rect 233252 16574 233280 150418
rect 233344 147286 233372 239006
rect 233528 238678 233556 239720
rect 233850 239714 233878 240108
rect 233942 239902 233970 240108
rect 234034 239970 234062 240108
rect 234022 239964 234074 239970
rect 234022 239906 234074 239912
rect 233930 239896 233982 239902
rect 233930 239838 233982 239844
rect 234126 239714 234154 240108
rect 234218 239970 234246 240108
rect 234206 239964 234258 239970
rect 234206 239906 234258 239912
rect 234310 239873 234338 240108
rect 234402 239902 234430 240108
rect 234390 239896 234442 239902
rect 234296 239864 234352 239873
rect 234390 239838 234442 239844
rect 234494 239850 234522 240108
rect 234586 239970 234614 240108
rect 234574 239964 234626 239970
rect 234574 239906 234626 239912
rect 234494 239822 234568 239850
rect 234296 239799 234352 239808
rect 233698 239663 233754 239672
rect 233804 239686 233878 239714
rect 233976 239692 234028 239698
rect 233804 239544 233832 239686
rect 233976 239634 234028 239640
rect 234080 239686 234154 239714
rect 234252 239760 234304 239766
rect 234252 239702 234304 239708
rect 234434 239728 234490 239737
rect 233988 239544 234016 239634
rect 233712 239516 233832 239544
rect 233896 239516 234016 239544
rect 233516 238672 233568 238678
rect 233516 238614 233568 238620
rect 233606 238640 233662 238649
rect 233606 238575 233662 238584
rect 233424 235952 233476 235958
rect 233424 235894 233476 235900
rect 233436 231810 233464 235894
rect 233424 231804 233476 231810
rect 233424 231746 233476 231752
rect 233516 230444 233568 230450
rect 233516 230386 233568 230392
rect 233528 229838 233556 230386
rect 233516 229832 233568 229838
rect 233516 229774 233568 229780
rect 233528 157214 233556 229774
rect 233620 220289 233648 238575
rect 233712 235958 233740 239516
rect 233790 239456 233846 239465
rect 233790 239391 233792 239400
rect 233844 239391 233846 239400
rect 233792 239362 233844 239368
rect 233792 238672 233844 238678
rect 233792 238614 233844 238620
rect 233700 235952 233752 235958
rect 233700 235894 233752 235900
rect 233700 232076 233752 232082
rect 233700 232018 233752 232024
rect 233712 224330 233740 232018
rect 233804 231441 233832 238614
rect 233896 236065 233924 239516
rect 233974 239456 234030 239465
rect 233974 239391 234030 239400
rect 233882 236056 233938 236065
rect 233882 235991 233938 236000
rect 233884 235952 233936 235958
rect 233884 235894 233936 235900
rect 233790 231432 233846 231441
rect 233790 231367 233846 231376
rect 233700 224324 233752 224330
rect 233700 224266 233752 224272
rect 233712 223650 233740 224266
rect 233700 223644 233752 223650
rect 233700 223586 233752 223592
rect 233606 220280 233662 220289
rect 233606 220215 233662 220224
rect 233516 157208 233568 157214
rect 233516 157150 233568 157156
rect 233332 147280 233384 147286
rect 233332 147222 233384 147228
rect 233896 141506 233924 235894
rect 233988 232937 234016 239391
rect 234080 236065 234108 239686
rect 234160 239624 234212 239630
rect 234160 239566 234212 239572
rect 234172 238649 234200 239566
rect 234158 238640 234214 238649
rect 234158 238575 234214 238584
rect 234160 237244 234212 237250
rect 234160 237186 234212 237192
rect 234066 236056 234122 236065
rect 234066 235991 234122 236000
rect 233974 232928 234030 232937
rect 233974 232863 234030 232872
rect 234068 231804 234120 231810
rect 234068 231746 234120 231752
rect 233976 230104 234028 230110
rect 233976 230046 234028 230052
rect 233988 150482 234016 230046
rect 234080 152386 234108 231746
rect 234172 227458 234200 237186
rect 234264 232082 234292 239702
rect 234344 239692 234396 239698
rect 234434 239663 234490 239672
rect 234344 239634 234396 239640
rect 234356 237250 234384 239634
rect 234448 239630 234476 239663
rect 234436 239624 234488 239630
rect 234436 239566 234488 239572
rect 234448 238678 234476 239566
rect 234436 238672 234488 238678
rect 234436 238614 234488 238620
rect 234540 238241 234568 239822
rect 234678 239816 234706 240108
rect 234770 239970 234798 240108
rect 234758 239964 234810 239970
rect 234758 239906 234810 239912
rect 234862 239873 234890 240108
rect 234848 239864 234904 239873
rect 234678 239788 234752 239816
rect 234954 239850 234982 240108
rect 235046 239970 235074 240108
rect 235034 239964 235086 239970
rect 235034 239906 235086 239912
rect 234954 239822 235028 239850
rect 234848 239799 234904 239808
rect 234620 238672 234672 238678
rect 234620 238614 234672 238620
rect 234526 238232 234582 238241
rect 234526 238167 234582 238176
rect 234434 238096 234490 238105
rect 234434 238031 234490 238040
rect 234448 237998 234476 238031
rect 234436 237992 234488 237998
rect 234436 237934 234488 237940
rect 234632 237930 234660 238614
rect 234620 237924 234672 237930
rect 234620 237866 234672 237872
rect 234344 237244 234396 237250
rect 234344 237186 234396 237192
rect 234724 237114 234752 239788
rect 234862 239748 234890 239799
rect 234816 239720 234890 239748
rect 234712 237108 234764 237114
rect 234712 237050 234764 237056
rect 234620 235544 234672 235550
rect 234620 235486 234672 235492
rect 234252 232076 234304 232082
rect 234252 232018 234304 232024
rect 234160 227452 234212 227458
rect 234160 227394 234212 227400
rect 234172 157078 234200 227394
rect 234160 157072 234212 157078
rect 234160 157014 234212 157020
rect 234068 152380 234120 152386
rect 234068 152322 234120 152328
rect 233976 150476 234028 150482
rect 233976 150418 234028 150424
rect 234632 141914 234660 235486
rect 234816 228478 234844 239720
rect 234896 239624 234948 239630
rect 234896 239566 234948 239572
rect 234908 239465 234936 239566
rect 234894 239456 234950 239465
rect 234894 239391 234950 239400
rect 234896 238264 234948 238270
rect 234896 238206 234948 238212
rect 234908 229770 234936 238206
rect 235000 236337 235028 239822
rect 235138 239816 235166 240108
rect 235230 239970 235258 240108
rect 235218 239964 235270 239970
rect 235218 239906 235270 239912
rect 235322 239850 235350 240108
rect 235414 239970 235442 240108
rect 235402 239964 235454 239970
rect 235402 239906 235454 239912
rect 235322 239822 235396 239850
rect 235092 239788 235166 239816
rect 235092 239737 235120 239788
rect 235264 239760 235316 239766
rect 235078 239728 235134 239737
rect 235264 239702 235316 239708
rect 235078 239663 235134 239672
rect 234986 236328 235042 236337
rect 234986 236263 235042 236272
rect 234896 229764 234948 229770
rect 234896 229706 234948 229712
rect 234804 228472 234856 228478
rect 234804 228414 234856 228420
rect 235092 226334 235120 239663
rect 235172 239624 235224 239630
rect 235172 239566 235224 239572
rect 235184 236745 235212 239566
rect 235276 238610 235304 239702
rect 235264 238604 235316 238610
rect 235264 238546 235316 238552
rect 235170 236736 235226 236745
rect 235170 236671 235226 236680
rect 235276 235006 235304 238546
rect 235368 237374 235396 239822
rect 235506 239816 235534 240108
rect 235598 239970 235626 240108
rect 235690 239970 235718 240108
rect 235782 239970 235810 240108
rect 235586 239964 235638 239970
rect 235586 239906 235638 239912
rect 235678 239964 235730 239970
rect 235678 239906 235730 239912
rect 235770 239964 235822 239970
rect 235770 239906 235822 239912
rect 235874 239816 235902 240108
rect 235966 239970 235994 240108
rect 235954 239964 236006 239970
rect 235954 239906 236006 239912
rect 236058 239902 236086 240108
rect 236046 239896 236098 239902
rect 236046 239838 236098 239844
rect 235506 239788 235672 239816
rect 235538 239728 235594 239737
rect 235448 239692 235500 239698
rect 235538 239663 235594 239672
rect 235448 239634 235500 239640
rect 235460 238785 235488 239634
rect 235552 239562 235580 239663
rect 235540 239556 235592 239562
rect 235540 239498 235592 239504
rect 235540 239420 235592 239426
rect 235540 239362 235592 239368
rect 235552 238950 235580 239362
rect 235540 238944 235592 238950
rect 235540 238886 235592 238892
rect 235446 238776 235502 238785
rect 235446 238711 235502 238720
rect 235540 238740 235592 238746
rect 235460 237998 235488 238711
rect 235540 238682 235592 238688
rect 235552 238610 235580 238682
rect 235540 238604 235592 238610
rect 235540 238546 235592 238552
rect 235448 237992 235500 237998
rect 235448 237934 235500 237940
rect 235368 237346 235580 237374
rect 235356 237312 235408 237318
rect 235356 237254 235408 237260
rect 235264 235000 235316 235006
rect 235264 234942 235316 234948
rect 235264 234252 235316 234258
rect 235264 234194 235316 234200
rect 235172 233980 235224 233986
rect 235172 233922 235224 233928
rect 235184 228342 235212 233922
rect 235172 228336 235224 228342
rect 235172 228278 235224 228284
rect 235184 227798 235212 228278
rect 235172 227792 235224 227798
rect 235172 227734 235224 227740
rect 234816 226306 235120 226334
rect 234816 213217 234844 226306
rect 234802 213208 234858 213217
rect 234802 213143 234858 213152
rect 235276 155718 235304 234194
rect 235368 234190 235396 237254
rect 235356 234184 235408 234190
rect 235356 234126 235408 234132
rect 235368 233730 235396 234126
rect 235368 233702 235488 233730
rect 235354 229800 235410 229809
rect 235354 229735 235410 229744
rect 235264 155712 235316 155718
rect 235264 155654 235316 155660
rect 235368 152862 235396 229735
rect 235460 157010 235488 233702
rect 235552 228818 235580 237346
rect 235644 234258 235672 239788
rect 235828 239788 235902 239816
rect 235724 239420 235776 239426
rect 235724 239362 235776 239368
rect 235736 237318 235764 239362
rect 235724 237312 235776 237318
rect 235724 237254 235776 237260
rect 235632 234252 235684 234258
rect 235632 234194 235684 234200
rect 235828 233986 235856 239788
rect 236000 239760 236052 239766
rect 235920 239720 236000 239748
rect 235920 239465 235948 239720
rect 236150 239748 236178 240108
rect 236104 239737 236178 239748
rect 236000 239702 236052 239708
rect 236090 239728 236178 239737
rect 236146 239720 236178 239728
rect 236090 239663 236146 239672
rect 236242 239680 236270 240108
rect 236334 239873 236362 240108
rect 236320 239864 236376 239873
rect 236320 239799 236376 239808
rect 236426 239748 236454 240108
rect 236518 239873 236546 240108
rect 236610 239970 236638 240108
rect 236598 239964 236650 239970
rect 236598 239906 236650 239912
rect 236702 239902 236730 240108
rect 236690 239896 236742 239902
rect 236504 239864 236560 239873
rect 236690 239838 236742 239844
rect 236504 239799 236560 239808
rect 236380 239720 236454 239748
rect 236794 239748 236822 240108
rect 236886 239970 236914 240108
rect 236874 239964 236926 239970
rect 236874 239906 236926 239912
rect 236978 239850 237006 240108
rect 237070 239970 237098 240108
rect 237058 239964 237110 239970
rect 237058 239906 237110 239912
rect 237162 239850 237190 240108
rect 236978 239834 237052 239850
rect 236978 239828 237064 239834
rect 236978 239822 237012 239828
rect 237012 239770 237064 239776
rect 237116 239822 237190 239850
rect 236920 239760 236972 239766
rect 236550 239728 236606 239737
rect 236242 239652 236316 239680
rect 236092 239624 236144 239630
rect 236092 239566 236144 239572
rect 236000 239488 236052 239494
rect 235906 239456 235962 239465
rect 236000 239430 236052 239436
rect 235906 239391 235962 239400
rect 236012 238746 236040 239430
rect 236000 238740 236052 238746
rect 236000 238682 236052 238688
rect 236104 238082 236132 239566
rect 236182 239456 236238 239465
rect 236182 239391 236238 239400
rect 236196 239154 236224 239391
rect 236184 239148 236236 239154
rect 236184 239090 236236 239096
rect 236012 238054 236132 238082
rect 236012 237522 236040 238054
rect 236092 237992 236144 237998
rect 236092 237934 236144 237940
rect 236000 237516 236052 237522
rect 236000 237458 236052 237464
rect 236012 235686 236040 237458
rect 236000 235680 236052 235686
rect 236000 235622 236052 235628
rect 235816 233980 235868 233986
rect 235816 233922 235868 233928
rect 235540 228812 235592 228818
rect 235540 228754 235592 228760
rect 235448 157004 235500 157010
rect 235448 156946 235500 156952
rect 235552 153105 235580 228754
rect 235632 227792 235684 227798
rect 235632 227734 235684 227740
rect 235644 154358 235672 227734
rect 235632 154352 235684 154358
rect 235632 154294 235684 154300
rect 235538 153096 235594 153105
rect 235538 153031 235594 153040
rect 235356 152856 235408 152862
rect 235356 152798 235408 152804
rect 235368 142154 235396 152798
rect 236000 151224 236052 151230
rect 236000 151166 236052 151172
rect 236012 150550 236040 151166
rect 236000 150544 236052 150550
rect 236000 150486 236052 150492
rect 235276 142126 235396 142154
rect 234620 141908 234672 141914
rect 234620 141850 234672 141856
rect 233884 141500 233936 141506
rect 233884 141442 233936 141448
rect 234710 98832 234766 98841
rect 234710 98767 234766 98776
rect 233252 16546 233464 16574
rect 232504 4140 232556 4146
rect 232504 4082 232556 4088
rect 232228 3868 232280 3874
rect 232228 3810 232280 3816
rect 232240 480 232268 3810
rect 233436 480 233464 16546
rect 234724 6914 234752 98767
rect 234632 6886 234752 6914
rect 234632 480 234660 6886
rect 235276 4078 235304 142126
rect 236012 16574 236040 150486
rect 236104 145858 236132 237934
rect 236288 237862 236316 239652
rect 236380 238678 236408 239720
rect 236794 239720 236920 239748
rect 236920 239702 236972 239708
rect 236550 239663 236606 239672
rect 236460 239556 236512 239562
rect 236460 239498 236512 239504
rect 236472 238785 236500 239498
rect 236458 238776 236514 238785
rect 236458 238711 236514 238720
rect 236368 238672 236420 238678
rect 236368 238614 236420 238620
rect 236458 238232 236514 238241
rect 236458 238167 236514 238176
rect 236276 237856 236328 237862
rect 236276 237798 236328 237804
rect 236366 237552 236422 237561
rect 236366 237487 236422 237496
rect 236184 237040 236236 237046
rect 236182 237008 236184 237017
rect 236236 237008 236238 237017
rect 236182 236943 236238 236952
rect 236182 236192 236238 236201
rect 236182 236127 236238 236136
rect 236196 213081 236224 236127
rect 236380 213761 236408 237487
rect 236472 228274 236500 238167
rect 236564 235482 236592 239663
rect 236828 239624 236880 239630
rect 236828 239566 236880 239572
rect 236920 239624 236972 239630
rect 236920 239566 236972 239572
rect 236734 238776 236790 238785
rect 236734 238711 236790 238720
rect 236644 238400 236696 238406
rect 236644 238342 236696 238348
rect 236656 237998 236684 238342
rect 236644 237992 236696 237998
rect 236644 237934 236696 237940
rect 236552 235476 236604 235482
rect 236552 235418 236604 235424
rect 236642 235240 236698 235249
rect 236642 235175 236698 235184
rect 236552 228472 236604 228478
rect 236552 228414 236604 228420
rect 236460 228268 236512 228274
rect 236460 228210 236512 228216
rect 236472 225622 236500 228210
rect 236564 227050 236592 228414
rect 236552 227044 236604 227050
rect 236552 226986 236604 226992
rect 236460 225616 236512 225622
rect 236460 225558 236512 225564
rect 236366 213752 236422 213761
rect 236366 213687 236422 213696
rect 236182 213072 236238 213081
rect 236182 213007 236238 213016
rect 236092 145852 236144 145858
rect 236092 145794 236144 145800
rect 236656 141545 236684 235175
rect 236748 233102 236776 238711
rect 236736 233096 236788 233102
rect 236736 233038 236788 233044
rect 236736 232892 236788 232898
rect 236840 232880 236868 239566
rect 236932 239154 236960 239566
rect 237012 239556 237064 239562
rect 237012 239498 237064 239504
rect 237024 239465 237052 239498
rect 237010 239456 237066 239465
rect 237010 239391 237066 239400
rect 237012 239352 237064 239358
rect 237012 239294 237064 239300
rect 236920 239148 236972 239154
rect 236920 239090 236972 239096
rect 236918 238232 236974 238241
rect 236918 238167 236974 238176
rect 236932 237794 236960 238167
rect 237024 237930 237052 239294
rect 237012 237924 237064 237930
rect 237012 237866 237064 237872
rect 236920 237788 236972 237794
rect 236920 237730 236972 237736
rect 237012 233096 237064 233102
rect 237012 233038 237064 233044
rect 236788 232852 236868 232880
rect 236736 232834 236788 232840
rect 236748 221474 236776 232834
rect 236920 232280 236972 232286
rect 236920 232222 236972 232228
rect 236932 227118 236960 232222
rect 237024 229094 237052 233038
rect 237116 232286 237144 239822
rect 237254 239748 237282 240108
rect 237346 239907 237374 240108
rect 237438 239970 237466 240108
rect 237530 239970 237558 240108
rect 237426 239964 237478 239970
rect 237332 239898 237388 239907
rect 237426 239906 237478 239912
rect 237518 239964 237570 239970
rect 237518 239906 237570 239912
rect 237622 239902 237650 240108
rect 237332 239833 237388 239842
rect 237610 239896 237662 239902
rect 237610 239838 237662 239844
rect 237714 239850 237742 240108
rect 237806 239970 237834 240108
rect 237794 239964 237846 239970
rect 237794 239906 237846 239912
rect 237898 239902 237926 240108
rect 237990 239902 238018 240108
rect 237886 239896 237938 239902
rect 237714 239822 237788 239850
rect 237886 239838 237938 239844
rect 237978 239896 238030 239902
rect 237978 239838 238030 239844
rect 237254 239720 237328 239748
rect 237300 239544 237328 239720
rect 237654 239728 237710 239737
rect 237564 239692 237616 239698
rect 237654 239663 237710 239672
rect 237564 239634 237616 239640
rect 237472 239624 237524 239630
rect 237472 239566 237524 239572
rect 237208 239516 237328 239544
rect 237208 237833 237236 239516
rect 237288 239420 237340 239426
rect 237288 239362 237340 239368
rect 237194 237824 237250 237833
rect 237194 237759 237250 237768
rect 237300 237153 237328 239362
rect 237380 239352 237432 239358
rect 237380 239294 237432 239300
rect 237286 237144 237342 237153
rect 237286 237079 237342 237088
rect 237288 232620 237340 232626
rect 237288 232562 237340 232568
rect 237104 232280 237156 232286
rect 237104 232222 237156 232228
rect 237024 229066 237144 229094
rect 237300 229090 237328 232562
rect 236920 227112 236972 227118
rect 236920 227054 236972 227060
rect 237012 226908 237064 226914
rect 237012 226850 237064 226856
rect 236826 226808 236882 226817
rect 236826 226743 236882 226752
rect 236736 221468 236788 221474
rect 236736 221410 236788 221416
rect 236734 218920 236790 218929
rect 236734 218855 236790 218864
rect 236748 143041 236776 218855
rect 236840 153921 236868 226743
rect 236918 224768 236974 224777
rect 236918 224703 236974 224712
rect 236826 153912 236882 153921
rect 236826 153847 236882 153856
rect 236932 150550 236960 224703
rect 237024 155446 237052 226850
rect 237116 222902 237144 229066
rect 237288 229084 237340 229090
rect 237288 229026 237340 229032
rect 237300 228886 237328 229026
rect 237288 228880 237340 228886
rect 237288 228822 237340 228828
rect 237392 227186 237420 239294
rect 237484 237046 237512 239566
rect 237472 237040 237524 237046
rect 237472 236982 237524 236988
rect 237472 236632 237524 236638
rect 237472 236574 237524 236580
rect 237484 235958 237512 236574
rect 237472 235952 237524 235958
rect 237472 235894 237524 235900
rect 237470 235784 237526 235793
rect 237470 235719 237526 235728
rect 237484 228954 237512 235719
rect 237576 234394 237604 239634
rect 237668 239562 237696 239663
rect 237656 239556 237708 239562
rect 237656 239498 237708 239504
rect 237668 238270 237696 239498
rect 237656 238264 237708 238270
rect 237656 238206 237708 238212
rect 237760 238066 237788 239822
rect 238082 239816 238110 240108
rect 238174 239970 238202 240108
rect 238266 239970 238294 240108
rect 238162 239964 238214 239970
rect 238162 239906 238214 239912
rect 238254 239964 238306 239970
rect 238254 239906 238306 239912
rect 238358 239816 238386 240108
rect 238450 239970 238478 240108
rect 238438 239964 238490 239970
rect 238438 239906 238490 239912
rect 238542 239907 238570 240108
rect 238634 239970 238662 240108
rect 238622 239964 238674 239970
rect 238528 239898 238584 239907
rect 238622 239906 238674 239912
rect 238726 239902 238754 240108
rect 238528 239833 238584 239842
rect 238714 239896 238766 239902
rect 238714 239838 238766 239844
rect 238082 239788 238156 239816
rect 238358 239788 238432 239816
rect 237932 239692 237984 239698
rect 237932 239634 237984 239640
rect 238024 239692 238076 239698
rect 238024 239634 238076 239640
rect 237840 239624 237892 239630
rect 237840 239566 237892 239572
rect 237852 239154 237880 239566
rect 237840 239148 237892 239154
rect 237840 239090 237892 239096
rect 237840 238740 237892 238746
rect 237840 238682 237892 238688
rect 237748 238060 237800 238066
rect 237748 238002 237800 238008
rect 237656 237924 237708 237930
rect 237656 237866 237708 237872
rect 237564 234388 237616 234394
rect 237564 234330 237616 234336
rect 237472 228948 237524 228954
rect 237472 228890 237524 228896
rect 237380 227180 237432 227186
rect 237380 227122 237432 227128
rect 237104 222896 237156 222902
rect 237104 222838 237156 222844
rect 237576 218754 237604 234330
rect 237668 228478 237696 237866
rect 237852 237368 237880 238682
rect 237760 237340 237880 237368
rect 237760 236638 237788 237340
rect 237944 237017 237972 239634
rect 238036 238746 238064 239634
rect 238128 239494 238156 239788
rect 238300 239692 238352 239698
rect 238220 239652 238300 239680
rect 238116 239488 238168 239494
rect 238116 239430 238168 239436
rect 238116 239148 238168 239154
rect 238116 239090 238168 239096
rect 238024 238740 238076 238746
rect 238024 238682 238076 238688
rect 238128 238116 238156 239090
rect 238220 238252 238248 239652
rect 238300 239634 238352 239640
rect 238298 239456 238354 239465
rect 238298 239391 238354 239400
rect 238312 239358 238340 239391
rect 238300 239352 238352 239358
rect 238300 239294 238352 239300
rect 238404 238320 238432 239788
rect 238484 239760 238536 239766
rect 238818 239748 238846 240108
rect 238910 239873 238938 240108
rect 238896 239864 238952 239873
rect 238896 239799 238952 239808
rect 239002 239748 239030 240108
rect 239094 239902 239122 240108
rect 239082 239896 239134 239902
rect 239082 239838 239134 239844
rect 239186 239850 239214 240108
rect 239278 239970 239306 240108
rect 239370 239970 239398 240108
rect 239462 239970 239490 240108
rect 239266 239964 239318 239970
rect 239266 239906 239318 239912
rect 239358 239964 239410 239970
rect 239358 239906 239410 239912
rect 239450 239964 239502 239970
rect 239450 239906 239502 239912
rect 239554 239873 239582 240108
rect 239540 239864 239596 239873
rect 239186 239834 239260 239850
rect 239186 239828 239272 239834
rect 239186 239822 239220 239828
rect 239540 239799 239596 239808
rect 239220 239770 239272 239776
rect 239312 239760 239364 239766
rect 238818 239720 238892 239748
rect 239002 239720 239076 239748
rect 238484 239702 238536 239708
rect 238496 238882 238524 239702
rect 238668 239692 238720 239698
rect 238668 239634 238720 239640
rect 238576 239624 238628 239630
rect 238576 239566 238628 239572
rect 238588 239154 238616 239566
rect 238680 239465 238708 239634
rect 238666 239456 238722 239465
rect 238666 239391 238722 239400
rect 238760 239420 238812 239426
rect 238760 239362 238812 239368
rect 238668 239352 238720 239358
rect 238668 239294 238720 239300
rect 238576 239148 238628 239154
rect 238576 239090 238628 239096
rect 238484 238876 238536 238882
rect 238484 238818 238536 238824
rect 238404 238292 238524 238320
rect 238220 238224 238432 238252
rect 238128 238088 238340 238116
rect 238024 237924 238076 237930
rect 238024 237866 238076 237872
rect 237930 237008 237986 237017
rect 237930 236943 237986 236952
rect 237748 236632 237800 236638
rect 237748 236574 237800 236580
rect 238036 230738 238064 237866
rect 238114 236736 238170 236745
rect 238114 236671 238170 236680
rect 237944 230710 238064 230738
rect 237656 228472 237708 228478
rect 237656 228414 237708 228420
rect 237944 224058 237972 230710
rect 238128 229094 238156 236671
rect 238208 236428 238260 236434
rect 238208 236370 238260 236376
rect 238036 229066 238156 229094
rect 237932 224052 237984 224058
rect 237932 223994 237984 224000
rect 237564 218748 237616 218754
rect 237564 218690 237616 218696
rect 237012 155440 237064 155446
rect 237012 155382 237064 155388
rect 236920 150544 236972 150550
rect 236920 150486 236972 150492
rect 236734 143032 236790 143041
rect 236734 142967 236790 142976
rect 236642 141536 236698 141545
rect 236642 141471 236698 141480
rect 238036 136406 238064 229066
rect 238116 227656 238168 227662
rect 238116 227598 238168 227604
rect 238128 144265 238156 227598
rect 238220 154154 238248 236370
rect 238312 224670 238340 238088
rect 238404 237726 238432 238224
rect 238392 237720 238444 237726
rect 238392 237662 238444 237668
rect 238404 237017 238432 237662
rect 238390 237008 238446 237017
rect 238390 236943 238446 236952
rect 238496 229378 238524 238292
rect 238588 236774 238616 239090
rect 238576 236768 238628 236774
rect 238576 236710 238628 236716
rect 238680 235521 238708 239294
rect 238772 235657 238800 239362
rect 238864 238610 238892 239720
rect 238944 239488 238996 239494
rect 238942 239456 238944 239465
rect 238996 239456 238998 239465
rect 238942 239391 238998 239400
rect 239048 239358 239076 239720
rect 239646 239748 239674 240108
rect 239738 239816 239766 240108
rect 239830 239970 239858 240108
rect 239818 239964 239870 239970
rect 239818 239906 239870 239912
rect 239738 239788 239812 239816
rect 239364 239720 239444 239748
rect 239646 239720 239720 239748
rect 239312 239702 239364 239708
rect 239220 239692 239272 239698
rect 239220 239634 239272 239640
rect 239036 239352 239088 239358
rect 239036 239294 239088 239300
rect 239036 238808 239088 238814
rect 239232 238762 239260 239634
rect 239312 239488 239364 239494
rect 239310 239456 239312 239465
rect 239364 239456 239366 239465
rect 239310 239391 239366 239400
rect 239036 238750 239088 238756
rect 238852 238604 238904 238610
rect 238852 238546 238904 238552
rect 239048 238406 239076 238750
rect 239140 238734 239260 238762
rect 239036 238400 239088 238406
rect 239036 238342 239088 238348
rect 238850 238232 238906 238241
rect 238850 238167 238906 238176
rect 238758 235648 238814 235657
rect 238758 235583 238814 235592
rect 238666 235512 238722 235521
rect 238666 235447 238722 235456
rect 238404 229350 238524 229378
rect 238300 224664 238352 224670
rect 238300 224606 238352 224612
rect 238404 224602 238432 229350
rect 238576 227316 238628 227322
rect 238576 227258 238628 227264
rect 238484 227180 238536 227186
rect 238484 227122 238536 227128
rect 238392 224596 238444 224602
rect 238392 224538 238444 224544
rect 238298 221504 238354 221513
rect 238298 221439 238354 221448
rect 238208 154148 238260 154154
rect 238208 154090 238260 154096
rect 238114 144256 238170 144265
rect 238114 144191 238170 144200
rect 238312 144129 238340 221439
rect 238404 149938 238432 224538
rect 238496 154329 238524 227122
rect 238588 159497 238616 227258
rect 238864 213897 238892 238167
rect 238942 237552 238998 237561
rect 238942 237487 238998 237496
rect 238956 232626 238984 237487
rect 239036 237448 239088 237454
rect 239036 237390 239088 237396
rect 239048 234462 239076 237390
rect 239140 237386 239168 238734
rect 239312 238128 239364 238134
rect 239312 238070 239364 238076
rect 239220 237856 239272 237862
rect 239220 237798 239272 237804
rect 239232 237590 239260 237798
rect 239220 237584 239272 237590
rect 239220 237526 239272 237532
rect 239324 237522 239352 238070
rect 239312 237516 239364 237522
rect 239312 237458 239364 237464
rect 239128 237380 239180 237386
rect 239128 237322 239180 237328
rect 239220 235408 239272 235414
rect 239220 235350 239272 235356
rect 239036 234456 239088 234462
rect 239036 234398 239088 234404
rect 239128 234116 239180 234122
rect 239128 234058 239180 234064
rect 238944 232620 238996 232626
rect 238944 232562 238996 232568
rect 239140 229906 239168 234058
rect 239128 229900 239180 229906
rect 239128 229842 239180 229848
rect 239232 226234 239260 235350
rect 239312 235204 239364 235210
rect 239312 235146 239364 235152
rect 239036 226228 239088 226234
rect 239036 226170 239088 226176
rect 239220 226228 239272 226234
rect 239220 226170 239272 226176
rect 239048 225826 239076 226170
rect 239036 225820 239088 225826
rect 239036 225762 239088 225768
rect 239324 224262 239352 235146
rect 239416 235142 239444 239720
rect 239588 239624 239640 239630
rect 239588 239566 239640 239572
rect 239496 238128 239548 238134
rect 239496 238070 239548 238076
rect 239404 235136 239456 235142
rect 239404 235078 239456 235084
rect 239416 230926 239444 235078
rect 239404 230920 239456 230926
rect 239404 230862 239456 230868
rect 239404 230240 239456 230246
rect 239404 230182 239456 230188
rect 239312 224256 239364 224262
rect 239312 224198 239364 224204
rect 238850 213888 238906 213897
rect 238850 213823 238906 213832
rect 238574 159488 238630 159497
rect 238574 159423 238630 159432
rect 238482 154320 238538 154329
rect 238482 154255 238538 154264
rect 238392 149932 238444 149938
rect 238392 149874 238444 149880
rect 239416 146878 239444 230182
rect 239404 146872 239456 146878
rect 239404 146814 239456 146820
rect 238298 144120 238354 144129
rect 238298 144055 238354 144064
rect 238024 136400 238076 136406
rect 238024 136342 238076 136348
rect 237380 129056 237432 129062
rect 237380 128998 237432 129004
rect 237392 16574 237420 128998
rect 236012 16546 236592 16574
rect 237392 16546 237696 16574
rect 235264 4072 235316 4078
rect 235264 4014 235316 4020
rect 235816 3936 235868 3942
rect 235816 3878 235868 3884
rect 235828 480 235856 3878
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 16546
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 237668 354 237696 16546
rect 239312 3800 239364 3806
rect 239312 3742 239364 3748
rect 239324 480 239352 3742
rect 239416 3398 239444 146814
rect 239508 141681 239536 238070
rect 239600 233374 239628 239566
rect 239692 234122 239720 239720
rect 239784 235414 239812 239788
rect 239922 239680 239950 240108
rect 240014 239970 240042 240108
rect 240002 239964 240054 239970
rect 240002 239906 240054 239912
rect 240106 239816 240134 240108
rect 240198 239970 240226 240108
rect 240186 239964 240238 239970
rect 240186 239906 240238 239912
rect 240290 239850 240318 240108
rect 240382 239873 240410 240108
rect 240474 239970 240502 240108
rect 240462 239964 240514 239970
rect 240462 239906 240514 239912
rect 240244 239822 240318 239850
rect 240368 239864 240424 239873
rect 240106 239788 240180 239816
rect 240048 239692 240100 239698
rect 239922 239652 239996 239680
rect 239772 235408 239824 235414
rect 239772 235350 239824 235356
rect 239680 234116 239732 234122
rect 239680 234058 239732 234064
rect 239968 233782 239996 239652
rect 240048 239634 240100 239640
rect 240060 235210 240088 239634
rect 240152 238785 240180 239788
rect 240138 238776 240194 238785
rect 240138 238711 240194 238720
rect 240244 237930 240272 239822
rect 240566 239816 240594 240108
rect 240658 239902 240686 240108
rect 240750 239970 240778 240108
rect 240738 239964 240790 239970
rect 240738 239906 240790 239912
rect 240646 239896 240698 239902
rect 240842 239873 240870 240108
rect 240934 239970 240962 240108
rect 241026 239970 241054 240108
rect 240922 239964 240974 239970
rect 240922 239906 240974 239912
rect 241014 239964 241066 239970
rect 241014 239906 241066 239912
rect 240646 239838 240698 239844
rect 240828 239864 240884 239873
rect 240368 239799 240424 239808
rect 240520 239788 240594 239816
rect 240828 239799 240884 239808
rect 240968 239828 241020 239834
rect 240324 239760 240376 239766
rect 240520 239748 240548 239788
rect 240968 239770 241020 239776
rect 240324 239702 240376 239708
rect 240428 239720 240548 239748
rect 240784 239760 240836 239766
rect 240336 238649 240364 239702
rect 240322 238640 240378 238649
rect 240322 238575 240378 238584
rect 240232 237924 240284 237930
rect 240232 237866 240284 237872
rect 240232 237788 240284 237794
rect 240232 237730 240284 237736
rect 240140 237720 240192 237726
rect 240140 237662 240192 237668
rect 240048 235204 240100 235210
rect 240048 235146 240100 235152
rect 239956 233776 240008 233782
rect 239956 233718 240008 233724
rect 239588 233368 239640 233374
rect 239588 233310 239640 233316
rect 239600 230474 239628 233310
rect 239600 230446 239720 230474
rect 239588 229560 239640 229566
rect 239588 229502 239640 229508
rect 239600 152794 239628 229502
rect 239692 228410 239720 230446
rect 239968 229974 239996 233718
rect 240152 233234 240180 237662
rect 240244 235822 240272 237730
rect 240232 235816 240284 235822
rect 240232 235758 240284 235764
rect 240060 233206 240180 233234
rect 240060 230246 240088 233206
rect 240048 230240 240100 230246
rect 240048 230182 240100 230188
rect 240428 230110 240456 239720
rect 240784 239702 240836 239708
rect 240876 239760 240928 239766
rect 240876 239702 240928 239708
rect 240692 239692 240744 239698
rect 240692 239634 240744 239640
rect 240600 239488 240652 239494
rect 240600 239430 240652 239436
rect 240508 238332 240560 238338
rect 240508 238274 240560 238280
rect 240520 237930 240548 238274
rect 240508 237924 240560 237930
rect 240508 237866 240560 237872
rect 240612 237368 240640 239430
rect 240704 238785 240732 239634
rect 240690 238776 240746 238785
rect 240690 238711 240746 238720
rect 240520 237340 240640 237368
rect 240416 230104 240468 230110
rect 240416 230046 240468 230052
rect 240520 230042 240548 237340
rect 240600 237244 240652 237250
rect 240600 237186 240652 237192
rect 240612 234598 240640 237186
rect 240600 234592 240652 234598
rect 240600 234534 240652 234540
rect 240704 233889 240732 238711
rect 240796 238542 240824 239702
rect 240784 238536 240836 238542
rect 240784 238478 240836 238484
rect 240796 235074 240824 238478
rect 240888 238241 240916 239702
rect 240874 238232 240930 238241
rect 240874 238167 240930 238176
rect 240784 235068 240836 235074
rect 240784 235010 240836 235016
rect 240888 234297 240916 238167
rect 240874 234288 240930 234297
rect 240874 234223 240930 234232
rect 240690 233880 240746 233889
rect 240690 233815 240746 233824
rect 240980 233234 241008 239770
rect 241118 239748 241146 240108
rect 241210 239907 241238 240108
rect 241196 239898 241252 239907
rect 241302 239902 241330 240108
rect 241196 239833 241252 239842
rect 241290 239896 241342 239902
rect 241290 239838 241342 239844
rect 241394 239748 241422 240108
rect 241486 239970 241514 240108
rect 241578 239970 241606 240108
rect 241670 239970 241698 240108
rect 241762 239970 241790 240108
rect 241474 239964 241526 239970
rect 241474 239906 241526 239912
rect 241566 239964 241618 239970
rect 241566 239906 241618 239912
rect 241658 239964 241710 239970
rect 241658 239906 241710 239912
rect 241750 239964 241802 239970
rect 241750 239906 241802 239912
rect 241702 239864 241758 239873
rect 241854 239850 241882 240108
rect 241946 239970 241974 240108
rect 241934 239964 241986 239970
rect 241934 239906 241986 239912
rect 241854 239822 241928 239850
rect 241702 239799 241758 239808
rect 241900 239816 241928 239822
rect 240690 233200 240746 233209
rect 240690 233135 240746 233144
rect 240796 233206 241008 233234
rect 241072 239720 241146 239748
rect 241348 239720 241422 239748
rect 240508 230036 240560 230042
rect 240508 229978 240560 229984
rect 239956 229968 240008 229974
rect 239956 229910 240008 229916
rect 239680 228404 239732 228410
rect 239680 228346 239732 228352
rect 239680 227520 239732 227526
rect 239680 227462 239732 227468
rect 239692 157185 239720 227462
rect 239772 226976 239824 226982
rect 239772 226918 239824 226924
rect 239784 159361 239812 226918
rect 240704 224777 240732 233135
rect 240796 232762 240824 233206
rect 240784 232756 240836 232762
rect 240784 232698 240836 232704
rect 240796 228750 240824 232698
rect 241072 232098 241100 239720
rect 241244 239692 241296 239698
rect 241244 239634 241296 239640
rect 241152 239216 241204 239222
rect 241152 239158 241204 239164
rect 241164 238950 241192 239158
rect 241152 238944 241204 238950
rect 241152 238886 241204 238892
rect 241150 238640 241206 238649
rect 241150 238575 241206 238584
rect 240980 232070 241100 232098
rect 240784 228744 240836 228750
rect 240784 228686 240836 228692
rect 240876 226840 240928 226846
rect 240876 226782 240928 226788
rect 240690 224768 240746 224777
rect 240690 224703 240746 224712
rect 240048 224528 240100 224534
rect 240048 224470 240100 224476
rect 240060 224262 240088 224470
rect 240784 224460 240836 224466
rect 240784 224402 240836 224408
rect 240048 224256 240100 224262
rect 240048 224198 240100 224204
rect 239770 159352 239826 159361
rect 239770 159287 239826 159296
rect 239678 157176 239734 157185
rect 239678 157111 239734 157120
rect 240140 156936 240192 156942
rect 240140 156878 240192 156884
rect 239588 152788 239640 152794
rect 239588 152730 239640 152736
rect 239494 141672 239550 141681
rect 239494 141607 239550 141616
rect 239404 3392 239456 3398
rect 239404 3334 239456 3340
rect 238086 354 238198 480
rect 237668 326 238198 354
rect 236982 -960 237094 326
rect 238086 -960 238198 326
rect 239282 -960 239394 480
rect 240152 354 240180 156878
rect 240796 151502 240824 224402
rect 240888 154193 240916 226782
rect 240980 224398 241008 232070
rect 241060 232008 241112 232014
rect 241060 231950 241112 231956
rect 240968 224392 241020 224398
rect 240968 224334 241020 224340
rect 240980 156942 241008 224334
rect 241072 224262 241100 231950
rect 241060 224256 241112 224262
rect 241060 224198 241112 224204
rect 241164 221649 241192 238575
rect 241256 236745 241284 239634
rect 241242 236736 241298 236745
rect 241242 236671 241298 236680
rect 241244 234048 241296 234054
rect 241244 233990 241296 233996
rect 241256 229094 241284 233990
rect 241348 232014 241376 239720
rect 241520 239692 241572 239698
rect 241520 239634 241572 239640
rect 241612 239692 241664 239698
rect 241612 239634 241664 239640
rect 241532 239358 241560 239634
rect 241520 239352 241572 239358
rect 241520 239294 241572 239300
rect 241428 239284 241480 239290
rect 241428 239226 241480 239232
rect 241440 238746 241468 239226
rect 241428 238740 241480 238746
rect 241428 238682 241480 238688
rect 241426 238640 241482 238649
rect 241426 238575 241482 238584
rect 241440 238105 241468 238575
rect 241520 238536 241572 238542
rect 241520 238478 241572 238484
rect 241532 238406 241560 238478
rect 241520 238400 241572 238406
rect 241520 238342 241572 238348
rect 241426 238096 241482 238105
rect 241426 238031 241482 238040
rect 241624 234614 241652 239634
rect 241716 237726 241744 239799
rect 241900 239788 241974 239816
rect 241796 239760 241848 239766
rect 241946 239714 241974 239788
rect 242038 239748 242066 240108
rect 242130 239873 242158 240108
rect 242116 239864 242172 239873
rect 242116 239799 242172 239808
rect 242038 239720 242112 239748
rect 241796 239702 241848 239708
rect 241704 237720 241756 237726
rect 241704 237662 241756 237668
rect 241704 236768 241756 236774
rect 241704 236710 241756 236716
rect 241440 234586 241652 234614
rect 241336 232008 241388 232014
rect 241336 231950 241388 231956
rect 241256 229066 241376 229094
rect 241242 226400 241298 226409
rect 241242 226335 241298 226344
rect 241150 221640 241206 221649
rect 241150 221575 241206 221584
rect 240968 156936 241020 156942
rect 240968 156878 241020 156884
rect 240874 154184 240930 154193
rect 240874 154119 240930 154128
rect 240784 151496 240836 151502
rect 240784 151438 240836 151444
rect 240796 2990 240824 151438
rect 241256 3262 241284 226335
rect 241348 152930 241376 229066
rect 241440 224466 241468 234586
rect 241716 234308 241744 236710
rect 241808 234433 241836 239702
rect 241900 239686 241974 239714
rect 241900 236745 241928 239686
rect 241980 239556 242032 239562
rect 241980 239498 242032 239504
rect 241886 236736 241942 236745
rect 241886 236671 241942 236680
rect 241888 236564 241940 236570
rect 241888 236506 241940 236512
rect 241794 234424 241850 234433
rect 241794 234359 241850 234368
rect 241716 234280 241836 234308
rect 241704 233912 241756 233918
rect 241704 233854 241756 233860
rect 241520 229628 241572 229634
rect 241520 229570 241572 229576
rect 241612 229628 241664 229634
rect 241612 229570 241664 229576
rect 241532 229362 241560 229570
rect 241520 229356 241572 229362
rect 241520 229298 241572 229304
rect 241428 224460 241480 224466
rect 241428 224402 241480 224408
rect 241520 224256 241572 224262
rect 241520 224198 241572 224204
rect 241336 152924 241388 152930
rect 241336 152866 241388 152872
rect 241532 151162 241560 224198
rect 241624 224194 241652 229570
rect 241716 225010 241744 233854
rect 241808 225554 241836 234280
rect 241900 226302 241928 236506
rect 241992 227089 242020 239498
rect 242084 236638 242112 239720
rect 242222 239714 242250 240108
rect 242314 239970 242342 240108
rect 242406 239970 242434 240108
rect 242498 239970 242526 240108
rect 242302 239964 242354 239970
rect 242302 239906 242354 239912
rect 242394 239964 242446 239970
rect 242394 239906 242446 239912
rect 242486 239964 242538 239970
rect 242486 239906 242538 239912
rect 242590 239816 242618 240108
rect 242176 239686 242250 239714
rect 242544 239788 242618 239816
rect 242072 236632 242124 236638
rect 242072 236574 242124 236580
rect 242176 229634 242204 239686
rect 242348 239556 242400 239562
rect 242348 239498 242400 239504
rect 242256 239148 242308 239154
rect 242256 239090 242308 239096
rect 242268 236774 242296 239090
rect 242256 236768 242308 236774
rect 242256 236710 242308 236716
rect 242256 236632 242308 236638
rect 242256 236574 242308 236580
rect 242164 229628 242216 229634
rect 242164 229570 242216 229576
rect 241978 227080 242034 227089
rect 241978 227015 242034 227024
rect 241992 226409 242020 227015
rect 241978 226400 242034 226409
rect 241978 226335 242034 226344
rect 241888 226296 241940 226302
rect 241888 226238 241940 226244
rect 241796 225548 241848 225554
rect 241796 225490 241848 225496
rect 241704 225004 241756 225010
rect 241704 224946 241756 224952
rect 241612 224188 241664 224194
rect 241612 224130 241664 224136
rect 241808 219434 241836 225490
rect 241900 225486 241928 226238
rect 241888 225480 241940 225486
rect 241888 225422 241940 225428
rect 242268 223281 242296 236574
rect 242360 234054 242388 239498
rect 242440 239488 242492 239494
rect 242440 239430 242492 239436
rect 242452 236570 242480 239430
rect 242544 239154 242572 239788
rect 242682 239748 242710 240108
rect 242774 239816 242802 240108
rect 242866 239970 242894 240108
rect 242854 239964 242906 239970
rect 242854 239906 242906 239912
rect 242958 239816 242986 240108
rect 243050 239970 243078 240108
rect 243038 239964 243090 239970
rect 243038 239906 243090 239912
rect 243142 239907 243170 240108
rect 243128 239898 243184 239907
rect 243128 239833 243184 239842
rect 243234 239816 243262 240108
rect 243326 239970 243354 240108
rect 243314 239964 243366 239970
rect 243314 239906 243366 239912
rect 243418 239816 243446 240108
rect 243510 239970 243538 240108
rect 243498 239964 243550 239970
rect 243498 239906 243550 239912
rect 243602 239850 243630 240108
rect 243694 239902 243722 240108
rect 242774 239788 242848 239816
rect 242958 239788 243032 239816
rect 243234 239788 243308 239816
rect 242636 239720 242710 239748
rect 242820 239748 242848 239788
rect 243004 239748 243032 239788
rect 242820 239720 242940 239748
rect 243004 239720 243124 239748
rect 243280 239737 243308 239788
rect 243372 239788 243446 239816
rect 243556 239822 243630 239850
rect 243682 239896 243734 239902
rect 243682 239838 243734 239844
rect 242532 239148 242584 239154
rect 242532 239090 242584 239096
rect 242532 239012 242584 239018
rect 242532 238954 242584 238960
rect 242544 238066 242572 238954
rect 242532 238060 242584 238066
rect 242532 238002 242584 238008
rect 242440 236564 242492 236570
rect 242440 236506 242492 236512
rect 242348 234048 242400 234054
rect 242348 233990 242400 233996
rect 242636 229974 242664 239720
rect 242912 239680 242940 239720
rect 242912 239652 243032 239680
rect 242808 239556 242860 239562
rect 242808 239498 242860 239504
rect 242900 239556 242952 239562
rect 242900 239498 242952 239504
rect 242716 239420 242768 239426
rect 242716 239362 242768 239368
rect 242728 233918 242756 239362
rect 242820 235550 242848 239498
rect 242912 239465 242940 239498
rect 242898 239456 242954 239465
rect 243004 239426 243032 239652
rect 242898 239391 242954 239400
rect 242992 239420 243044 239426
rect 242992 239362 243044 239368
rect 242900 239080 242952 239086
rect 242900 239022 242952 239028
rect 242912 238678 242940 239022
rect 242900 238672 242952 238678
rect 242900 238614 242952 238620
rect 243096 235929 243124 239720
rect 243266 239728 243322 239737
rect 243176 239692 243228 239698
rect 243266 239663 243322 239672
rect 243176 239634 243228 239640
rect 243082 235920 243138 235929
rect 243082 235855 243138 235864
rect 242808 235544 242860 235550
rect 242808 235486 242860 235492
rect 242820 234161 242848 235486
rect 243096 235385 243124 235855
rect 243188 235414 243216 239634
rect 243268 239624 243320 239630
rect 243268 239566 243320 239572
rect 243280 239465 243308 239566
rect 243266 239456 243322 239465
rect 243266 239391 243322 239400
rect 243268 239352 243320 239358
rect 243268 239294 243320 239300
rect 243280 236881 243308 239294
rect 243266 236872 243322 236881
rect 243266 236807 243322 236816
rect 243176 235408 243228 235414
rect 243082 235376 243138 235385
rect 243176 235350 243228 235356
rect 243082 235311 243138 235320
rect 243084 235204 243136 235210
rect 243084 235146 243136 235152
rect 242806 234152 242862 234161
rect 242806 234087 242862 234096
rect 242716 233912 242768 233918
rect 242716 233854 242768 233860
rect 242992 233436 243044 233442
rect 242992 233378 243044 233384
rect 242624 229968 242676 229974
rect 242624 229910 242676 229916
rect 242636 229094 242664 229910
rect 242636 229066 242756 229094
rect 242532 225480 242584 225486
rect 242532 225422 242584 225428
rect 242254 223272 242310 223281
rect 242254 223207 242310 223216
rect 241808 219406 242204 219434
rect 242176 159594 242204 219406
rect 242164 159588 242216 159594
rect 242164 159530 242216 159536
rect 241520 151156 241572 151162
rect 241520 151098 241572 151104
rect 241532 150482 241560 151098
rect 241520 150476 241572 150482
rect 241520 150418 241572 150424
rect 242164 150476 242216 150482
rect 242164 150418 242216 150424
rect 241520 134632 241572 134638
rect 241520 134574 241572 134580
rect 241532 16574 241560 134574
rect 241532 16546 241744 16574
rect 241244 3256 241296 3262
rect 241244 3198 241296 3204
rect 240784 2984 240836 2990
rect 240784 2926 240836 2932
rect 241716 480 241744 16546
rect 242176 2922 242204 150418
rect 242268 142089 242296 223207
rect 242544 213314 242572 225422
rect 242624 225412 242676 225418
rect 242624 225354 242676 225360
rect 242636 225010 242664 225354
rect 242624 225004 242676 225010
rect 242624 224946 242676 224952
rect 242532 213308 242584 213314
rect 242532 213250 242584 213256
rect 242636 184210 242664 224946
rect 242624 184204 242676 184210
rect 242624 184146 242676 184152
rect 242728 151638 242756 229066
rect 242806 225040 242862 225049
rect 242806 224975 242862 224984
rect 242716 151632 242768 151638
rect 242716 151574 242768 151580
rect 242728 150482 242756 151574
rect 242716 150476 242768 150482
rect 242716 150418 242768 150424
rect 242254 142080 242310 142089
rect 242254 142015 242310 142024
rect 242820 4078 242848 224975
rect 243004 222154 243032 233378
rect 243096 225962 243124 235146
rect 243372 233617 243400 239788
rect 243450 239728 243506 239737
rect 243450 239663 243506 239672
rect 243464 234530 243492 239663
rect 243556 235210 243584 239822
rect 243636 239760 243688 239766
rect 243786 239748 243814 240108
rect 243636 239702 243688 239708
rect 243740 239720 243814 239748
rect 243544 235204 243596 235210
rect 243544 235146 243596 235152
rect 243452 234524 243504 234530
rect 243452 234466 243504 234472
rect 243358 233608 243414 233617
rect 243358 233543 243414 233552
rect 243084 225956 243136 225962
rect 243084 225898 243136 225904
rect 243096 225486 243124 225898
rect 243084 225480 243136 225486
rect 243084 225422 243136 225428
rect 242992 222148 243044 222154
rect 242992 222090 243044 222096
rect 243464 147422 243492 234466
rect 243648 233442 243676 239702
rect 243740 238338 243768 239720
rect 243878 239680 243906 240108
rect 243970 239748 243998 240108
rect 244062 239850 244090 240108
rect 244154 239970 244182 240108
rect 244142 239964 244194 239970
rect 244142 239906 244194 239912
rect 244062 239822 244136 239850
rect 243970 239720 244044 239748
rect 243832 239652 243906 239680
rect 243728 238332 243780 238338
rect 243728 238274 243780 238280
rect 243728 238196 243780 238202
rect 243728 238138 243780 238144
rect 243740 237726 243768 238138
rect 243728 237720 243780 237726
rect 243728 237662 243780 237668
rect 243728 237312 243780 237318
rect 243728 237254 243780 237260
rect 243740 233918 243768 237254
rect 243832 237182 243860 239652
rect 244016 239578 244044 239720
rect 243924 239550 244044 239578
rect 243820 237176 243872 237182
rect 243820 237118 243872 237124
rect 243820 235476 243872 235482
rect 243820 235418 243872 235424
rect 243728 233912 243780 233918
rect 243728 233854 243780 233860
rect 243636 233436 243688 233442
rect 243636 233378 243688 233384
rect 243740 230178 243768 233854
rect 243728 230172 243780 230178
rect 243728 230114 243780 230120
rect 243544 225480 243596 225486
rect 243544 225422 243596 225428
rect 243556 151434 243584 225422
rect 243728 224120 243780 224126
rect 243728 224062 243780 224068
rect 243636 222148 243688 222154
rect 243636 222090 243688 222096
rect 243648 221678 243676 222090
rect 243636 221672 243688 221678
rect 243636 221614 243688 221620
rect 243648 158914 243676 221614
rect 243636 158908 243688 158914
rect 243636 158850 243688 158856
rect 243544 151428 243596 151434
rect 243544 151370 243596 151376
rect 243452 147416 243504 147422
rect 243452 147358 243504 147364
rect 243464 146946 243492 147358
rect 243452 146940 243504 146946
rect 243452 146882 243504 146888
rect 242808 4072 242860 4078
rect 242808 4014 242860 4020
rect 243556 3874 243584 151370
rect 243636 150476 243688 150482
rect 243636 150418 243688 150424
rect 243648 3942 243676 150418
rect 243740 148714 243768 224062
rect 243728 148708 243780 148714
rect 243728 148650 243780 148656
rect 243636 3936 243688 3942
rect 243636 3878 243688 3884
rect 243544 3868 243596 3874
rect 243544 3810 243596 3816
rect 243740 3806 243768 148650
rect 243832 143274 243860 235418
rect 243924 219026 243952 239550
rect 244004 239488 244056 239494
rect 244004 239430 244056 239436
rect 244016 237318 244044 239430
rect 244004 237312 244056 237318
rect 244004 237254 244056 237260
rect 244004 236632 244056 236638
rect 244004 236574 244056 236580
rect 244016 224126 244044 236574
rect 244108 231470 244136 239822
rect 244246 239816 244274 240108
rect 244200 239788 244274 239816
rect 244200 237454 244228 239788
rect 244338 239748 244366 240108
rect 244430 239970 244458 240108
rect 244418 239964 244470 239970
rect 244418 239906 244470 239912
rect 244522 239850 244550 240108
rect 244614 239970 244642 240108
rect 244706 239970 244734 240108
rect 244798 239970 244826 240108
rect 244602 239964 244654 239970
rect 244602 239906 244654 239912
rect 244694 239964 244746 239970
rect 244694 239906 244746 239912
rect 244786 239964 244838 239970
rect 244786 239906 244838 239912
rect 244292 239720 244366 239748
rect 244476 239822 244550 239850
rect 244738 239864 244794 239873
rect 244188 237448 244240 237454
rect 244188 237390 244240 237396
rect 244292 237300 244320 239720
rect 244476 239544 244504 239822
rect 244890 239816 244918 240108
rect 244982 239834 245010 240108
rect 245074 239970 245102 240108
rect 245062 239964 245114 239970
rect 245062 239906 245114 239912
rect 244738 239799 244740 239808
rect 244792 239799 244794 239808
rect 244740 239770 244792 239776
rect 244844 239788 244918 239816
rect 244970 239828 245022 239834
rect 244556 239760 244608 239766
rect 244556 239702 244608 239708
rect 244200 237272 244320 237300
rect 244384 239516 244504 239544
rect 244200 232694 244228 237272
rect 244384 237232 244412 239516
rect 244462 239456 244518 239465
rect 244462 239391 244518 239400
rect 244292 237204 244412 237232
rect 244292 234326 244320 237204
rect 244372 237108 244424 237114
rect 244372 237050 244424 237056
rect 244280 234320 244332 234326
rect 244280 234262 244332 234268
rect 244188 232688 244240 232694
rect 244188 232630 244240 232636
rect 244096 231464 244148 231470
rect 244096 231406 244148 231412
rect 244200 231282 244228 232630
rect 244108 231254 244228 231282
rect 244004 224120 244056 224126
rect 244004 224062 244056 224068
rect 243912 219020 243964 219026
rect 243912 218962 243964 218968
rect 243924 213489 243952 218962
rect 243910 213480 243966 213489
rect 243910 213415 243966 213424
rect 244108 148850 244136 231254
rect 244280 230444 244332 230450
rect 244280 230386 244332 230392
rect 244292 230314 244320 230386
rect 244188 230308 244240 230314
rect 244188 230250 244240 230256
rect 244280 230308 244332 230314
rect 244280 230250 244332 230256
rect 244200 229158 244228 230250
rect 244188 229152 244240 229158
rect 244188 229094 244240 229100
rect 244200 225758 244228 229094
rect 244188 225752 244240 225758
rect 244188 225694 244240 225700
rect 244384 213246 244412 237050
rect 244476 227594 244504 239391
rect 244568 233234 244596 239702
rect 244648 239692 244700 239698
rect 244648 239634 244700 239640
rect 244660 236638 244688 239634
rect 244752 238241 244780 239770
rect 244738 238232 244794 238241
rect 244738 238167 244794 238176
rect 244740 237040 244792 237046
rect 244740 236982 244792 236988
rect 244648 236632 244700 236638
rect 244648 236574 244700 236580
rect 244648 236020 244700 236026
rect 244648 235962 244700 235968
rect 244660 234598 244688 235962
rect 244752 235618 244780 236982
rect 244740 235612 244792 235618
rect 244740 235554 244792 235560
rect 244752 235346 244780 235554
rect 244740 235340 244792 235346
rect 244740 235282 244792 235288
rect 244648 234592 244700 234598
rect 244648 234534 244700 234540
rect 244568 233206 244688 233234
rect 244660 229770 244688 233206
rect 244844 229906 244872 239788
rect 245166 239816 245194 240108
rect 244970 239770 245022 239776
rect 245120 239788 245194 239816
rect 245120 239714 245148 239788
rect 245258 239748 245286 240108
rect 245350 239970 245378 240108
rect 245442 239970 245470 240108
rect 245338 239964 245390 239970
rect 245338 239906 245390 239912
rect 245430 239964 245482 239970
rect 245430 239906 245482 239912
rect 245382 239864 245438 239873
rect 245382 239799 245438 239808
rect 244924 239692 244976 239698
rect 245074 239686 245148 239714
rect 245212 239720 245286 239748
rect 245074 239680 245102 239686
rect 244924 239634 244976 239640
rect 245028 239652 245102 239680
rect 244936 237046 244964 239634
rect 244924 237040 244976 237046
rect 244924 236982 244976 236988
rect 244924 236768 244976 236774
rect 244924 236710 244976 236716
rect 244936 235754 244964 236710
rect 244924 235748 244976 235754
rect 244924 235690 244976 235696
rect 244832 229900 244884 229906
rect 244832 229842 244884 229848
rect 244648 229764 244700 229770
rect 244648 229706 244700 229712
rect 244464 227588 244516 227594
rect 244464 227530 244516 227536
rect 244372 213240 244424 213246
rect 244372 213182 244424 213188
rect 244936 150074 244964 235690
rect 245028 228206 245056 239652
rect 245108 239352 245160 239358
rect 245108 239294 245160 239300
rect 245120 237114 245148 239294
rect 245108 237108 245160 237114
rect 245108 237050 245160 237056
rect 245212 236774 245240 239720
rect 245292 239624 245344 239630
rect 245292 239566 245344 239572
rect 245304 239465 245332 239566
rect 245396 239562 245424 239799
rect 245534 239748 245562 240108
rect 245626 239850 245654 240108
rect 245718 239970 245746 240108
rect 245706 239964 245758 239970
rect 245706 239906 245758 239912
rect 245810 239902 245838 240108
rect 245798 239896 245850 239902
rect 245626 239822 245700 239850
rect 245798 239838 245850 239844
rect 245902 239850 245930 240108
rect 245994 239970 246022 240108
rect 245982 239964 246034 239970
rect 245982 239906 246034 239912
rect 246086 239850 246114 240108
rect 246178 239970 246206 240108
rect 246166 239964 246218 239970
rect 246166 239906 246218 239912
rect 245902 239822 245976 239850
rect 245534 239720 245608 239748
rect 245672 239737 245700 239822
rect 245752 239760 245804 239766
rect 245476 239624 245528 239630
rect 245476 239566 245528 239572
rect 245384 239556 245436 239562
rect 245384 239498 245436 239504
rect 245290 239456 245346 239465
rect 245290 239391 245346 239400
rect 245382 238640 245438 238649
rect 245382 238575 245438 238584
rect 245200 236768 245252 236774
rect 245200 236710 245252 236716
rect 245108 236292 245160 236298
rect 245108 236234 245160 236240
rect 245120 230450 245148 236234
rect 245396 234614 245424 238575
rect 245488 238066 245516 239566
rect 245476 238060 245528 238066
rect 245476 238002 245528 238008
rect 245580 236298 245608 239720
rect 245658 239728 245714 239737
rect 245752 239702 245804 239708
rect 245844 239760 245896 239766
rect 245844 239702 245896 239708
rect 245658 239663 245714 239672
rect 245660 239216 245712 239222
rect 245660 239158 245712 239164
rect 245672 238542 245700 239158
rect 245660 238536 245712 238542
rect 245660 238478 245712 238484
rect 245568 236292 245620 236298
rect 245568 236234 245620 236240
rect 245568 234864 245620 234870
rect 245568 234806 245620 234812
rect 245304 234586 245424 234614
rect 245108 230444 245160 230450
rect 245108 230386 245160 230392
rect 245200 230308 245252 230314
rect 245200 230250 245252 230256
rect 245212 229906 245240 230250
rect 245200 229900 245252 229906
rect 245200 229842 245252 229848
rect 245016 228200 245068 228206
rect 245016 228142 245068 228148
rect 245016 168428 245068 168434
rect 245016 168370 245068 168376
rect 244924 150068 244976 150074
rect 244924 150010 244976 150016
rect 244096 148844 244148 148850
rect 244096 148786 244148 148792
rect 245028 148646 245056 168370
rect 245016 148640 245068 148646
rect 245016 148582 245068 148588
rect 243820 143268 243872 143274
rect 243820 143210 243872 143216
rect 243832 141574 243860 143210
rect 245212 141846 245240 229842
rect 245304 168434 245332 234586
rect 245384 233300 245436 233306
rect 245384 233242 245436 233248
rect 245292 168428 245344 168434
rect 245292 168370 245344 168376
rect 245396 151570 245424 233242
rect 245476 229764 245528 229770
rect 245476 229706 245528 229712
rect 245488 229634 245516 229706
rect 245476 229628 245528 229634
rect 245476 229570 245528 229576
rect 245384 151564 245436 151570
rect 245384 151506 245436 151512
rect 245396 151162 245424 151506
rect 245384 151156 245436 151162
rect 245384 151098 245436 151104
rect 245488 146062 245516 229570
rect 245580 225826 245608 234806
rect 245764 234462 245792 239702
rect 245856 234870 245884 239702
rect 245844 234864 245896 234870
rect 245844 234806 245896 234812
rect 245752 234456 245804 234462
rect 245752 234398 245804 234404
rect 245764 233306 245792 234398
rect 245752 233300 245804 233306
rect 245752 233242 245804 233248
rect 245948 233209 245976 239822
rect 246040 239822 246114 239850
rect 245934 233200 245990 233209
rect 245934 233135 245990 233144
rect 246040 229770 246068 239822
rect 246270 239816 246298 240108
rect 246362 239907 246390 240108
rect 246348 239898 246404 239907
rect 246454 239902 246482 240108
rect 246348 239833 246404 239842
rect 246442 239896 246494 239902
rect 246442 239838 246494 239844
rect 246224 239788 246298 239816
rect 246120 239760 246172 239766
rect 246120 239702 246172 239708
rect 246132 233238 246160 239702
rect 246120 233232 246172 233238
rect 246120 233174 246172 233180
rect 246224 233034 246252 239788
rect 246396 239760 246448 239766
rect 246394 239728 246396 239737
rect 246448 239728 246450 239737
rect 246304 239692 246356 239698
rect 246394 239663 246450 239672
rect 246546 239680 246574 240108
rect 246638 239970 246666 240108
rect 246730 239970 246758 240108
rect 246626 239964 246678 239970
rect 246626 239906 246678 239912
rect 246718 239964 246770 239970
rect 246718 239906 246770 239912
rect 246822 239816 246850 240108
rect 246684 239788 246850 239816
rect 246546 239652 246620 239680
rect 246304 239634 246356 239640
rect 246316 239154 246344 239634
rect 246488 239556 246540 239562
rect 246488 239498 246540 239504
rect 246396 239488 246448 239494
rect 246396 239430 246448 239436
rect 246304 239148 246356 239154
rect 246304 239090 246356 239096
rect 246408 233850 246436 239430
rect 246500 234802 246528 239498
rect 246488 234796 246540 234802
rect 246488 234738 246540 234744
rect 246396 233844 246448 233850
rect 246396 233786 246448 233792
rect 246212 233028 246264 233034
rect 246212 232970 246264 232976
rect 246224 230874 246252 232970
rect 246132 230846 246252 230874
rect 246028 229764 246080 229770
rect 246028 229706 246080 229712
rect 246132 225894 246160 230846
rect 246592 229906 246620 239652
rect 246684 238610 246712 239788
rect 246914 239748 246942 240108
rect 247006 239873 247034 240108
rect 246992 239864 247048 239873
rect 246992 239799 247048 239808
rect 247098 239748 247126 240108
rect 246776 239720 246942 239748
rect 247052 239720 247126 239748
rect 246672 238604 246724 238610
rect 246672 238546 246724 238552
rect 246672 233232 246724 233238
rect 246672 233174 246724 233180
rect 246212 229900 246264 229906
rect 246212 229842 246264 229848
rect 246580 229900 246632 229906
rect 246580 229842 246632 229848
rect 246120 225888 246172 225894
rect 246120 225830 246172 225836
rect 245568 225820 245620 225826
rect 245568 225762 245620 225768
rect 246224 224954 246252 229842
rect 246580 229764 246632 229770
rect 246580 229706 246632 229712
rect 246488 226160 246540 226166
rect 246488 226102 246540 226108
rect 246500 225690 246528 226102
rect 246488 225684 246540 225690
rect 246488 225626 246540 225632
rect 246224 224926 246344 224954
rect 246316 161022 246344 224926
rect 246396 219292 246448 219298
rect 246396 219234 246448 219240
rect 246304 161016 246356 161022
rect 246304 160958 246356 160964
rect 246304 152924 246356 152930
rect 246304 152866 246356 152872
rect 245476 146056 245528 146062
rect 245476 145998 245528 146004
rect 245200 141840 245252 141846
rect 245200 141782 245252 141788
rect 243820 141568 243872 141574
rect 243820 141510 243872 141516
rect 245212 141506 245240 141782
rect 245200 141500 245252 141506
rect 245200 141442 245252 141448
rect 246028 133748 246080 133754
rect 246028 133690 246080 133696
rect 246040 133346 246068 133690
rect 246028 133340 246080 133346
rect 246028 133282 246080 133288
rect 244278 122224 244334 122233
rect 244278 122159 244334 122168
rect 244292 16574 244320 122159
rect 244292 16546 245240 16574
rect 243728 3800 243780 3806
rect 243728 3742 243780 3748
rect 242900 3664 242952 3670
rect 242900 3606 242952 3612
rect 242164 2916 242216 2922
rect 242164 2858 242216 2864
rect 242912 480 242940 3606
rect 244096 2916 244148 2922
rect 244096 2858 244148 2864
rect 244108 480 244136 2858
rect 245212 480 245240 16546
rect 246316 3330 246344 152866
rect 246408 143313 246436 219234
rect 246500 151298 246528 225626
rect 246592 217326 246620 229706
rect 246684 224954 246712 233174
rect 246776 226166 246804 239720
rect 246948 239420 247000 239426
rect 246948 239362 247000 239368
rect 246856 238808 246908 238814
rect 246856 238750 246908 238756
rect 246868 238542 246896 238750
rect 246856 238536 246908 238542
rect 246856 238478 246908 238484
rect 246856 234796 246908 234802
rect 246856 234738 246908 234744
rect 246764 226160 246816 226166
rect 246764 226102 246816 226108
rect 246868 226098 246896 234738
rect 246960 230178 246988 239362
rect 247052 239358 247080 239720
rect 247190 239680 247218 240108
rect 247282 239816 247310 240108
rect 247374 239970 247402 240108
rect 247362 239964 247414 239970
rect 247362 239906 247414 239912
rect 247466 239816 247494 240108
rect 247558 239873 247586 240108
rect 247650 239902 247678 240108
rect 247742 239970 247770 240108
rect 247834 239970 247862 240108
rect 247926 239970 247954 240108
rect 247730 239964 247782 239970
rect 247730 239906 247782 239912
rect 247822 239964 247874 239970
rect 247822 239906 247874 239912
rect 247914 239964 247966 239970
rect 247914 239906 247966 239912
rect 248018 239902 248046 240108
rect 248110 239902 248138 240108
rect 247638 239896 247690 239902
rect 247282 239788 247356 239816
rect 247144 239652 247218 239680
rect 247040 239352 247092 239358
rect 247040 239294 247092 239300
rect 246948 230172 247000 230178
rect 246948 230114 247000 230120
rect 246856 226092 246908 226098
rect 246856 226034 246908 226040
rect 246856 225888 246908 225894
rect 246856 225830 246908 225836
rect 246684 224926 246804 224954
rect 246776 219162 246804 224926
rect 246764 219156 246816 219162
rect 246764 219098 246816 219104
rect 246580 217320 246632 217326
rect 246580 217262 246632 217268
rect 246592 157146 246620 217262
rect 246776 171154 246804 219098
rect 246764 171148 246816 171154
rect 246764 171090 246816 171096
rect 246776 161474 246804 171090
rect 246684 161446 246804 161474
rect 246580 157140 246632 157146
rect 246580 157082 246632 157088
rect 246488 151292 246540 151298
rect 246488 151234 246540 151240
rect 246684 145926 246712 161446
rect 246672 145920 246724 145926
rect 246672 145862 246724 145868
rect 246394 143304 246450 143313
rect 246394 143239 246450 143248
rect 246868 140554 246896 225830
rect 246856 140548 246908 140554
rect 246856 140490 246908 140496
rect 246960 133346 246988 230114
rect 247144 215966 247172 239652
rect 247328 239465 247356 239788
rect 247420 239788 247494 239816
rect 247544 239864 247600 239873
rect 247638 239838 247690 239844
rect 248006 239896 248058 239902
rect 248006 239838 248058 239844
rect 248098 239896 248150 239902
rect 248098 239838 248150 239844
rect 247544 239799 247600 239808
rect 248202 239816 248230 240108
rect 248294 239970 248322 240108
rect 248282 239964 248334 239970
rect 248282 239906 248334 239912
rect 248386 239816 248414 240108
rect 248478 239970 248506 240108
rect 248466 239964 248518 239970
rect 248466 239906 248518 239912
rect 248570 239850 248598 240108
rect 248662 239873 248690 240108
rect 248524 239822 248598 239850
rect 248648 239864 248704 239873
rect 248202 239788 248276 239816
rect 248386 239788 248460 239816
rect 247314 239456 247370 239465
rect 247314 239391 247370 239400
rect 247420 238388 247448 239788
rect 247914 239760 247966 239766
rect 247966 239720 248092 239748
rect 247914 239702 247966 239708
rect 247960 239624 248012 239630
rect 247960 239566 248012 239572
rect 247500 239556 247552 239562
rect 247500 239498 247552 239504
rect 247684 239556 247736 239562
rect 247684 239498 247736 239504
rect 247868 239556 247920 239562
rect 247868 239498 247920 239504
rect 247328 238360 247448 238388
rect 247328 234734 247356 238360
rect 247512 236858 247540 239498
rect 247420 236830 247540 236858
rect 247316 234728 247368 234734
rect 247316 234670 247368 234676
rect 247420 231538 247448 236830
rect 247696 236722 247724 239498
rect 247880 239465 247908 239498
rect 247866 239456 247922 239465
rect 247866 239391 247922 239400
rect 247776 239148 247828 239154
rect 247776 239090 247828 239096
rect 247788 238882 247816 239090
rect 247776 238876 247828 238882
rect 247776 238818 247828 238824
rect 247880 237114 247908 239391
rect 247868 237108 247920 237114
rect 247868 237050 247920 237056
rect 247972 236994 248000 239566
rect 247512 236694 247724 236722
rect 247880 236966 248000 236994
rect 247408 231532 247460 231538
rect 247408 231474 247460 231480
rect 247420 230790 247448 231474
rect 247408 230784 247460 230790
rect 247408 230726 247460 230732
rect 247512 222902 247540 236694
rect 247880 236434 247908 236966
rect 247960 236632 248012 236638
rect 247960 236574 248012 236580
rect 247868 236428 247920 236434
rect 247868 236370 247920 236376
rect 247776 234728 247828 234734
rect 247776 234670 247828 234676
rect 247682 233880 247738 233889
rect 247682 233815 247738 233824
rect 247500 222896 247552 222902
rect 247500 222838 247552 222844
rect 247132 215960 247184 215966
rect 247132 215902 247184 215908
rect 247696 158506 247724 233815
rect 247788 226030 247816 234670
rect 247776 226024 247828 226030
rect 247776 225966 247828 225972
rect 247776 222896 247828 222902
rect 247776 222838 247828 222844
rect 247684 158500 247736 158506
rect 247684 158442 247736 158448
rect 247788 152998 247816 222838
rect 247868 215960 247920 215966
rect 247868 215902 247920 215908
rect 247776 152992 247828 152998
rect 247776 152934 247828 152940
rect 247880 151366 247908 215902
rect 247972 203658 248000 236574
rect 248064 232490 248092 239720
rect 248142 239728 248198 239737
rect 248142 239663 248144 239672
rect 248196 239663 248198 239672
rect 248144 239634 248196 239640
rect 248156 238134 248184 239634
rect 248144 238128 248196 238134
rect 248144 238070 248196 238076
rect 248248 237232 248276 239788
rect 248328 239692 248380 239698
rect 248328 239634 248380 239640
rect 248156 237204 248276 237232
rect 248052 232484 248104 232490
rect 248052 232426 248104 232432
rect 248156 231266 248184 237204
rect 248236 237108 248288 237114
rect 248236 237050 248288 237056
rect 248144 231260 248196 231266
rect 248144 231202 248196 231208
rect 248248 230874 248276 237050
rect 248340 236638 248368 239634
rect 248432 237250 248460 239788
rect 248420 237244 248472 237250
rect 248420 237186 248472 237192
rect 248524 236722 248552 239822
rect 248648 239799 248704 239808
rect 248754 239816 248782 240108
rect 248846 239970 248874 240108
rect 248834 239964 248886 239970
rect 248834 239906 248886 239912
rect 248938 239902 248966 240108
rect 249030 239902 249058 240108
rect 248926 239896 248978 239902
rect 248926 239838 248978 239844
rect 249018 239896 249070 239902
rect 249018 239838 249070 239844
rect 249122 239850 249150 240108
rect 249214 239970 249242 240108
rect 249202 239964 249254 239970
rect 249202 239906 249254 239912
rect 249122 239822 249196 239850
rect 248754 239788 248828 239816
rect 248604 239692 248656 239698
rect 248604 239634 248656 239640
rect 248432 236694 248552 236722
rect 248328 236632 248380 236638
rect 248328 236574 248380 236580
rect 248326 234288 248382 234297
rect 248326 234223 248382 234232
rect 248064 230846 248276 230874
rect 248064 229106 248092 230846
rect 248144 230784 248196 230790
rect 248144 230726 248196 230732
rect 248156 229242 248184 230726
rect 248340 229362 248368 234223
rect 248432 229770 248460 236694
rect 248616 235482 248644 239634
rect 248800 239544 248828 239788
rect 249064 239760 249116 239766
rect 248878 239728 248934 239737
rect 249064 239702 249116 239708
rect 248878 239663 248880 239672
rect 248932 239663 248934 239672
rect 248972 239692 249024 239698
rect 248880 239634 248932 239640
rect 248972 239634 249024 239640
rect 248800 239516 248920 239544
rect 248696 239488 248748 239494
rect 248696 239430 248748 239436
rect 248604 235476 248656 235482
rect 248604 235418 248656 235424
rect 248708 233234 248736 239430
rect 248788 239420 248840 239426
rect 248788 239362 248840 239368
rect 248800 236722 248828 239362
rect 248892 238338 248920 239516
rect 248984 238814 249012 239634
rect 249076 239426 249104 239702
rect 249064 239420 249116 239426
rect 249064 239362 249116 239368
rect 249168 238898 249196 239822
rect 249306 239816 249334 240108
rect 249398 239970 249426 240108
rect 249386 239964 249438 239970
rect 249386 239906 249438 239912
rect 249306 239788 249380 239816
rect 249352 239698 249380 239788
rect 249340 239692 249392 239698
rect 249490 239680 249518 240108
rect 249582 239902 249610 240108
rect 249674 239902 249702 240108
rect 249570 239896 249622 239902
rect 249570 239838 249622 239844
rect 249662 239896 249714 239902
rect 249766 239873 249794 240108
rect 249858 239902 249886 240108
rect 249950 239970 249978 240108
rect 249938 239964 249990 239970
rect 249938 239906 249990 239912
rect 249846 239896 249898 239902
rect 249662 239838 249714 239844
rect 249752 239864 249808 239873
rect 249846 239838 249898 239844
rect 250042 239816 250070 240108
rect 249752 239799 249808 239808
rect 249996 239788 250070 239816
rect 249800 239760 249852 239766
rect 249892 239760 249944 239766
rect 249800 239702 249852 239708
rect 249890 239728 249892 239737
rect 249944 239728 249946 239737
rect 249490 239652 249564 239680
rect 249340 239634 249392 239640
rect 249340 239556 249392 239562
rect 249340 239498 249392 239504
rect 249248 239420 249300 239426
rect 249248 239362 249300 239368
rect 249076 238870 249196 238898
rect 248972 238808 249024 238814
rect 248972 238750 249024 238756
rect 248880 238332 248932 238338
rect 248880 238274 248932 238280
rect 249076 237930 249104 238870
rect 249156 238808 249208 238814
rect 249156 238750 249208 238756
rect 249064 237924 249116 237930
rect 249064 237866 249116 237872
rect 248800 236694 248920 236722
rect 248786 236464 248842 236473
rect 248786 236399 248842 236408
rect 248524 233206 248736 233234
rect 248420 229764 248472 229770
rect 248420 229706 248472 229712
rect 248328 229356 248380 229362
rect 248328 229298 248380 229304
rect 248156 229214 248368 229242
rect 248064 229078 248276 229106
rect 247960 203652 248012 203658
rect 247960 203594 248012 203600
rect 247972 156874 248000 203594
rect 248248 175302 248276 229078
rect 248236 175296 248288 175302
rect 248236 175238 248288 175244
rect 248248 161474 248276 175238
rect 248064 161446 248276 161474
rect 247960 156868 248012 156874
rect 247960 156810 248012 156816
rect 247868 151360 247920 151366
rect 247868 151302 247920 151308
rect 248064 148782 248092 161446
rect 248052 148776 248104 148782
rect 248052 148718 248104 148724
rect 246948 133340 247000 133346
rect 246948 133282 247000 133288
rect 247040 132320 247092 132326
rect 247040 132262 247092 132268
rect 247052 131918 247080 132262
rect 248340 131918 248368 229214
rect 248524 220386 248552 233206
rect 248800 228585 248828 236399
rect 248786 228576 248842 228585
rect 248786 228511 248842 228520
rect 248892 227066 248920 236694
rect 248972 236632 249024 236638
rect 248972 236574 249024 236580
rect 248984 231402 249012 236574
rect 249168 234598 249196 238750
rect 249260 236978 249288 239362
rect 249352 238134 249380 239498
rect 249536 239465 249564 239652
rect 249708 239556 249760 239562
rect 249708 239498 249760 239504
rect 249616 239488 249668 239494
rect 249522 239456 249578 239465
rect 249616 239430 249668 239436
rect 249522 239391 249578 239400
rect 249340 238128 249392 238134
rect 249340 238070 249392 238076
rect 249248 236972 249300 236978
rect 249248 236914 249300 236920
rect 249156 234592 249208 234598
rect 249156 234534 249208 234540
rect 249536 233234 249564 239391
rect 249444 233206 249564 233234
rect 248972 231396 249024 231402
rect 248972 231338 249024 231344
rect 249340 230172 249392 230178
rect 249340 230114 249392 230120
rect 249352 229634 249380 230114
rect 249340 229628 249392 229634
rect 249340 229570 249392 229576
rect 248970 228576 249026 228585
rect 248970 228511 249026 228520
rect 248984 227390 249012 228511
rect 249338 228440 249394 228449
rect 249338 228375 249394 228384
rect 248972 227384 249024 227390
rect 248972 227326 249024 227332
rect 249352 227254 249380 228375
rect 249340 227248 249392 227254
rect 249340 227190 249392 227196
rect 248616 227038 248920 227066
rect 248616 222154 248644 227038
rect 248696 226772 248748 226778
rect 248696 226714 248748 226720
rect 248708 224806 248736 226714
rect 249444 224954 249472 233206
rect 249524 229764 249576 229770
rect 249524 229706 249576 229712
rect 249076 224926 249472 224954
rect 248696 224800 248748 224806
rect 248696 224742 248748 224748
rect 248604 222148 248656 222154
rect 248604 222090 248656 222096
rect 248512 220380 248564 220386
rect 248512 220322 248564 220328
rect 249076 141778 249104 224926
rect 249432 224800 249484 224806
rect 249432 224742 249484 224748
rect 249340 222148 249392 222154
rect 249340 222090 249392 222096
rect 249352 221474 249380 222090
rect 249340 221468 249392 221474
rect 249340 221410 249392 221416
rect 249156 220380 249208 220386
rect 249156 220322 249208 220328
rect 249168 220114 249196 220322
rect 249156 220108 249208 220114
rect 249156 220050 249208 220056
rect 249168 148442 249196 220050
rect 249248 218068 249300 218074
rect 249248 218010 249300 218016
rect 249260 148578 249288 218010
rect 249352 157962 249380 221410
rect 249444 161129 249472 224742
rect 249536 218754 249564 229706
rect 249628 226778 249656 239430
rect 249720 236638 249748 239498
rect 249708 236632 249760 236638
rect 249708 236574 249760 236580
rect 249812 232966 249840 239702
rect 249890 239663 249946 239672
rect 249890 236736 249946 236745
rect 249890 236671 249946 236680
rect 249800 232960 249852 232966
rect 249800 232902 249852 232908
rect 249812 231860 249840 232902
rect 249720 231832 249840 231860
rect 249616 226772 249668 226778
rect 249616 226714 249668 226720
rect 249720 224954 249748 231832
rect 249800 230444 249852 230450
rect 249800 230386 249852 230392
rect 249812 229702 249840 230386
rect 249800 229696 249852 229702
rect 249800 229638 249852 229644
rect 249628 224926 249748 224954
rect 249524 218748 249576 218754
rect 249524 218690 249576 218696
rect 249536 218074 249564 218690
rect 249524 218068 249576 218074
rect 249524 218010 249576 218016
rect 249430 161120 249486 161129
rect 249430 161055 249486 161064
rect 249340 157956 249392 157962
rect 249340 157898 249392 157904
rect 249248 148572 249300 148578
rect 249248 148514 249300 148520
rect 249156 148436 249208 148442
rect 249156 148378 249208 148384
rect 249432 148368 249484 148374
rect 249432 148310 249484 148316
rect 249444 147422 249472 148310
rect 249432 147416 249484 147422
rect 249432 147358 249484 147364
rect 249064 141772 249116 141778
rect 249064 141714 249116 141720
rect 249628 136474 249656 224926
rect 249904 219434 249932 236671
rect 249812 219406 249932 219434
rect 249812 204950 249840 219406
rect 249996 219298 250024 239788
rect 250134 239748 250162 240108
rect 250088 239720 250162 239748
rect 250226 239748 250254 240108
rect 250318 239907 250346 240108
rect 250304 239898 250360 239907
rect 250304 239833 250360 239842
rect 250410 239748 250438 240108
rect 250226 239720 250300 239748
rect 250088 231985 250116 239720
rect 250272 239680 250300 239720
rect 250180 239652 250300 239680
rect 250364 239720 250438 239748
rect 250180 239426 250208 239652
rect 250168 239420 250220 239426
rect 250168 239362 250220 239368
rect 250168 238876 250220 238882
rect 250168 238818 250220 238824
rect 250180 238542 250208 238818
rect 250168 238536 250220 238542
rect 250168 238478 250220 238484
rect 250364 233234 250392 239720
rect 250502 239680 250530 240108
rect 250594 239970 250622 240108
rect 250686 239970 250714 240108
rect 250582 239964 250634 239970
rect 250582 239906 250634 239912
rect 250674 239964 250726 239970
rect 250674 239906 250726 239912
rect 250778 239850 250806 240108
rect 250180 233206 250392 233234
rect 250456 239652 250530 239680
rect 250640 239822 250806 239850
rect 250180 232830 250208 233206
rect 250168 232824 250220 232830
rect 250168 232766 250220 232772
rect 250074 231976 250130 231985
rect 250074 231911 250130 231920
rect 250456 230450 250484 239652
rect 250536 239556 250588 239562
rect 250536 239498 250588 239504
rect 250548 234326 250576 239498
rect 250536 234320 250588 234326
rect 250536 234262 250588 234268
rect 250444 230444 250496 230450
rect 250444 230386 250496 230392
rect 250534 222184 250590 222193
rect 250534 222119 250590 222128
rect 249984 219292 250036 219298
rect 249984 219234 250036 219240
rect 249800 204944 249852 204950
rect 249800 204886 249852 204892
rect 250444 204944 250496 204950
rect 250444 204886 250496 204892
rect 250456 157486 250484 204886
rect 250444 157480 250496 157486
rect 250444 157422 250496 157428
rect 250444 153876 250496 153882
rect 250444 153818 250496 153824
rect 249708 147416 249760 147422
rect 249708 147358 249760 147364
rect 249616 136468 249668 136474
rect 249616 136410 249668 136416
rect 249628 136066 249656 136410
rect 249616 136060 249668 136066
rect 249616 136002 249668 136008
rect 247040 131912 247092 131918
rect 247040 131854 247092 131860
rect 248328 131912 248380 131918
rect 248328 131854 248380 131860
rect 247682 112432 247738 112441
rect 247682 112367 247738 112376
rect 246396 4140 246448 4146
rect 246396 4082 246448 4088
rect 246304 3324 246356 3330
rect 246304 3266 246356 3272
rect 246408 480 246436 4082
rect 247592 2984 247644 2990
rect 247592 2926 247644 2932
rect 247604 480 247632 2926
rect 247696 2922 247724 112367
rect 249720 3194 249748 147358
rect 250456 4146 250484 153818
rect 250548 149977 250576 222119
rect 250640 213246 250668 239822
rect 250720 239760 250772 239766
rect 250720 239702 250772 239708
rect 250732 238649 250760 239702
rect 250870 239680 250898 240108
rect 250962 239748 250990 240108
rect 251054 239902 251082 240108
rect 251042 239896 251094 239902
rect 251042 239838 251094 239844
rect 251146 239816 251174 240108
rect 251238 239970 251266 240108
rect 251330 239970 251358 240108
rect 251422 239970 251450 240108
rect 251514 239970 251542 240108
rect 251226 239964 251278 239970
rect 251226 239906 251278 239912
rect 251318 239964 251370 239970
rect 251318 239906 251370 239912
rect 251410 239964 251462 239970
rect 251410 239906 251462 239912
rect 251502 239964 251554 239970
rect 251502 239906 251554 239912
rect 251606 239850 251634 240108
rect 251698 239970 251726 240108
rect 251790 239970 251818 240108
rect 251882 239970 251910 240108
rect 251686 239964 251738 239970
rect 251686 239906 251738 239912
rect 251778 239964 251830 239970
rect 251778 239906 251830 239912
rect 251870 239964 251922 239970
rect 251870 239906 251922 239912
rect 251822 239864 251878 239873
rect 251606 239822 251680 239850
rect 251146 239788 251220 239816
rect 250962 239737 251036 239748
rect 250962 239728 251050 239737
rect 250962 239720 250994 239728
rect 250870 239652 250944 239680
rect 250994 239663 251050 239672
rect 250812 239420 250864 239426
rect 250812 239362 250864 239368
rect 250718 238640 250774 238649
rect 250718 238575 250774 238584
rect 250824 237969 250852 239362
rect 250810 237960 250866 237969
rect 250810 237895 250866 237904
rect 250916 233986 250944 239652
rect 250996 239624 251048 239630
rect 251192 239612 251220 239788
rect 251548 239760 251600 239766
rect 251454 239728 251510 239737
rect 251548 239702 251600 239708
rect 251454 239663 251510 239672
rect 250996 239566 251048 239572
rect 251100 239584 251220 239612
rect 251272 239624 251324 239630
rect 251008 238785 251036 239566
rect 250994 238776 251050 238785
rect 250994 238711 251050 238720
rect 250996 238536 251048 238542
rect 250996 238478 251048 238484
rect 250904 233980 250956 233986
rect 250904 233922 250956 233928
rect 250902 232792 250958 232801
rect 250902 232727 250958 232736
rect 250916 231985 250944 232727
rect 250902 231976 250958 231985
rect 250902 231911 250958 231920
rect 250628 213240 250680 213246
rect 250628 213182 250680 213188
rect 250534 149968 250590 149977
rect 250534 149903 250590 149912
rect 250640 146742 250668 213182
rect 250628 146736 250680 146742
rect 250628 146678 250680 146684
rect 250916 145994 250944 231911
rect 251008 231674 251036 238478
rect 251100 233714 251128 239584
rect 251272 239566 251324 239572
rect 251180 239488 251232 239494
rect 251180 239430 251232 239436
rect 251192 238542 251220 239430
rect 251180 238536 251232 238542
rect 251180 238478 251232 238484
rect 251180 237312 251232 237318
rect 251180 237254 251232 237260
rect 251088 233708 251140 233714
rect 251088 233650 251140 233656
rect 251088 233164 251140 233170
rect 251088 233106 251140 233112
rect 251100 232830 251128 233106
rect 251088 232824 251140 232830
rect 251088 232766 251140 232772
rect 250996 231668 251048 231674
rect 250996 231610 251048 231616
rect 250904 145988 250956 145994
rect 250904 145930 250956 145936
rect 250916 145654 250944 145930
rect 250904 145648 250956 145654
rect 250904 145590 250956 145596
rect 251008 135250 251036 231610
rect 250996 135244 251048 135250
rect 250996 135186 251048 135192
rect 251008 134638 251036 135186
rect 250996 134632 251048 134638
rect 250996 134574 251048 134580
rect 251100 125526 251128 232766
rect 251192 214849 251220 237254
rect 251284 229770 251312 239566
rect 251468 237998 251496 239663
rect 251560 239442 251588 239702
rect 251652 239562 251680 239822
rect 251732 239828 251784 239834
rect 251974 239850 252002 240108
rect 252066 239902 252094 240108
rect 251822 239799 251878 239808
rect 251928 239822 252002 239850
rect 252054 239896 252106 239902
rect 252054 239838 252106 239844
rect 251732 239770 251784 239776
rect 251640 239556 251692 239562
rect 251640 239498 251692 239504
rect 251560 239414 251680 239442
rect 251548 239352 251600 239358
rect 251548 239294 251600 239300
rect 251456 237992 251508 237998
rect 251456 237934 251508 237940
rect 251456 237856 251508 237862
rect 251456 237798 251508 237804
rect 251468 237318 251496 237798
rect 251456 237312 251508 237318
rect 251456 237254 251508 237260
rect 251560 237046 251588 239294
rect 251652 237862 251680 239414
rect 251744 238746 251772 239770
rect 251836 239766 251864 239799
rect 251824 239760 251876 239766
rect 251928 239737 251956 239822
rect 252158 239816 252186 240108
rect 252250 239970 252278 240108
rect 252238 239964 252290 239970
rect 252238 239906 252290 239912
rect 252342 239850 252370 240108
rect 252434 239902 252462 240108
rect 252296 239822 252370 239850
rect 252422 239896 252474 239902
rect 252422 239838 252474 239844
rect 252158 239788 252232 239816
rect 251824 239702 251876 239708
rect 251914 239728 251970 239737
rect 251914 239663 251970 239672
rect 251916 239624 251968 239630
rect 251968 239584 252140 239612
rect 251916 239566 251968 239572
rect 251824 239556 251876 239562
rect 251824 239498 251876 239504
rect 251732 238740 251784 238746
rect 251732 238682 251784 238688
rect 251732 238060 251784 238066
rect 251732 238002 251784 238008
rect 251640 237856 251692 237862
rect 251640 237798 251692 237804
rect 251548 237040 251600 237046
rect 251548 236982 251600 236988
rect 251744 236978 251772 238002
rect 251732 236972 251784 236978
rect 251732 236914 251784 236920
rect 251272 229764 251324 229770
rect 251272 229706 251324 229712
rect 251836 226166 251864 239498
rect 252008 239488 252060 239494
rect 252008 239430 252060 239436
rect 252020 235210 252048 239430
rect 252112 236473 252140 239584
rect 252098 236464 252154 236473
rect 252098 236399 252154 236408
rect 252008 235204 252060 235210
rect 252008 235146 252060 235152
rect 252204 233234 252232 239788
rect 252112 233206 252232 233234
rect 252112 227594 252140 233206
rect 252296 232626 252324 239822
rect 252376 239760 252428 239766
rect 252526 239748 252554 240108
rect 252618 239907 252646 240108
rect 252710 239970 252738 240108
rect 252698 239964 252750 239970
rect 252604 239898 252660 239907
rect 252698 239906 252750 239912
rect 252604 239833 252660 239842
rect 252802 239816 252830 240108
rect 252894 239970 252922 240108
rect 252986 239970 253014 240108
rect 252882 239964 252934 239970
rect 252882 239906 252934 239912
rect 252974 239964 253026 239970
rect 252974 239906 253026 239912
rect 253078 239850 253106 240108
rect 252376 239702 252428 239708
rect 252480 239720 252554 239748
rect 252756 239788 252830 239816
rect 253032 239822 253106 239850
rect 252756 239737 252784 239788
rect 252742 239728 252798 239737
rect 252284 232620 252336 232626
rect 252284 232562 252336 232568
rect 252388 231854 252416 239702
rect 252480 232558 252508 239720
rect 252742 239663 252798 239672
rect 252836 239692 252888 239698
rect 252836 239634 252888 239640
rect 252744 239624 252796 239630
rect 252744 239566 252796 239572
rect 252560 239556 252612 239562
rect 252560 239498 252612 239504
rect 252572 239465 252600 239498
rect 252558 239456 252614 239465
rect 252558 239391 252614 239400
rect 252560 239352 252612 239358
rect 252560 239294 252612 239300
rect 252572 235940 252600 239294
rect 252572 235912 252692 235940
rect 252468 232552 252520 232558
rect 252468 232494 252520 232500
rect 252204 231826 252416 231854
rect 252560 231872 252612 231878
rect 252100 227588 252152 227594
rect 252100 227530 252152 227536
rect 251824 226160 251876 226166
rect 251824 226102 251876 226108
rect 251272 224188 251324 224194
rect 251272 224130 251324 224136
rect 251178 214840 251234 214849
rect 251178 214775 251234 214784
rect 251284 150958 251312 224130
rect 251836 158710 251864 226102
rect 252112 224954 252140 227530
rect 251928 224926 252140 224954
rect 251824 158704 251876 158710
rect 251824 158646 251876 158652
rect 251272 150952 251324 150958
rect 251272 150894 251324 150900
rect 251284 150482 251312 150894
rect 251272 150476 251324 150482
rect 251272 150418 251324 150424
rect 251824 150476 251876 150482
rect 251824 150418 251876 150424
rect 251088 125520 251140 125526
rect 251088 125462 251140 125468
rect 251100 124982 251128 125462
rect 251088 124976 251140 124982
rect 251088 124918 251140 124924
rect 251270 95976 251326 95985
rect 251270 95911 251326 95920
rect 251284 16574 251312 95911
rect 251284 16546 251772 16574
rect 250444 4140 250496 4146
rect 250444 4082 250496 4088
rect 249984 4004 250036 4010
rect 249984 3946 250036 3952
rect 249708 3188 249760 3194
rect 249708 3130 249760 3136
rect 247684 2916 247736 2922
rect 247684 2858 247736 2864
rect 248788 2916 248840 2922
rect 248788 2858 248840 2864
rect 248800 480 248828 2858
rect 249996 480 250024 3946
rect 251744 3482 251772 16546
rect 251836 3670 251864 150418
rect 251928 148510 251956 224926
rect 252008 224800 252060 224806
rect 252008 224742 252060 224748
rect 252020 158302 252048 224742
rect 252204 222018 252232 231826
rect 252560 231814 252612 231820
rect 252572 231441 252600 231814
rect 252558 231432 252614 231441
rect 252558 231367 252614 231376
rect 252466 230072 252522 230081
rect 252466 230007 252522 230016
rect 252376 229764 252428 229770
rect 252376 229706 252428 229712
rect 252388 224806 252416 229706
rect 252376 224800 252428 224806
rect 252376 224742 252428 224748
rect 252192 222012 252244 222018
rect 252192 221954 252244 221960
rect 252204 219434 252232 221954
rect 252112 219406 252232 219434
rect 252008 158296 252060 158302
rect 252008 158238 252060 158244
rect 252112 158234 252140 219406
rect 252100 158228 252152 158234
rect 252100 158170 252152 158176
rect 251916 148504 251968 148510
rect 251916 148446 251968 148452
rect 252480 124166 252508 230007
rect 252560 229764 252612 229770
rect 252560 229706 252612 229712
rect 252572 214606 252600 229706
rect 252664 222086 252692 235912
rect 252756 222154 252784 239566
rect 252848 238490 252876 239634
rect 252928 239488 252980 239494
rect 253032 239465 253060 239822
rect 253170 239748 253198 240108
rect 253262 239970 253290 240108
rect 253250 239964 253302 239970
rect 253250 239906 253302 239912
rect 253354 239850 253382 240108
rect 253308 239822 253382 239850
rect 253308 239748 253336 239822
rect 253124 239720 253198 239748
rect 253262 239720 253336 239748
rect 253446 239748 253474 240108
rect 253538 239902 253566 240108
rect 253630 239902 253658 240108
rect 253526 239896 253578 239902
rect 253526 239838 253578 239844
rect 253618 239896 253670 239902
rect 253618 239838 253670 239844
rect 253572 239760 253624 239766
rect 253446 239720 253520 239748
rect 252928 239430 252980 239436
rect 253018 239456 253074 239465
rect 252940 238678 252968 239430
rect 253018 239391 253074 239400
rect 252928 238672 252980 238678
rect 252928 238614 252980 238620
rect 252848 238462 252968 238490
rect 252836 237992 252888 237998
rect 252836 237934 252888 237940
rect 252848 236638 252876 237934
rect 252836 236632 252888 236638
rect 252940 236609 252968 238462
rect 252836 236574 252888 236580
rect 252926 236600 252982 236609
rect 252926 236535 252982 236544
rect 252940 230858 252968 236535
rect 253032 235249 253060 239391
rect 253124 236745 253152 239720
rect 253262 239578 253290 239720
rect 253388 239624 253440 239630
rect 253262 239550 253336 239578
rect 253388 239566 253440 239572
rect 253308 238105 253336 239550
rect 253294 238096 253350 238105
rect 253294 238031 253350 238040
rect 253400 237289 253428 239566
rect 253386 237280 253442 237289
rect 253386 237215 253442 237224
rect 253110 236736 253166 236745
rect 253110 236671 253166 236680
rect 253492 236570 253520 239720
rect 253722 239748 253750 240108
rect 253572 239702 253624 239708
rect 253676 239720 253750 239748
rect 253584 237454 253612 239702
rect 253572 237448 253624 237454
rect 253572 237390 253624 237396
rect 253572 237312 253624 237318
rect 253572 237254 253624 237260
rect 253584 237114 253612 237254
rect 253572 237108 253624 237114
rect 253572 237050 253624 237056
rect 253480 236564 253532 236570
rect 253480 236506 253532 236512
rect 253676 235958 253704 239720
rect 253814 239680 253842 240108
rect 253906 239970 253934 240108
rect 253894 239964 253946 239970
rect 253894 239906 253946 239912
rect 253998 239850 254026 240108
rect 253768 239652 253842 239680
rect 253952 239822 254026 239850
rect 253112 235952 253164 235958
rect 253112 235894 253164 235900
rect 253664 235952 253716 235958
rect 253664 235894 253716 235900
rect 253018 235240 253074 235249
rect 253018 235175 253074 235184
rect 252928 230852 252980 230858
rect 252928 230794 252980 230800
rect 253124 222834 253152 235894
rect 253662 235784 253718 235793
rect 253662 235719 253718 235728
rect 253480 235340 253532 235346
rect 253480 235282 253532 235288
rect 253492 233238 253520 235282
rect 253572 233504 253624 233510
rect 253572 233446 253624 233452
rect 253480 233232 253532 233238
rect 253480 233174 253532 233180
rect 253204 232960 253256 232966
rect 253204 232902 253256 232908
rect 253216 232830 253244 232902
rect 253204 232824 253256 232830
rect 253204 232766 253256 232772
rect 253584 231334 253612 233446
rect 253572 231328 253624 231334
rect 253572 231270 253624 231276
rect 253584 229634 253612 231270
rect 253572 229628 253624 229634
rect 253572 229570 253624 229576
rect 253676 224954 253704 235719
rect 253768 229770 253796 239652
rect 253848 239556 253900 239562
rect 253848 239498 253900 239504
rect 253860 239465 253888 239498
rect 253846 239456 253902 239465
rect 253846 239391 253902 239400
rect 253848 239352 253900 239358
rect 253848 239294 253900 239300
rect 253860 235346 253888 239294
rect 253848 235340 253900 235346
rect 253848 235282 253900 235288
rect 253952 235090 253980 239822
rect 254090 239748 254118 240108
rect 254182 239902 254210 240108
rect 254274 239970 254302 240108
rect 254262 239964 254314 239970
rect 254262 239906 254314 239912
rect 254170 239896 254222 239902
rect 254366 239850 254394 240108
rect 254170 239838 254222 239844
rect 254320 239822 254394 239850
rect 254458 239850 254486 240108
rect 254550 239970 254578 240108
rect 254538 239964 254590 239970
rect 254538 239906 254590 239912
rect 254458 239822 254532 239850
rect 254090 239720 254164 239748
rect 254032 239420 254084 239426
rect 254032 239362 254084 239368
rect 253860 235062 253980 235090
rect 253860 233510 253888 235062
rect 254044 234938 254072 239362
rect 254032 234932 254084 234938
rect 254032 234874 254084 234880
rect 253848 233504 253900 233510
rect 253848 233446 253900 233452
rect 253848 233232 253900 233238
rect 253848 233174 253900 233180
rect 254032 233232 254084 233238
rect 254032 233174 254084 233180
rect 253860 232966 253888 233174
rect 253848 232960 253900 232966
rect 253848 232902 253900 232908
rect 253756 229764 253808 229770
rect 253756 229706 253808 229712
rect 253756 229628 253808 229634
rect 253756 229570 253808 229576
rect 253400 224926 253704 224954
rect 253112 222828 253164 222834
rect 253112 222770 253164 222776
rect 252744 222148 252796 222154
rect 252744 222090 252796 222096
rect 253204 222148 253256 222154
rect 253204 222090 253256 222096
rect 252652 222080 252704 222086
rect 252652 222022 252704 222028
rect 253216 221746 253244 222090
rect 253296 221944 253348 221950
rect 253296 221886 253348 221892
rect 253204 221740 253256 221746
rect 253204 221682 253256 221688
rect 253110 218104 253166 218113
rect 253110 218039 253166 218048
rect 252560 214600 252612 214606
rect 253124 214577 253152 218039
rect 252560 214542 252612 214548
rect 253110 214568 253166 214577
rect 253110 214503 253166 214512
rect 252560 213308 252612 213314
rect 252560 213250 252612 213256
rect 252572 155514 252600 213250
rect 253216 158166 253244 221682
rect 253204 158160 253256 158166
rect 253204 158102 253256 158108
rect 252560 155508 252612 155514
rect 252560 155450 252612 155456
rect 253204 155508 253256 155514
rect 253204 155450 253256 155456
rect 252572 154970 252600 155450
rect 252560 154964 252612 154970
rect 252560 154906 252612 154912
rect 252468 124160 252520 124166
rect 252468 124102 252520 124108
rect 252480 123554 252508 124102
rect 252468 123548 252520 123554
rect 252468 123490 252520 123496
rect 253112 3936 253164 3942
rect 253112 3878 253164 3884
rect 253216 3890 253244 155450
rect 253308 151337 253336 221886
rect 253294 151328 253350 151337
rect 253294 151263 253350 151272
rect 253296 146940 253348 146946
rect 253296 146882 253348 146888
rect 253308 4010 253336 146882
rect 253400 117298 253428 224926
rect 253480 222080 253532 222086
rect 253480 222022 253532 222028
rect 253492 221814 253520 222022
rect 253480 221808 253532 221814
rect 253480 221750 253532 221756
rect 253492 147150 253520 221750
rect 253572 214600 253624 214606
rect 253572 214542 253624 214548
rect 253480 147144 253532 147150
rect 253480 147086 253532 147092
rect 253584 146810 253612 214542
rect 253768 147218 253796 229570
rect 253756 147212 253808 147218
rect 253756 147154 253808 147160
rect 253572 146804 253624 146810
rect 253572 146746 253624 146752
rect 253860 126818 253888 232902
rect 254044 232558 254072 233174
rect 254032 232552 254084 232558
rect 254032 232494 254084 232500
rect 254032 229764 254084 229770
rect 254032 229706 254084 229712
rect 253938 223136 253994 223145
rect 253938 223071 253994 223080
rect 253952 221882 253980 223071
rect 253940 221876 253992 221882
rect 253940 221818 253992 221824
rect 254044 221406 254072 229706
rect 254136 222154 254164 239720
rect 254320 239578 254348 239822
rect 254400 239760 254452 239766
rect 254400 239702 254452 239708
rect 254228 239550 254348 239578
rect 254228 223242 254256 239550
rect 254308 239488 254360 239494
rect 254308 239430 254360 239436
rect 254320 231854 254348 239430
rect 254412 237114 254440 239702
rect 254400 237108 254452 237114
rect 254400 237050 254452 237056
rect 254412 236910 254440 237050
rect 254400 236904 254452 236910
rect 254400 236846 254452 236852
rect 254504 232393 254532 239822
rect 254642 239816 254670 240108
rect 254734 239873 254762 240108
rect 254596 239788 254670 239816
rect 254720 239864 254776 239873
rect 254720 239799 254776 239808
rect 254490 232384 254546 232393
rect 254490 232319 254546 232328
rect 254320 231826 254440 231854
rect 254308 229696 254360 229702
rect 254308 229638 254360 229644
rect 254216 223236 254268 223242
rect 254216 223178 254268 223184
rect 254320 223106 254348 229638
rect 254412 223145 254440 231826
rect 254596 229702 254624 239788
rect 254826 239748 254854 240108
rect 254780 239720 254854 239748
rect 254918 239748 254946 240108
rect 255010 239902 255038 240108
rect 254998 239896 255050 239902
rect 254998 239838 255050 239844
rect 255102 239850 255130 240108
rect 255194 239970 255222 240108
rect 255182 239964 255234 239970
rect 255182 239906 255234 239912
rect 255102 239834 255176 239850
rect 255102 239828 255188 239834
rect 255102 239822 255136 239828
rect 255136 239770 255188 239776
rect 255286 239748 255314 240108
rect 254918 239720 254992 239748
rect 254676 239692 254728 239698
rect 254676 239634 254728 239640
rect 254688 237998 254716 239634
rect 254676 237992 254728 237998
rect 254676 237934 254728 237940
rect 254676 237448 254728 237454
rect 254676 237390 254728 237396
rect 254584 229696 254636 229702
rect 254584 229638 254636 229644
rect 254688 224954 254716 237390
rect 254780 235142 254808 239720
rect 254964 239442 254992 239720
rect 255134 239728 255190 239737
rect 255134 239663 255190 239672
rect 255240 239720 255314 239748
rect 255378 239748 255406 240108
rect 255470 239970 255498 240108
rect 255458 239964 255510 239970
rect 255458 239906 255510 239912
rect 255562 239816 255590 240108
rect 255654 239902 255682 240108
rect 255642 239896 255694 239902
rect 255642 239838 255694 239844
rect 255516 239788 255590 239816
rect 255746 239816 255774 240108
rect 255838 239970 255866 240108
rect 255826 239964 255878 239970
rect 255826 239906 255878 239912
rect 255930 239816 255958 240108
rect 256022 239902 256050 240108
rect 256114 239907 256142 240108
rect 256010 239896 256062 239902
rect 256010 239838 256062 239844
rect 256100 239898 256156 239907
rect 256100 239833 256156 239842
rect 255746 239788 255820 239816
rect 255378 239720 255452 239748
rect 254872 239414 254992 239442
rect 254872 237833 254900 239414
rect 254952 239352 255004 239358
rect 254952 239294 255004 239300
rect 254858 237824 254914 237833
rect 254858 237759 254914 237768
rect 254768 235136 254820 235142
rect 254768 235078 254820 235084
rect 254964 229770 254992 239294
rect 255148 238882 255176 239663
rect 255136 238876 255188 238882
rect 255136 238818 255188 238824
rect 255240 238728 255268 239720
rect 255320 239624 255372 239630
rect 255320 239566 255372 239572
rect 255056 238700 255268 238728
rect 254952 229764 255004 229770
rect 254952 229706 255004 229712
rect 254688 224926 254992 224954
rect 254860 223236 254912 223242
rect 254860 223178 254912 223184
rect 254398 223136 254454 223145
rect 254308 223100 254360 223106
rect 254398 223071 254454 223080
rect 254308 223042 254360 223048
rect 254124 222148 254176 222154
rect 254124 222090 254176 222096
rect 254032 221400 254084 221406
rect 254032 221342 254084 221348
rect 254320 219434 254348 223042
rect 254676 222148 254728 222154
rect 254676 222090 254728 222096
rect 254688 221882 254716 222090
rect 254768 222012 254820 222018
rect 254768 221954 254820 221960
rect 254676 221876 254728 221882
rect 254676 221818 254728 221824
rect 254320 219406 254624 219434
rect 254596 147082 254624 219406
rect 254688 147354 254716 221818
rect 254780 221406 254808 221954
rect 254768 221400 254820 221406
rect 254768 221342 254820 221348
rect 254780 151473 254808 221342
rect 254872 161090 254900 223178
rect 254964 222154 254992 224926
rect 254952 222148 255004 222154
rect 254952 222090 255004 222096
rect 254964 221950 254992 222090
rect 254952 221944 255004 221950
rect 254952 221886 255004 221892
rect 255056 219201 255084 238700
rect 255134 238640 255190 238649
rect 255134 238575 255190 238584
rect 255228 238604 255280 238610
rect 255148 238542 255176 238575
rect 255228 238546 255280 238552
rect 255136 238536 255188 238542
rect 255136 238478 255188 238484
rect 255148 230654 255176 238478
rect 255240 238270 255268 238546
rect 255228 238264 255280 238270
rect 255228 238206 255280 238212
rect 255332 236026 255360 239566
rect 255424 238066 255452 239720
rect 255412 238060 255464 238066
rect 255412 238002 255464 238008
rect 255410 237960 255466 237969
rect 255410 237895 255466 237904
rect 255320 236020 255372 236026
rect 255320 235962 255372 235968
rect 255228 234932 255280 234938
rect 255228 234874 255280 234880
rect 255240 233209 255268 234874
rect 255226 233200 255282 233209
rect 255226 233135 255282 233144
rect 255136 230648 255188 230654
rect 255136 230590 255188 230596
rect 255042 219192 255098 219201
rect 255042 219127 255098 219136
rect 255056 214985 255084 219127
rect 255042 214976 255098 214985
rect 255042 214911 255098 214920
rect 254860 161084 254912 161090
rect 254860 161026 254912 161032
rect 254766 151464 254822 151473
rect 254766 151399 254822 151408
rect 254676 147348 254728 147354
rect 254676 147290 254728 147296
rect 254584 147076 254636 147082
rect 254584 147018 254636 147024
rect 255240 131102 255268 233135
rect 255424 157690 255452 237895
rect 255516 230790 255544 239788
rect 255596 239692 255648 239698
rect 255596 239634 255648 239640
rect 255688 239692 255740 239698
rect 255688 239634 255740 239640
rect 255608 237833 255636 239634
rect 255700 239193 255728 239634
rect 255686 239184 255742 239193
rect 255686 239119 255742 239128
rect 255688 238876 255740 238882
rect 255688 238818 255740 238824
rect 255594 237824 255650 237833
rect 255594 237759 255650 237768
rect 255608 235278 255636 237759
rect 255700 236842 255728 238818
rect 255688 236836 255740 236842
rect 255688 236778 255740 236784
rect 255792 236745 255820 239788
rect 255884 239788 255958 239816
rect 255884 238785 255912 239788
rect 256056 239760 256108 239766
rect 256054 239728 256056 239737
rect 256206 239748 256234 240108
rect 256108 239728 256110 239737
rect 255964 239692 256016 239698
rect 256054 239663 256110 239672
rect 256160 239720 256234 239748
rect 255964 239634 256016 239640
rect 255976 239465 256004 239634
rect 255962 239456 256018 239465
rect 255962 239391 256018 239400
rect 255976 238882 256004 239391
rect 255964 238876 256016 238882
rect 255964 238818 256016 238824
rect 255870 238776 255926 238785
rect 255870 238711 255926 238720
rect 256160 238660 256188 239720
rect 256298 239714 256326 240108
rect 256390 239970 256418 240108
rect 256378 239964 256430 239970
rect 256378 239906 256430 239912
rect 256482 239816 256510 240108
rect 256436 239788 256510 239816
rect 256574 239816 256602 240108
rect 256666 239970 256694 240108
rect 256758 239970 256786 240108
rect 256850 239970 256878 240108
rect 256654 239964 256706 239970
rect 256654 239906 256706 239912
rect 256746 239964 256798 239970
rect 256746 239906 256798 239912
rect 256838 239964 256890 239970
rect 256838 239906 256890 239912
rect 256700 239828 256752 239834
rect 256574 239788 256648 239816
rect 256298 239686 256372 239714
rect 256240 239556 256292 239562
rect 256240 239498 256292 239504
rect 255884 238632 256188 238660
rect 255778 236736 255834 236745
rect 255778 236671 255834 236680
rect 255688 236020 255740 236026
rect 255688 235962 255740 235968
rect 255596 235272 255648 235278
rect 255596 235214 255648 235220
rect 255596 231872 255648 231878
rect 255596 231814 255648 231820
rect 255504 230784 255556 230790
rect 255504 230726 255556 230732
rect 255504 229764 255556 229770
rect 255504 229706 255556 229712
rect 255516 221950 255544 229706
rect 255608 223174 255636 231814
rect 255700 231441 255728 235962
rect 255884 231854 255912 238632
rect 256252 238592 256280 239498
rect 255792 231826 255912 231854
rect 255976 238564 256280 238592
rect 255976 231854 256004 238564
rect 255976 231826 256280 231854
rect 255686 231432 255742 231441
rect 255686 231367 255742 231376
rect 255792 230489 255820 231826
rect 255778 230480 255834 230489
rect 255778 230415 255834 230424
rect 256146 230480 256202 230489
rect 256146 230415 256202 230424
rect 256160 229566 256188 230415
rect 256148 229560 256200 229566
rect 256148 229502 256200 229508
rect 255596 223168 255648 223174
rect 255596 223110 255648 223116
rect 256148 223168 256200 223174
rect 256148 223110 256200 223116
rect 256054 222048 256110 222057
rect 256054 221983 256110 221992
rect 255504 221944 255556 221950
rect 255504 221886 255556 221892
rect 255964 221944 256016 221950
rect 255964 221886 256016 221892
rect 255412 157684 255464 157690
rect 255412 157626 255464 157632
rect 255976 146674 256004 221886
rect 256068 148753 256096 221983
rect 256160 161158 256188 223110
rect 256252 220289 256280 231826
rect 256344 229770 256372 239686
rect 256436 231198 256464 239788
rect 256516 238740 256568 238746
rect 256516 238682 256568 238688
rect 256528 237250 256556 238682
rect 256516 237244 256568 237250
rect 256516 237186 256568 237192
rect 256620 231878 256648 239788
rect 256700 239770 256752 239776
rect 256792 239828 256844 239834
rect 256792 239770 256844 239776
rect 256712 238542 256740 239770
rect 256804 239578 256832 239770
rect 256942 239748 256970 240108
rect 257034 239902 257062 240108
rect 257126 239970 257154 240108
rect 257114 239964 257166 239970
rect 257114 239906 257166 239912
rect 257022 239896 257074 239902
rect 257218 239850 257246 240108
rect 257022 239838 257074 239844
rect 257172 239822 257246 239850
rect 256942 239720 257016 239748
rect 257172 239737 257200 239822
rect 256804 239550 256924 239578
rect 256792 239488 256844 239494
rect 256792 239430 256844 239436
rect 256700 238536 256752 238542
rect 256700 238478 256752 238484
rect 256804 234818 256832 239430
rect 256712 234790 256832 234818
rect 256608 231872 256660 231878
rect 256608 231814 256660 231820
rect 256424 231192 256476 231198
rect 256424 231134 256476 231140
rect 256516 230784 256568 230790
rect 256516 230726 256568 230732
rect 256332 229764 256384 229770
rect 256332 229706 256384 229712
rect 256238 220280 256294 220289
rect 256238 220215 256294 220224
rect 256252 214713 256280 220215
rect 256528 219230 256556 230726
rect 256712 227390 256740 234790
rect 256792 234728 256844 234734
rect 256792 234670 256844 234676
rect 256700 227384 256752 227390
rect 256700 227326 256752 227332
rect 256712 223574 256740 227326
rect 256620 223546 256740 223574
rect 256516 219224 256568 219230
rect 256516 219166 256568 219172
rect 256238 214704 256294 214713
rect 256238 214639 256294 214648
rect 256528 183598 256556 219166
rect 256240 183592 256292 183598
rect 256240 183534 256292 183540
rect 256516 183592 256568 183598
rect 256516 183534 256568 183540
rect 256148 161152 256200 161158
rect 256148 161094 256200 161100
rect 256252 158846 256280 183534
rect 256240 158840 256292 158846
rect 256240 158782 256292 158788
rect 256054 148744 256110 148753
rect 256054 148679 256110 148688
rect 255964 146668 256016 146674
rect 255964 146610 256016 146616
rect 255318 142896 255374 142905
rect 255318 142831 255320 142840
rect 255372 142831 255374 142840
rect 255320 142802 255372 142808
rect 255228 131096 255280 131102
rect 255228 131038 255280 131044
rect 255240 130422 255268 131038
rect 255228 130416 255280 130422
rect 255228 130358 255280 130364
rect 256056 128240 256108 128246
rect 256056 128182 256108 128188
rect 256068 127702 256096 128182
rect 256620 127702 256648 223546
rect 256804 223378 256832 234670
rect 256896 232014 256924 239550
rect 256884 232008 256936 232014
rect 256884 231950 256936 231956
rect 256884 231872 256936 231878
rect 256884 231814 256936 231820
rect 256896 223446 256924 231814
rect 256988 231577 257016 239720
rect 257158 239728 257214 239737
rect 257310 239714 257338 240108
rect 257402 239902 257430 240108
rect 257494 239970 257522 240108
rect 257482 239964 257534 239970
rect 257482 239906 257534 239912
rect 257390 239896 257442 239902
rect 257390 239838 257442 239844
rect 257586 239816 257614 240108
rect 257540 239788 257614 239816
rect 257678 239816 257706 240108
rect 257770 239970 257798 240108
rect 257758 239964 257810 239970
rect 257758 239906 257810 239912
rect 257862 239850 257890 240108
rect 257954 239970 257982 240108
rect 257942 239964 257994 239970
rect 257942 239906 257994 239912
rect 258046 239902 258074 240108
rect 257816 239822 257890 239850
rect 258034 239896 258086 239902
rect 258138 239873 258166 240108
rect 258034 239838 258086 239844
rect 258124 239864 258180 239873
rect 257678 239788 257752 239816
rect 257310 239686 257384 239714
rect 257158 239663 257214 239672
rect 257068 239624 257120 239630
rect 257068 239566 257120 239572
rect 257080 237374 257108 239566
rect 257172 238610 257200 239663
rect 257252 239624 257304 239630
rect 257252 239566 257304 239572
rect 257264 238785 257292 239566
rect 257250 238776 257306 238785
rect 257250 238711 257306 238720
rect 257160 238604 257212 238610
rect 257160 238546 257212 238552
rect 257080 237346 257292 237374
rect 257264 235793 257292 237346
rect 257356 236910 257384 239686
rect 257436 239692 257488 239698
rect 257436 239634 257488 239640
rect 257344 236904 257396 236910
rect 257344 236846 257396 236852
rect 257356 236706 257384 236846
rect 257344 236700 257396 236706
rect 257344 236642 257396 236648
rect 257250 235784 257306 235793
rect 257250 235719 257306 235728
rect 257264 235385 257292 235719
rect 257250 235376 257306 235385
rect 257250 235311 257306 235320
rect 256974 231568 257030 231577
rect 256974 231503 257030 231512
rect 256988 231130 257016 231503
rect 256976 231124 257028 231130
rect 256976 231066 257028 231072
rect 257448 226334 257476 239634
rect 257540 239034 257568 239788
rect 257620 239692 257672 239698
rect 257620 239634 257672 239640
rect 257632 239465 257660 239634
rect 257724 239562 257752 239788
rect 257712 239556 257764 239562
rect 257712 239498 257764 239504
rect 257618 239456 257674 239465
rect 257674 239414 257752 239442
rect 257618 239391 257674 239400
rect 257540 239006 257660 239034
rect 257528 238876 257580 238882
rect 257528 238818 257580 238824
rect 257540 235113 257568 238818
rect 257526 235104 257582 235113
rect 257526 235039 257582 235048
rect 257632 227050 257660 239006
rect 257724 237368 257752 239414
rect 257816 237590 257844 239822
rect 258124 239799 258180 239808
rect 257896 239760 257948 239766
rect 258230 239748 258258 240108
rect 258322 239902 258350 240108
rect 258414 239970 258442 240108
rect 258402 239964 258454 239970
rect 258402 239906 258454 239912
rect 258310 239896 258362 239902
rect 258310 239838 258362 239844
rect 258506 239816 258534 240108
rect 258598 239902 258626 240108
rect 258690 239902 258718 240108
rect 258782 239970 258810 240108
rect 258874 239970 258902 240108
rect 258770 239964 258822 239970
rect 258770 239906 258822 239912
rect 258862 239964 258914 239970
rect 258862 239906 258914 239912
rect 258586 239896 258638 239902
rect 258586 239838 258638 239844
rect 258678 239896 258730 239902
rect 258966 239850 258994 240108
rect 259058 239902 259086 240108
rect 259150 239970 259178 240108
rect 259138 239964 259190 239970
rect 259138 239906 259190 239912
rect 258678 239838 258730 239844
rect 257896 239702 257948 239708
rect 258092 239720 258258 239748
rect 258414 239788 258534 239816
rect 258920 239822 258994 239850
rect 259046 239896 259098 239902
rect 259046 239838 259098 239844
rect 257804 237584 257856 237590
rect 257804 237526 257856 237532
rect 257724 237340 257844 237368
rect 257712 236836 257764 236842
rect 257712 236778 257764 236784
rect 257724 230518 257752 236778
rect 257712 230512 257764 230518
rect 257712 230454 257764 230460
rect 257620 227044 257672 227050
rect 257620 226986 257672 226992
rect 257448 226306 257752 226334
rect 256884 223440 256936 223446
rect 256884 223382 256936 223388
rect 257344 223440 257396 223446
rect 257344 223382 257396 223388
rect 256792 223372 256844 223378
rect 256792 223314 256844 223320
rect 257356 145790 257384 223382
rect 257436 223372 257488 223378
rect 257436 223314 257488 223320
rect 257448 161265 257476 223314
rect 257724 223310 257752 226306
rect 257712 223304 257764 223310
rect 257712 223246 257764 223252
rect 257724 219434 257752 223246
rect 257540 219406 257752 219434
rect 257540 202201 257568 219406
rect 257526 202192 257582 202201
rect 257526 202127 257582 202136
rect 257816 187746 257844 237340
rect 257908 234734 257936 239702
rect 257988 239556 258040 239562
rect 257988 239498 258040 239504
rect 258000 238728 258028 239498
rect 258092 239465 258120 239720
rect 258172 239624 258224 239630
rect 258414 239612 258442 239788
rect 258724 239760 258776 239766
rect 258538 239728 258594 239737
rect 258776 239708 258856 239714
rect 258724 239702 258856 239708
rect 258736 239686 258856 239702
rect 258538 239663 258540 239672
rect 258592 239663 258594 239672
rect 258540 239634 258592 239640
rect 258724 239624 258776 239630
rect 258414 239584 258488 239612
rect 258172 239566 258224 239572
rect 258078 239456 258134 239465
rect 258078 239391 258134 239400
rect 258184 239034 258212 239566
rect 258460 239544 258488 239584
rect 258724 239566 258776 239572
rect 258460 239516 258580 239544
rect 258356 239488 258408 239494
rect 258356 239430 258408 239436
rect 258092 239006 258212 239034
rect 258092 238882 258120 239006
rect 258080 238876 258132 238882
rect 258080 238818 258132 238824
rect 258172 238740 258224 238746
rect 258000 238700 258120 238728
rect 257988 238604 258040 238610
rect 257988 238546 258040 238552
rect 257896 234728 257948 234734
rect 257896 234670 257948 234676
rect 257896 234592 257948 234598
rect 257896 234534 257948 234540
rect 257908 233850 257936 234534
rect 257896 233844 257948 233850
rect 257896 233786 257948 233792
rect 257528 187740 257580 187746
rect 257528 187682 257580 187688
rect 257804 187740 257856 187746
rect 257804 187682 257856 187688
rect 257434 161256 257490 161265
rect 257434 161191 257490 161200
rect 257540 150113 257568 187682
rect 258000 186386 258028 238546
rect 258092 231878 258120 238700
rect 258172 238682 258224 238688
rect 258080 231872 258132 231878
rect 258080 231814 258132 231820
rect 257620 186380 257672 186386
rect 257620 186322 257672 186328
rect 257988 186380 258040 186386
rect 257988 186322 258040 186328
rect 257632 160993 257660 186322
rect 257618 160984 257674 160993
rect 257618 160919 257674 160928
rect 257526 150104 257582 150113
rect 257526 150039 257582 150048
rect 257344 145784 257396 145790
rect 257344 145726 257396 145732
rect 258184 145722 258212 238682
rect 258262 238368 258318 238377
rect 258262 238303 258318 238312
rect 258276 236842 258304 238303
rect 258368 238105 258396 239430
rect 258448 239420 258500 239426
rect 258448 239362 258500 239368
rect 258354 238096 258410 238105
rect 258354 238031 258410 238040
rect 258264 236836 258316 236842
rect 258264 236778 258316 236784
rect 258264 236700 258316 236706
rect 258264 236642 258316 236648
rect 258276 227254 258304 236642
rect 258264 227248 258316 227254
rect 258264 227190 258316 227196
rect 258368 223574 258396 238031
rect 258460 237930 258488 239362
rect 258448 237924 258500 237930
rect 258448 237866 258500 237872
rect 258552 237374 258580 239516
rect 258460 237346 258580 237374
rect 258632 237380 258684 237386
rect 258460 236502 258488 237346
rect 258736 237374 258764 239566
rect 258828 239465 258856 239686
rect 258814 239456 258870 239465
rect 258814 239391 258870 239400
rect 258828 238746 258856 239391
rect 258816 238740 258868 238746
rect 258816 238682 258868 238688
rect 258736 237346 258856 237374
rect 258632 237322 258684 237328
rect 258448 236496 258500 236502
rect 258448 236438 258500 236444
rect 258460 234666 258488 236438
rect 258448 234660 258500 234666
rect 258448 234602 258500 234608
rect 258644 223650 258672 237322
rect 258724 234320 258776 234326
rect 258724 234262 258776 234268
rect 258736 233986 258764 234262
rect 258724 233980 258776 233986
rect 258724 233922 258776 233928
rect 258828 231169 258856 237346
rect 258920 236706 258948 239822
rect 259242 239816 259270 240108
rect 259196 239788 259270 239816
rect 259000 239760 259052 239766
rect 259000 239702 259052 239708
rect 259012 236960 259040 239702
rect 259092 239624 259144 239630
rect 259092 239566 259144 239572
rect 259104 238785 259132 239566
rect 259090 238776 259146 238785
rect 259090 238711 259146 238720
rect 259012 236932 259132 236960
rect 258998 236736 259054 236745
rect 258908 236700 258960 236706
rect 258998 236671 259054 236680
rect 258908 236642 258960 236648
rect 258814 231160 258870 231169
rect 258814 231095 258870 231104
rect 258632 223644 258684 223650
rect 258632 223586 258684 223592
rect 258368 223546 258580 223574
rect 258172 145716 258224 145722
rect 258172 145658 258224 145664
rect 258552 140729 258580 223546
rect 258644 219434 258672 223586
rect 258816 223576 258868 223582
rect 258816 223518 258868 223524
rect 258644 219406 258764 219434
rect 258736 145586 258764 219406
rect 258828 148889 258856 223518
rect 259012 219434 259040 236671
rect 259104 233234 259132 236932
rect 259196 233345 259224 239788
rect 259334 239748 259362 240108
rect 259426 239902 259454 240108
rect 259518 239902 259546 240108
rect 259414 239896 259466 239902
rect 259414 239838 259466 239844
rect 259506 239896 259558 239902
rect 259506 239838 259558 239844
rect 259288 239720 259362 239748
rect 259460 239760 259512 239766
rect 259458 239728 259460 239737
rect 259512 239728 259514 239737
rect 259288 237386 259316 239720
rect 259610 239714 259638 240108
rect 259702 239970 259730 240108
rect 259690 239964 259742 239970
rect 259690 239906 259742 239912
rect 259794 239748 259822 240108
rect 259886 239970 259914 240108
rect 259978 239970 260006 240108
rect 259874 239964 259926 239970
rect 259874 239906 259926 239912
rect 259966 239964 260018 239970
rect 259966 239906 260018 239912
rect 260070 239850 260098 240108
rect 260162 239970 260190 240108
rect 260150 239964 260202 239970
rect 260150 239906 260202 239912
rect 260070 239822 260144 239850
rect 259794 239720 259868 239748
rect 259610 239686 259684 239714
rect 259458 239663 259514 239672
rect 259368 239624 259420 239630
rect 259368 239566 259420 239572
rect 259380 238202 259408 239566
rect 259368 238196 259420 238202
rect 259368 238138 259420 238144
rect 259276 237380 259328 237386
rect 259276 237322 259328 237328
rect 259276 236904 259328 236910
rect 259276 236846 259328 236852
rect 259288 234326 259316 236846
rect 259276 234320 259328 234326
rect 259276 234262 259328 234268
rect 259182 233336 259238 233345
rect 259182 233271 259238 233280
rect 259104 233206 259224 233234
rect 259196 223582 259224 233206
rect 259274 232384 259330 232393
rect 259274 232319 259330 232328
rect 259288 230654 259316 232319
rect 259380 231606 259408 238138
rect 259368 231600 259420 231606
rect 259368 231542 259420 231548
rect 259472 230722 259500 239663
rect 259552 239624 259604 239630
rect 259656 239612 259684 239686
rect 259656 239584 259776 239612
rect 259552 239566 259604 239572
rect 259564 238542 259592 239566
rect 259748 239465 259776 239584
rect 259734 239456 259790 239465
rect 259644 239420 259696 239426
rect 259734 239391 259790 239400
rect 259644 239362 259696 239368
rect 259552 238536 259604 238542
rect 259656 238513 259684 239362
rect 259736 239352 259788 239358
rect 259736 239294 259788 239300
rect 259748 238610 259776 239294
rect 259736 238604 259788 238610
rect 259736 238546 259788 238552
rect 259552 238478 259604 238484
rect 259642 238504 259698 238513
rect 259642 238439 259698 238448
rect 259460 230716 259512 230722
rect 259460 230658 259512 230664
rect 259276 230648 259328 230654
rect 259276 230590 259328 230596
rect 259288 225894 259316 230590
rect 259656 226982 259684 238439
rect 259734 238368 259790 238377
rect 259734 238303 259736 238312
rect 259788 238303 259790 238312
rect 259736 238274 259788 238280
rect 259840 235890 259868 239720
rect 260012 239692 260064 239698
rect 259932 239652 260012 239680
rect 259828 235884 259880 235890
rect 259828 235826 259880 235832
rect 259734 232248 259790 232257
rect 259734 232183 259790 232192
rect 259644 226976 259696 226982
rect 259644 226918 259696 226924
rect 259748 226914 259776 232183
rect 259828 229628 259880 229634
rect 259828 229570 259880 229576
rect 259736 226908 259788 226914
rect 259736 226850 259788 226856
rect 259276 225888 259328 225894
rect 259276 225830 259328 225836
rect 259184 223576 259236 223582
rect 259184 223518 259236 223524
rect 259368 223508 259420 223514
rect 259368 223450 259420 223456
rect 259380 223174 259408 223450
rect 259368 223168 259420 223174
rect 259368 223110 259420 223116
rect 258920 219406 259040 219434
rect 258920 157758 258948 219406
rect 258908 157752 258960 157758
rect 258908 157694 258960 157700
rect 258814 148880 258870 148889
rect 258814 148815 258870 148824
rect 258724 145580 258776 145586
rect 258724 145522 258776 145528
rect 259840 144634 259868 229570
rect 259932 227526 259960 239652
rect 260012 239634 260064 239640
rect 260012 239556 260064 239562
rect 260012 239498 260064 239504
rect 260024 228410 260052 239498
rect 260116 234598 260144 239822
rect 260254 239816 260282 240108
rect 260208 239788 260282 239816
rect 260104 234592 260156 234598
rect 260104 234534 260156 234540
rect 260012 228404 260064 228410
rect 260012 228346 260064 228352
rect 260024 227662 260052 228346
rect 260012 227656 260064 227662
rect 260208 227644 260236 239788
rect 260346 239612 260374 240108
rect 260438 239970 260466 240108
rect 260426 239964 260478 239970
rect 260426 239906 260478 239912
rect 260530 239873 260558 240108
rect 260622 239902 260650 240108
rect 260610 239896 260662 239902
rect 260516 239864 260572 239873
rect 260610 239838 260662 239844
rect 260516 239799 260572 239808
rect 260472 239760 260524 239766
rect 260472 239702 260524 239708
rect 260714 239714 260742 240108
rect 260806 239873 260834 240108
rect 260898 239970 260926 240108
rect 260886 239964 260938 239970
rect 260886 239906 260938 239912
rect 260792 239864 260848 239873
rect 260990 239850 261018 240108
rect 260944 239822 261018 239850
rect 260848 239808 260880 239816
rect 260792 239799 260880 239808
rect 260806 239788 260880 239799
rect 260346 239584 260420 239612
rect 260288 239488 260340 239494
rect 260288 239430 260340 239436
rect 260300 239358 260328 239430
rect 260288 239352 260340 239358
rect 260288 239294 260340 239300
rect 260392 238785 260420 239584
rect 260484 239544 260512 239702
rect 260714 239686 260788 239714
rect 260656 239624 260708 239630
rect 260656 239566 260708 239572
rect 260484 239516 260604 239544
rect 260470 239456 260526 239465
rect 260470 239391 260526 239400
rect 260378 238776 260434 238785
rect 260378 238711 260434 238720
rect 260378 238640 260434 238649
rect 260378 238575 260434 238584
rect 260392 238134 260420 238575
rect 260288 238128 260340 238134
rect 260288 238070 260340 238076
rect 260380 238128 260432 238134
rect 260380 238070 260432 238076
rect 260300 231062 260328 238070
rect 260484 236473 260512 239391
rect 260576 238898 260604 239516
rect 260668 239465 260696 239566
rect 260654 239456 260710 239465
rect 260654 239391 260710 239400
rect 260576 238870 260696 238898
rect 260564 238808 260616 238814
rect 260564 238750 260616 238756
rect 260576 238105 260604 238750
rect 260668 238649 260696 238870
rect 260654 238640 260710 238649
rect 260654 238575 260710 238584
rect 260760 238490 260788 239686
rect 260668 238462 260788 238490
rect 260562 238096 260618 238105
rect 260562 238031 260618 238040
rect 260470 236464 260526 236473
rect 260470 236399 260526 236408
rect 260668 234784 260696 238462
rect 260746 238368 260802 238377
rect 260746 238303 260802 238312
rect 260576 234756 260696 234784
rect 260288 231056 260340 231062
rect 260288 230998 260340 231004
rect 260012 227598 260064 227604
rect 260116 227616 260236 227644
rect 259920 227520 259972 227526
rect 259920 227462 259972 227468
rect 259932 227361 259960 227462
rect 259918 227352 259974 227361
rect 259918 227287 259974 227296
rect 260116 223417 260144 227616
rect 260576 227526 260604 234756
rect 260564 227520 260616 227526
rect 260564 227462 260616 227468
rect 260576 226334 260604 227462
rect 260300 226306 260604 226334
rect 260196 224936 260248 224942
rect 260196 224878 260248 224884
rect 260102 223408 260158 223417
rect 260102 223343 260158 223352
rect 259828 144628 259880 144634
rect 259828 144570 259880 144576
rect 260116 144566 260144 223343
rect 260208 161401 260236 224878
rect 260300 206378 260328 226306
rect 260288 206372 260340 206378
rect 260288 206314 260340 206320
rect 260760 175234 260788 238303
rect 260852 229634 260880 239788
rect 260944 238864 260972 239822
rect 261082 239816 261110 240108
rect 261174 239970 261202 240108
rect 261266 239970 261294 240108
rect 261162 239964 261214 239970
rect 261162 239906 261214 239912
rect 261254 239964 261306 239970
rect 261254 239906 261306 239912
rect 261358 239816 261386 240108
rect 261450 239873 261478 240108
rect 261082 239788 261156 239816
rect 261024 239692 261076 239698
rect 261024 239634 261076 239640
rect 261036 239494 261064 239634
rect 261024 239488 261076 239494
rect 261024 239430 261076 239436
rect 261128 238882 261156 239788
rect 261312 239788 261386 239816
rect 261436 239864 261492 239873
rect 261436 239799 261492 239808
rect 261312 239714 261340 239788
rect 261542 239748 261570 240108
rect 261634 239902 261662 240108
rect 261622 239896 261674 239902
rect 261622 239838 261674 239844
rect 261726 239816 261754 240108
rect 261818 239970 261846 240108
rect 261806 239964 261858 239970
rect 261806 239906 261858 239912
rect 261910 239816 261938 240108
rect 262002 239970 262030 240108
rect 261990 239964 262042 239970
rect 261990 239906 262042 239912
rect 262094 239816 262122 240108
rect 262186 239970 262214 240108
rect 262174 239964 262226 239970
rect 262174 239906 262226 239912
rect 262278 239850 262306 240108
rect 262370 239902 262398 240108
rect 261726 239788 261800 239816
rect 261910 239788 261984 239816
rect 261390 239728 261446 239737
rect 261312 239686 261390 239714
rect 261390 239663 261446 239672
rect 261496 239720 261570 239748
rect 261666 239728 261722 239737
rect 261300 239624 261352 239630
rect 261300 239566 261352 239572
rect 261208 239488 261260 239494
rect 261208 239430 261260 239436
rect 261116 238876 261168 238882
rect 260944 238836 261064 238864
rect 261036 238762 261064 238836
rect 261116 238818 261168 238824
rect 261036 238734 261156 238762
rect 261022 238640 261078 238649
rect 261022 238575 261078 238584
rect 261036 238377 261064 238575
rect 261022 238368 261078 238377
rect 261022 238303 261078 238312
rect 261024 237380 261076 237386
rect 261024 237322 261076 237328
rect 261036 237114 261064 237322
rect 261024 237108 261076 237114
rect 261024 237050 261076 237056
rect 261024 236972 261076 236978
rect 261024 236914 261076 236920
rect 261036 236298 261064 236914
rect 261024 236292 261076 236298
rect 261024 236234 261076 236240
rect 261128 231854 261156 238734
rect 261220 236094 261248 239430
rect 261312 238746 261340 239566
rect 261392 238876 261444 238882
rect 261392 238818 261444 238824
rect 261300 238740 261352 238746
rect 261300 238682 261352 238688
rect 261298 238640 261354 238649
rect 261298 238575 261354 238584
rect 261312 237998 261340 238575
rect 261300 237992 261352 237998
rect 261300 237934 261352 237940
rect 261404 236201 261432 238818
rect 261390 236192 261446 236201
rect 261496 236162 261524 239720
rect 261666 239663 261722 239672
rect 261680 239630 261708 239663
rect 261668 239624 261720 239630
rect 261668 239566 261720 239572
rect 261576 238808 261628 238814
rect 261576 238750 261628 238756
rect 261588 238406 261616 238750
rect 261576 238400 261628 238406
rect 261576 238342 261628 238348
rect 261576 237856 261628 237862
rect 261576 237798 261628 237804
rect 261588 237658 261616 237798
rect 261576 237652 261628 237658
rect 261576 237594 261628 237600
rect 261680 237538 261708 239566
rect 261588 237510 261708 237538
rect 261390 236127 261446 236136
rect 261484 236156 261536 236162
rect 261484 236098 261536 236104
rect 261208 236088 261260 236094
rect 261588 236042 261616 237510
rect 261772 236842 261800 239788
rect 261852 239692 261904 239698
rect 261852 239634 261904 239640
rect 261760 236836 261812 236842
rect 261760 236778 261812 236784
rect 261864 236722 261892 239634
rect 261956 239465 261984 239788
rect 262048 239788 262122 239816
rect 262232 239822 262306 239850
rect 262358 239896 262410 239902
rect 262358 239838 262410 239844
rect 261942 239456 261998 239465
rect 261942 239391 261998 239400
rect 261208 236030 261260 236036
rect 260944 231826 261156 231854
rect 261496 236014 261616 236042
rect 261680 236694 261892 236722
rect 260840 229628 260892 229634
rect 260840 229570 260892 229576
rect 260944 226914 260972 231826
rect 260932 226908 260984 226914
rect 260932 226850 260984 226856
rect 260930 226264 260986 226273
rect 260930 226199 260986 226208
rect 260944 225622 260972 226199
rect 260932 225616 260984 225622
rect 260932 225558 260984 225564
rect 260840 184204 260892 184210
rect 260840 184146 260892 184152
rect 260288 175228 260340 175234
rect 260288 175170 260340 175176
rect 260748 175228 260800 175234
rect 260748 175170 260800 175176
rect 260300 173942 260328 175170
rect 260288 173936 260340 173942
rect 260288 173878 260340 173884
rect 260300 162081 260328 173878
rect 260286 162072 260342 162081
rect 260286 162007 260342 162016
rect 260194 161392 260250 161401
rect 260194 161327 260250 161336
rect 260852 150142 260880 184146
rect 260840 150136 260892 150142
rect 260840 150078 260892 150084
rect 260104 144560 260156 144566
rect 260104 144502 260156 144508
rect 258538 140720 258594 140729
rect 258538 140655 258594 140664
rect 259550 130384 259606 130393
rect 259550 130319 259606 130328
rect 256056 127696 256108 127702
rect 255318 127664 255374 127673
rect 256056 127638 256108 127644
rect 256608 127696 256660 127702
rect 256608 127638 256660 127644
rect 255318 127599 255374 127608
rect 253480 126812 253532 126818
rect 253480 126754 253532 126760
rect 253848 126812 253900 126818
rect 253848 126754 253900 126760
rect 253492 126342 253520 126754
rect 253480 126336 253532 126342
rect 253480 126278 253532 126284
rect 253388 117292 253440 117298
rect 253388 117234 253440 117240
rect 253400 116618 253428 117234
rect 253388 116612 253440 116618
rect 253388 116554 253440 116560
rect 255332 16574 255360 127599
rect 255332 16546 255912 16574
rect 253296 4004 253348 4010
rect 253296 3946 253348 3952
rect 251824 3664 251876 3670
rect 251824 3606 251876 3612
rect 251744 3454 252416 3482
rect 251180 3256 251232 3262
rect 251180 3198 251232 3204
rect 251192 480 251220 3198
rect 252388 480 252416 3454
rect 253124 3262 253152 3878
rect 253216 3862 253612 3890
rect 253584 3398 253612 3862
rect 254676 3664 254728 3670
rect 254676 3606 254728 3612
rect 254768 3664 254820 3670
rect 254768 3606 254820 3612
rect 253480 3392 253532 3398
rect 253480 3334 253532 3340
rect 253572 3392 253624 3398
rect 253572 3334 253624 3340
rect 253112 3256 253164 3262
rect 253112 3198 253164 3204
rect 253492 480 253520 3334
rect 254688 480 254716 3606
rect 254780 3194 254808 3606
rect 254768 3188 254820 3194
rect 254768 3130 254820 3136
rect 255884 480 255912 16546
rect 259564 6914 259592 130319
rect 260852 16574 260880 150078
rect 260944 146169 260972 225558
rect 260930 146160 260986 146169
rect 260930 146095 260986 146104
rect 261496 124098 261524 236014
rect 261680 233073 261708 236694
rect 261852 236292 261904 236298
rect 261852 236234 261904 236240
rect 261864 235226 261892 236234
rect 262048 235346 262076 239788
rect 262128 239556 262180 239562
rect 262128 239498 262180 239504
rect 262140 238241 262168 239498
rect 262232 238456 262260 239822
rect 262312 239760 262364 239766
rect 262462 239748 262490 240108
rect 262554 239902 262582 240108
rect 262542 239896 262594 239902
rect 262646 239873 262674 240108
rect 262738 239970 262766 240108
rect 262726 239964 262778 239970
rect 262726 239906 262778 239912
rect 262542 239838 262594 239844
rect 262632 239864 262688 239873
rect 262632 239799 262688 239808
rect 262312 239702 262364 239708
rect 262416 239720 262490 239748
rect 262738 239748 262766 239906
rect 262830 239816 262858 240108
rect 262922 239970 262950 240108
rect 263014 239970 263042 240108
rect 263106 239970 263134 240108
rect 262910 239964 262962 239970
rect 262910 239906 262962 239912
rect 263002 239964 263054 239970
rect 263002 239906 263054 239912
rect 263094 239964 263146 239970
rect 263094 239906 263146 239912
rect 263198 239873 263226 240108
rect 263290 239970 263318 240108
rect 263278 239964 263330 239970
rect 263278 239906 263330 239912
rect 263184 239864 263240 239873
rect 262956 239828 263008 239834
rect 262830 239788 262904 239816
rect 262738 239720 262812 239748
rect 262324 238592 262352 239702
rect 262416 239465 262444 239720
rect 262496 239556 262548 239562
rect 262496 239498 262548 239504
rect 262402 239456 262458 239465
rect 262402 239391 262458 239400
rect 262324 238564 262444 238592
rect 262232 238428 262352 238456
rect 262220 238332 262272 238338
rect 262220 238274 262272 238280
rect 262126 238232 262182 238241
rect 262126 238167 262182 238176
rect 262036 235340 262088 235346
rect 262036 235282 262088 235288
rect 261772 235198 261892 235226
rect 261666 233064 261722 233073
rect 261666 232999 261722 233008
rect 261576 232008 261628 232014
rect 261576 231950 261628 231956
rect 261588 231130 261616 231950
rect 261576 231124 261628 231130
rect 261576 231066 261628 231072
rect 261588 136610 261616 231066
rect 261680 205018 261708 232999
rect 261772 227730 261800 235198
rect 261850 235104 261906 235113
rect 261850 235039 261906 235048
rect 261760 227724 261812 227730
rect 261760 227666 261812 227672
rect 261668 205012 261720 205018
rect 261668 204954 261720 204960
rect 261864 161945 261892 235039
rect 262232 221542 262260 238274
rect 262324 236978 262352 238428
rect 262312 236972 262364 236978
rect 262312 236914 262364 236920
rect 262310 230888 262366 230897
rect 262310 230823 262366 230832
rect 262324 228954 262352 230823
rect 262312 228948 262364 228954
rect 262312 228890 262364 228896
rect 262324 222766 262352 228890
rect 262416 226778 262444 238564
rect 262508 234569 262536 239498
rect 262588 239488 262640 239494
rect 262588 239430 262640 239436
rect 262600 238785 262628 239430
rect 262586 238776 262642 238785
rect 262586 238711 262642 238720
rect 262680 238740 262732 238746
rect 262680 238682 262732 238688
rect 262692 238626 262720 238682
rect 262600 238598 262720 238626
rect 262600 236910 262628 238598
rect 262588 236904 262640 236910
rect 262588 236846 262640 236852
rect 262784 236688 262812 239720
rect 262876 237114 262904 239788
rect 262956 239770 263008 239776
rect 263048 239828 263100 239834
rect 263382 239850 263410 240108
rect 263474 239970 263502 240108
rect 263462 239964 263514 239970
rect 263462 239906 263514 239912
rect 263184 239799 263240 239808
rect 263336 239822 263410 239850
rect 263048 239770 263100 239776
rect 262864 237108 262916 237114
rect 262864 237050 262916 237056
rect 262692 236660 262812 236688
rect 262494 234560 262550 234569
rect 262494 234495 262550 234504
rect 262404 226772 262456 226778
rect 262404 226714 262456 226720
rect 262416 224942 262444 226714
rect 262404 224936 262456 224942
rect 262404 224878 262456 224884
rect 262312 222760 262364 222766
rect 262312 222702 262364 222708
rect 262220 221536 262272 221542
rect 262220 221478 262272 221484
rect 262692 219434 262720 236660
rect 262772 236564 262824 236570
rect 262772 236506 262824 236512
rect 262784 232558 262812 236506
rect 262864 235408 262916 235414
rect 262864 235350 262916 235356
rect 262772 232552 262824 232558
rect 262772 232494 262824 232500
rect 262876 231810 262904 235350
rect 262864 231804 262916 231810
rect 262864 231746 262916 231752
rect 262862 230208 262918 230217
rect 262862 230143 262918 230152
rect 262416 219406 262720 219434
rect 261850 161936 261906 161945
rect 261850 161871 261906 161880
rect 262416 144226 262444 219406
rect 262404 144220 262456 144226
rect 262404 144162 262456 144168
rect 262876 139369 262904 230143
rect 262968 227322 262996 239770
rect 263060 238762 263088 239770
rect 263140 239692 263192 239698
rect 263140 239634 263192 239640
rect 263152 239426 263180 239634
rect 263140 239420 263192 239426
rect 263140 239362 263192 239368
rect 263060 238734 263180 238762
rect 263048 238264 263100 238270
rect 263048 238206 263100 238212
rect 262956 227316 263008 227322
rect 262956 227258 263008 227264
rect 263060 224942 263088 238206
rect 263152 235278 263180 238734
rect 263140 235272 263192 235278
rect 263336 235249 263364 239822
rect 263566 239816 263594 240108
rect 263520 239788 263594 239816
rect 263658 239816 263686 240108
rect 263750 239970 263778 240108
rect 263738 239964 263790 239970
rect 263738 239906 263790 239912
rect 263842 239902 263870 240108
rect 263830 239896 263882 239902
rect 263830 239838 263882 239844
rect 263934 239850 263962 240108
rect 264026 239970 264054 240108
rect 264014 239964 264066 239970
rect 264014 239906 264066 239912
rect 264118 239873 264146 240108
rect 264104 239864 264160 239873
rect 263934 239822 264008 239850
rect 263658 239788 263732 239816
rect 263416 239760 263468 239766
rect 263416 239702 263468 239708
rect 263428 237930 263456 239702
rect 263416 237924 263468 237930
rect 263416 237866 263468 237872
rect 263520 237697 263548 239788
rect 263598 239728 263654 239737
rect 263598 239663 263600 239672
rect 263652 239663 263654 239672
rect 263600 239634 263652 239640
rect 263600 239420 263652 239426
rect 263600 239362 263652 239368
rect 263612 238338 263640 239362
rect 263704 238746 263732 239788
rect 263876 239760 263928 239766
rect 263876 239702 263928 239708
rect 263784 239692 263836 239698
rect 263784 239634 263836 239640
rect 263692 238740 263744 238746
rect 263692 238682 263744 238688
rect 263600 238332 263652 238338
rect 263600 238274 263652 238280
rect 263598 238232 263654 238241
rect 263598 238167 263654 238176
rect 263506 237688 263562 237697
rect 263506 237623 263562 237632
rect 263508 237584 263560 237590
rect 263508 237526 263560 237532
rect 263140 235214 263192 235220
rect 263322 235240 263378 235249
rect 263322 235175 263378 235184
rect 263520 227118 263548 237526
rect 263508 227112 263560 227118
rect 263508 227054 263560 227060
rect 263048 224936 263100 224942
rect 263048 224878 263100 224884
rect 263046 223544 263102 223553
rect 262956 223508 263008 223514
rect 263046 223479 263102 223488
rect 262956 223450 263008 223456
rect 262968 223310 262996 223450
rect 262956 223304 263008 223310
rect 262956 223246 263008 223252
rect 262956 222760 263008 222766
rect 262956 222702 263008 222708
rect 262968 154465 262996 222702
rect 263060 163577 263088 223479
rect 263612 165073 263640 238167
rect 263796 237697 263824 239634
rect 263782 237688 263838 237697
rect 263692 237652 263744 237658
rect 263782 237623 263838 237632
rect 263692 237594 263744 237600
rect 263704 166297 263732 237594
rect 263796 233889 263824 237623
rect 263782 233880 263838 233889
rect 263782 233815 263838 233824
rect 263784 233708 263836 233714
rect 263784 233650 263836 233656
rect 263796 229022 263824 233650
rect 263888 233234 263916 239702
rect 263980 238610 264008 239822
rect 264104 239799 264160 239808
rect 264210 239714 264238 240108
rect 264302 239816 264330 240108
rect 264394 239970 264422 240108
rect 264382 239964 264434 239970
rect 264382 239906 264434 239912
rect 264486 239816 264514 240108
rect 264302 239788 264376 239816
rect 264210 239686 264284 239714
rect 264060 239624 264112 239630
rect 264060 239566 264112 239572
rect 264152 239624 264204 239630
rect 264152 239566 264204 239572
rect 263968 238604 264020 238610
rect 263968 238546 264020 238552
rect 264072 236609 264100 239566
rect 264164 238785 264192 239566
rect 264150 238776 264206 238785
rect 264150 238711 264206 238720
rect 264256 237590 264284 239686
rect 264244 237584 264296 237590
rect 264244 237526 264296 237532
rect 264058 236600 264114 236609
rect 264058 236535 264114 236544
rect 263888 233206 264008 233234
rect 263980 229094 264008 233206
rect 264348 231854 264376 239788
rect 264440 239788 264514 239816
rect 264440 238202 264468 239788
rect 264578 239714 264606 240108
rect 264670 239873 264698 240108
rect 264656 239864 264712 239873
rect 264762 239850 264790 240108
rect 264854 239970 264882 240108
rect 264946 239970 264974 240108
rect 264842 239964 264894 239970
rect 264842 239906 264894 239912
rect 264934 239964 264986 239970
rect 264934 239906 264986 239912
rect 264762 239822 264928 239850
rect 264656 239799 264712 239808
rect 264900 239737 264928 239822
rect 264886 239728 264942 239737
rect 264578 239686 264698 239714
rect 264520 239624 264572 239630
rect 264670 239612 264698 239686
rect 264796 239692 264848 239698
rect 265038 239714 265066 240108
rect 265130 239902 265158 240108
rect 265118 239896 265170 239902
rect 265118 239838 265170 239844
rect 265038 239686 265112 239714
rect 264886 239663 264942 239672
rect 264796 239634 264848 239640
rect 264520 239566 264572 239572
rect 264624 239584 264698 239612
rect 264428 238196 264480 238202
rect 264428 238138 264480 238144
rect 264532 237300 264560 239566
rect 264624 237374 264652 239584
rect 264702 239456 264758 239465
rect 264702 239391 264704 239400
rect 264756 239391 264758 239400
rect 264704 239362 264756 239368
rect 264716 237658 264744 239362
rect 264704 237652 264756 237658
rect 264704 237594 264756 237600
rect 264624 237346 264744 237374
rect 264532 237272 264652 237300
rect 264348 231826 264468 231854
rect 264440 229094 264468 231826
rect 263980 229066 264376 229094
rect 264440 229066 264560 229094
rect 263784 229016 263836 229022
rect 263784 228958 263836 228964
rect 263796 227866 263824 228958
rect 263784 227860 263836 227866
rect 263784 227802 263836 227808
rect 264244 227860 264296 227866
rect 264244 227802 264296 227808
rect 264152 223644 264204 223650
rect 264152 223586 264204 223592
rect 264164 223514 264192 223586
rect 264152 223508 264204 223514
rect 264152 223450 264204 223456
rect 263690 166288 263746 166297
rect 263690 166223 263746 166232
rect 263598 165064 263654 165073
rect 263598 164999 263654 165008
rect 263046 163568 263102 163577
rect 263046 163503 263102 163512
rect 264256 159186 264284 227802
rect 264348 226273 264376 229066
rect 264428 228880 264480 228886
rect 264428 228822 264480 228828
rect 264334 226264 264390 226273
rect 264334 226199 264390 226208
rect 264348 180033 264376 226199
rect 264440 206310 264468 228822
rect 264532 228750 264560 229066
rect 264520 228744 264572 228750
rect 264520 228686 264572 228692
rect 264532 207738 264560 228686
rect 264624 226817 264652 237272
rect 264716 233714 264744 237346
rect 264704 233708 264756 233714
rect 264704 233650 264756 233656
rect 264808 228886 264836 239634
rect 264886 239456 264942 239465
rect 264886 239391 264942 239400
rect 264900 239358 264928 239391
rect 264888 239352 264940 239358
rect 264888 239294 264940 239300
rect 265084 238610 265112 239686
rect 265222 239680 265250 240108
rect 265314 239748 265342 240108
rect 265406 239873 265434 240108
rect 265498 239902 265526 240108
rect 265590 239970 265618 240108
rect 265682 239970 265710 240108
rect 265578 239964 265630 239970
rect 265578 239906 265630 239912
rect 265670 239964 265722 239970
rect 265670 239906 265722 239912
rect 265486 239896 265538 239902
rect 265392 239864 265448 239873
rect 265774 239850 265802 240108
rect 265486 239838 265538 239844
rect 265392 239799 265448 239808
rect 265624 239828 265676 239834
rect 265624 239770 265676 239776
rect 265728 239822 265802 239850
rect 265532 239760 265584 239766
rect 265314 239720 265388 239748
rect 265222 239652 265296 239680
rect 265162 238776 265218 238785
rect 265162 238711 265218 238720
rect 264980 238604 265032 238610
rect 264980 238546 265032 238552
rect 265072 238604 265124 238610
rect 265072 238546 265124 238552
rect 264992 237454 265020 238546
rect 265072 238332 265124 238338
rect 265072 238274 265124 238280
rect 265084 237658 265112 238274
rect 265072 237652 265124 237658
rect 265072 237594 265124 237600
rect 264980 237448 265032 237454
rect 264980 237390 265032 237396
rect 264978 236736 265034 236745
rect 264978 236671 265034 236680
rect 264796 228880 264848 228886
rect 264796 228822 264848 228828
rect 264610 226808 264666 226817
rect 264610 226743 264666 226752
rect 264520 207732 264572 207738
rect 264520 207674 264572 207680
rect 264428 206304 264480 206310
rect 264428 206246 264480 206252
rect 264992 191049 265020 236671
rect 265072 235204 265124 235210
rect 265072 235146 265124 235152
rect 265084 232354 265112 235146
rect 265072 232348 265124 232354
rect 265072 232290 265124 232296
rect 265176 227186 265204 238711
rect 265268 231849 265296 239652
rect 265360 238116 265388 239720
rect 265530 239728 265532 239737
rect 265584 239728 265586 239737
rect 265440 239692 265492 239698
rect 265530 239663 265586 239672
rect 265440 239634 265492 239640
rect 265452 238338 265480 239634
rect 265440 238332 265492 238338
rect 265440 238274 265492 238280
rect 265360 238088 265480 238116
rect 265348 237652 265400 237658
rect 265348 237594 265400 237600
rect 265254 231840 265310 231849
rect 265254 231775 265310 231784
rect 265164 227180 265216 227186
rect 265164 227122 265216 227128
rect 264978 191040 265034 191049
rect 264978 190975 265034 190984
rect 264334 180024 264390 180033
rect 264334 179959 264390 179968
rect 264244 159180 264296 159186
rect 264244 159122 264296 159128
rect 262954 154456 263010 154465
rect 262954 154391 263010 154400
rect 264244 142928 264296 142934
rect 264244 142870 264296 142876
rect 262862 139360 262918 139369
rect 262862 139295 262918 139304
rect 261576 136604 261628 136610
rect 261576 136546 261628 136552
rect 262128 136604 262180 136610
rect 262128 136546 262180 136552
rect 262140 135998 262168 136546
rect 262128 135992 262180 135998
rect 262128 135934 262180 135940
rect 261484 124092 261536 124098
rect 261484 124034 261536 124040
rect 262128 124092 262180 124098
rect 262128 124034 262180 124040
rect 262140 123486 262168 124034
rect 262128 123480 262180 123486
rect 262128 123422 262180 123428
rect 262220 111104 262272 111110
rect 262220 111046 262272 111052
rect 262232 16574 262260 111046
rect 260852 16546 261800 16574
rect 262232 16546 262536 16574
rect 259472 6886 259592 6914
rect 258264 3392 258316 3398
rect 258264 3334 258316 3340
rect 257068 3324 257120 3330
rect 257068 3266 257120 3272
rect 257080 480 257108 3266
rect 258276 480 258304 3334
rect 259472 480 259500 6886
rect 260656 3188 260708 3194
rect 260656 3130 260708 3136
rect 260668 480 260696 3130
rect 261772 480 261800 16546
rect 240478 354 240590 480
rect 240152 326 240590 354
rect 240478 -960 240590 326
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 354 262536 16546
rect 264152 4140 264204 4146
rect 264152 4082 264204 4088
rect 264164 480 264192 4082
rect 264256 3398 264284 142870
rect 265360 141710 265388 237594
rect 265452 236706 265480 238088
rect 265544 237658 265572 239663
rect 265532 237652 265584 237658
rect 265532 237594 265584 237600
rect 265440 236700 265492 236706
rect 265440 236642 265492 236648
rect 265532 236632 265584 236638
rect 265532 236574 265584 236580
rect 265544 229770 265572 236574
rect 265532 229764 265584 229770
rect 265532 229706 265584 229712
rect 265636 228993 265664 239770
rect 265728 237153 265756 239822
rect 265866 239714 265894 240108
rect 265820 239686 265894 239714
rect 265958 239714 265986 240108
rect 266050 239902 266078 240108
rect 266038 239896 266090 239902
rect 266036 239864 266038 239873
rect 266090 239864 266092 239873
rect 266036 239799 266092 239808
rect 266142 239748 266170 240108
rect 266234 239902 266262 240108
rect 266222 239896 266274 239902
rect 266222 239838 266274 239844
rect 266096 239720 266170 239748
rect 266326 239737 266354 240108
rect 266312 239728 266368 239737
rect 265958 239686 266032 239714
rect 265820 238490 265848 239686
rect 265900 239624 265952 239630
rect 265900 239566 265952 239572
rect 265912 239426 265940 239566
rect 265900 239420 265952 239426
rect 265900 239362 265952 239368
rect 265820 238462 265940 238490
rect 265808 238196 265860 238202
rect 265808 238138 265860 238144
rect 265714 237144 265770 237153
rect 265714 237079 265770 237088
rect 265820 235385 265848 238138
rect 265912 236366 265940 238462
rect 265900 236360 265952 236366
rect 265900 236302 265952 236308
rect 265806 235376 265862 235385
rect 265806 235311 265862 235320
rect 265714 231840 265770 231849
rect 265714 231775 265770 231784
rect 265622 228984 265678 228993
rect 265544 228942 265622 228970
rect 265544 223990 265572 228942
rect 265622 228919 265678 228928
rect 265622 228848 265678 228857
rect 265622 228783 265678 228792
rect 265532 223984 265584 223990
rect 265532 223926 265584 223932
rect 265636 166433 265664 228783
rect 265728 177313 265756 231775
rect 266004 228857 266032 239686
rect 266096 233889 266124 239720
rect 266312 239663 266368 239672
rect 266418 239612 266446 240108
rect 266188 239584 266446 239612
rect 266510 239612 266538 240108
rect 266602 239714 266630 240108
rect 266694 239816 266722 240108
rect 266786 239970 266814 240108
rect 266774 239964 266826 239970
rect 266774 239906 266826 239912
rect 266878 239816 266906 240108
rect 266694 239788 266768 239816
rect 266602 239686 266676 239714
rect 266510 239584 266584 239612
rect 266188 238785 266216 239584
rect 266556 238814 266584 239584
rect 266648 239426 266676 239686
rect 266636 239420 266688 239426
rect 266636 239362 266688 239368
rect 266360 238808 266412 238814
rect 266174 238776 266230 238785
rect 266360 238750 266412 238756
rect 266544 238808 266596 238814
rect 266544 238750 266596 238756
rect 266174 238711 266230 238720
rect 266372 238241 266400 238750
rect 266452 238332 266504 238338
rect 266452 238274 266504 238280
rect 266358 238232 266414 238241
rect 266358 238167 266414 238176
rect 266176 237652 266228 237658
rect 266176 237594 266228 237600
rect 266082 233880 266138 233889
rect 266082 233815 266138 233824
rect 265990 228848 266046 228857
rect 265990 228783 266046 228792
rect 265808 223984 265860 223990
rect 265808 223926 265860 223932
rect 265820 207670 265848 223926
rect 265808 207664 265860 207670
rect 265808 207606 265860 207612
rect 265714 177304 265770 177313
rect 265714 177239 265770 177248
rect 265622 166424 265678 166433
rect 265622 166359 265678 166368
rect 266188 163441 266216 237594
rect 266464 171737 266492 238274
rect 266556 219434 266584 238750
rect 266636 238740 266688 238746
rect 266636 238682 266688 238688
rect 266648 236745 266676 238682
rect 266740 238218 266768 239788
rect 266832 239788 266906 239816
rect 266832 239737 266860 239788
rect 266818 239728 266874 239737
rect 266818 239663 266874 239672
rect 266832 238338 266860 239663
rect 266970 239630 266998 240108
rect 267062 239970 267090 240108
rect 267050 239964 267102 239970
rect 267050 239906 267102 239912
rect 267154 239850 267182 240108
rect 267246 239970 267274 240108
rect 267234 239964 267286 239970
rect 267338 239952 267366 240108
rect 267568 240106 267596 240230
rect 267556 240100 267608 240106
rect 267556 240042 267608 240048
rect 267338 239924 267412 239952
rect 267234 239906 267286 239912
rect 267154 239822 267320 239850
rect 267096 239760 267148 239766
rect 267096 239702 267148 239708
rect 267188 239760 267240 239766
rect 267188 239702 267240 239708
rect 266958 239624 267010 239630
rect 266958 239566 267010 239572
rect 266820 238332 266872 238338
rect 266820 238274 266872 238280
rect 266740 238190 266952 238218
rect 266820 238128 266872 238134
rect 266820 238070 266872 238076
rect 266728 237992 266780 237998
rect 266728 237934 266780 237940
rect 266740 237522 266768 237934
rect 266832 237522 266860 238070
rect 266728 237516 266780 237522
rect 266728 237458 266780 237464
rect 266820 237516 266872 237522
rect 266820 237458 266872 237464
rect 266924 237153 266952 238190
rect 267004 238196 267056 238202
rect 267004 238138 267056 238144
rect 267016 237833 267044 238138
rect 267002 237824 267058 237833
rect 267002 237759 267058 237768
rect 266910 237144 266966 237153
rect 266910 237079 266966 237088
rect 266912 236836 266964 236842
rect 266912 236778 266964 236784
rect 266634 236736 266690 236745
rect 266634 236671 266690 236680
rect 266820 236360 266872 236366
rect 266820 236302 266872 236308
rect 266832 234025 266860 236302
rect 266924 235521 266952 236778
rect 266910 235512 266966 235521
rect 266910 235447 266966 235456
rect 267108 235260 267136 239702
rect 267200 239494 267228 239702
rect 267292 239494 267320 239822
rect 267188 239488 267240 239494
rect 267188 239430 267240 239436
rect 267280 239488 267332 239494
rect 267280 239430 267332 239436
rect 267280 238740 267332 238746
rect 267280 238682 267332 238688
rect 267292 237386 267320 238682
rect 267280 237380 267332 237386
rect 267280 237322 267332 237328
rect 267280 236088 267332 236094
rect 267280 236030 267332 236036
rect 267108 235232 267228 235260
rect 267002 235104 267058 235113
rect 267002 235039 267058 235048
rect 266818 234016 266874 234025
rect 266818 233951 266874 233960
rect 266556 219406 266768 219434
rect 266740 202162 266768 219406
rect 266728 202156 266780 202162
rect 266728 202098 266780 202104
rect 266450 171728 266506 171737
rect 266450 171663 266506 171672
rect 267016 169153 267044 235039
rect 267200 230432 267228 235232
rect 267292 235210 267320 236030
rect 267280 235204 267332 235210
rect 267280 235146 267332 235152
rect 267200 230404 267320 230432
rect 267186 229936 267242 229945
rect 267186 229871 267242 229880
rect 267096 225412 267148 225418
rect 267096 225354 267148 225360
rect 267108 173233 267136 225354
rect 267200 175982 267228 229871
rect 267292 227497 267320 230404
rect 267384 228721 267412 239924
rect 267556 239420 267608 239426
rect 267660 239408 267688 260063
rect 267738 250472 267794 250481
rect 267738 250407 267794 250416
rect 267752 241641 267780 250407
rect 268014 247616 268070 247625
rect 268014 247551 268070 247560
rect 267922 246392 267978 246401
rect 267922 246327 267978 246336
rect 267738 241632 267794 241641
rect 267738 241567 267794 241576
rect 267740 240916 267792 240922
rect 267740 240858 267792 240864
rect 267752 240666 267780 240858
rect 267752 240638 267872 240666
rect 267738 240272 267794 240281
rect 267738 240207 267794 240216
rect 267752 239834 267780 240207
rect 267740 239828 267792 239834
rect 267740 239770 267792 239776
rect 267740 239488 267792 239494
rect 267740 239430 267792 239436
rect 267608 239380 267688 239408
rect 267556 239362 267608 239368
rect 267464 238332 267516 238338
rect 267464 238274 267516 238280
rect 267370 228712 267426 228721
rect 267370 228647 267426 228656
rect 267278 227488 267334 227497
rect 267278 227423 267334 227432
rect 267188 175976 267240 175982
rect 267188 175918 267240 175924
rect 267292 173369 267320 227423
rect 267384 225418 267412 228647
rect 267372 225412 267424 225418
rect 267372 225354 267424 225360
rect 267476 182889 267504 238274
rect 267462 182880 267518 182889
rect 267462 182815 267518 182824
rect 267278 173360 267334 173369
rect 267278 173295 267334 173304
rect 267094 173224 267150 173233
rect 267094 173159 267150 173168
rect 267002 169144 267058 169153
rect 267002 169079 267058 169088
rect 267568 164937 267596 239362
rect 267648 234592 267700 234598
rect 267648 234534 267700 234540
rect 267660 233714 267688 234534
rect 267648 233708 267700 233714
rect 267648 233650 267700 233656
rect 267752 223574 267780 239430
rect 267844 238814 267872 240638
rect 267936 240582 267964 246327
rect 267924 240576 267976 240582
rect 267924 240518 267976 240524
rect 267924 240304 267976 240310
rect 267924 240246 267976 240252
rect 267936 240145 267964 240246
rect 267922 240136 267978 240145
rect 267922 240071 267978 240080
rect 268028 240009 268056 247551
rect 268290 243672 268346 243681
rect 268290 243607 268346 243616
rect 268106 242312 268162 242321
rect 268106 242247 268162 242256
rect 268120 240088 268148 242247
rect 268198 241632 268254 241641
rect 268198 241567 268254 241576
rect 268212 240378 268240 241567
rect 268304 240446 268332 243607
rect 268292 240440 268344 240446
rect 268292 240382 268344 240388
rect 268200 240372 268252 240378
rect 268200 240314 268252 240320
rect 268200 240100 268252 240106
rect 268120 240060 268200 240088
rect 268200 240042 268252 240048
rect 268014 240000 268070 240009
rect 268014 239935 268070 239944
rect 268108 239964 268160 239970
rect 268108 239906 268160 239912
rect 268016 239692 268068 239698
rect 268016 239634 268068 239640
rect 267832 238808 267884 238814
rect 267832 238750 267884 238756
rect 267922 235512 267978 235521
rect 267922 235447 267978 235456
rect 267830 235240 267886 235249
rect 267830 235175 267886 235184
rect 267660 223546 267780 223574
rect 267660 178673 267688 223546
rect 267646 178664 267702 178673
rect 267646 178599 267702 178608
rect 267554 164928 267610 164937
rect 267554 164863 267610 164872
rect 266174 163432 266230 163441
rect 266174 163367 266230 163376
rect 267844 155553 267872 235175
rect 267936 155689 267964 235447
rect 268028 229945 268056 239634
rect 268120 235113 268148 239906
rect 268212 238338 268240 240042
rect 268396 239986 268424 285110
rect 268936 285058 268988 285064
rect 268936 284980 268988 284986
rect 268936 284922 268988 284928
rect 268474 265568 268530 265577
rect 268474 265503 268530 265512
rect 268488 243681 268516 265503
rect 268566 257408 268622 257417
rect 268566 257343 268622 257352
rect 268474 243672 268530 243681
rect 268474 243607 268530 243616
rect 268474 243536 268530 243545
rect 268474 243471 268530 243480
rect 268304 239958 268424 239986
rect 268200 238332 268252 238338
rect 268200 238274 268252 238280
rect 268304 238082 268332 239958
rect 268488 239766 268516 243471
rect 268476 239760 268528 239766
rect 268476 239702 268528 239708
rect 268580 238474 268608 257343
rect 268948 251174 268976 284922
rect 268672 251146 268976 251174
rect 268672 238785 268700 251146
rect 268750 247888 268806 247897
rect 268750 247823 268806 247832
rect 268764 239494 268792 247823
rect 269040 247034 269068 287642
rect 269120 265668 269172 265674
rect 269120 265610 269172 265616
rect 269132 265577 269160 265610
rect 269118 265568 269174 265577
rect 269118 265503 269174 265512
rect 269120 257440 269172 257446
rect 269118 257408 269120 257417
rect 269172 257408 269174 257417
rect 269118 257343 269174 257352
rect 269040 247006 269160 247034
rect 268842 246528 268898 246537
rect 268842 246463 268898 246472
rect 268856 240854 268884 246463
rect 268936 244996 268988 245002
rect 268936 244938 268988 244944
rect 268844 240848 268896 240854
rect 268844 240790 268896 240796
rect 268842 240680 268898 240689
rect 268842 240615 268898 240624
rect 268856 240378 268884 240615
rect 268844 240372 268896 240378
rect 268844 240314 268896 240320
rect 268752 239488 268804 239494
rect 268752 239430 268804 239436
rect 268658 238776 268714 238785
rect 268658 238711 268714 238720
rect 268568 238468 268620 238474
rect 268568 238410 268620 238416
rect 268382 238368 268438 238377
rect 268382 238303 268438 238312
rect 268476 238332 268528 238338
rect 268212 238066 268332 238082
rect 268200 238060 268332 238066
rect 268252 238054 268332 238060
rect 268200 238002 268252 238008
rect 268304 237374 268332 238054
rect 268396 237998 268424 238303
rect 268476 238274 268528 238280
rect 268384 237992 268436 237998
rect 268384 237934 268436 237940
rect 268212 237346 268332 237374
rect 268106 235104 268162 235113
rect 268106 235039 268162 235048
rect 268212 231854 268240 237346
rect 268488 237318 268516 238274
rect 268660 238060 268712 238066
rect 268660 238002 268712 238008
rect 268476 237312 268528 237318
rect 268476 237254 268528 237260
rect 268672 236774 268700 238002
rect 268948 237862 268976 244938
rect 269028 241664 269080 241670
rect 269028 241606 269080 241612
rect 268936 237856 268988 237862
rect 268936 237798 268988 237804
rect 269040 237794 269068 241606
rect 269132 240718 269160 247006
rect 269212 241120 269264 241126
rect 269212 241062 269264 241068
rect 269224 240786 269252 241062
rect 269212 240780 269264 240786
rect 269212 240722 269264 240728
rect 269120 240712 269172 240718
rect 269120 240654 269172 240660
rect 269132 238542 269160 240654
rect 269212 240576 269264 240582
rect 269316 240553 269344 318650
rect 269396 318436 269448 318442
rect 269396 318378 269448 318384
rect 269408 317626 269436 318378
rect 269396 317620 269448 317626
rect 269396 317562 269448 317568
rect 269212 240518 269264 240524
rect 269302 240544 269358 240553
rect 269224 239562 269252 240518
rect 269302 240479 269358 240488
rect 269212 239556 269264 239562
rect 269212 239498 269264 239504
rect 269408 239290 269436 317562
rect 269592 308514 269620 385591
rect 269684 313857 269712 387087
rect 269764 374332 269816 374338
rect 269764 374274 269816 374280
rect 269670 313848 269726 313857
rect 269670 313783 269726 313792
rect 269670 308816 269726 308825
rect 269670 308751 269726 308760
rect 269580 308508 269632 308514
rect 269580 308450 269632 308456
rect 269580 257372 269632 257378
rect 269580 257314 269632 257320
rect 269486 250744 269542 250753
rect 269486 250679 269542 250688
rect 269500 240854 269528 250679
rect 269592 241505 269620 257314
rect 269578 241496 269634 241505
rect 269578 241431 269634 241440
rect 269488 240848 269540 240854
rect 269488 240790 269540 240796
rect 269580 240644 269632 240650
rect 269580 240586 269632 240592
rect 269486 240272 269542 240281
rect 269486 240207 269542 240216
rect 269500 240174 269528 240207
rect 269488 240168 269540 240174
rect 269488 240110 269540 240116
rect 269488 239420 269540 239426
rect 269488 239362 269540 239368
rect 269396 239284 269448 239290
rect 269396 239226 269448 239232
rect 269120 238536 269172 238542
rect 269120 238478 269172 238484
rect 269120 238264 269172 238270
rect 269120 238206 269172 238212
rect 269028 237788 269080 237794
rect 269028 237730 269080 237736
rect 268844 237380 268896 237386
rect 268844 237322 268896 237328
rect 268660 236768 268712 236774
rect 268660 236710 268712 236716
rect 268292 235884 268344 235890
rect 268292 235826 268344 235832
rect 268304 235414 268332 235826
rect 268292 235408 268344 235414
rect 268292 235350 268344 235356
rect 268856 231854 268884 237322
rect 268934 237280 268990 237289
rect 268934 237215 268990 237224
rect 268212 231826 268332 231854
rect 268014 229936 268070 229945
rect 268014 229871 268070 229880
rect 268304 219434 268332 231826
rect 268764 231826 268884 231854
rect 268764 229094 268792 231826
rect 268948 230568 268976 237215
rect 269132 235793 269160 238206
rect 269118 235784 269174 235793
rect 269118 235719 269174 235728
rect 269500 235482 269528 239362
rect 269592 236774 269620 240586
rect 269580 236768 269632 236774
rect 269580 236710 269632 236716
rect 269578 235648 269634 235657
rect 269578 235583 269634 235592
rect 269592 235482 269620 235583
rect 269488 235476 269540 235482
rect 269488 235418 269540 235424
rect 269580 235476 269632 235482
rect 269580 235418 269632 235424
rect 269028 235136 269080 235142
rect 269028 235078 269080 235084
rect 269040 230994 269068 235078
rect 269684 233238 269712 308751
rect 269776 292194 269804 374274
rect 269868 321638 269896 392566
rect 269948 383104 270000 383110
rect 269948 383046 270000 383052
rect 269856 321632 269908 321638
rect 269856 321574 269908 321580
rect 269960 318442 269988 383046
rect 270144 320385 270172 396714
rect 270328 325694 270356 397967
rect 270406 395312 270462 395321
rect 270406 395247 270462 395256
rect 270236 325666 270356 325694
rect 270130 320376 270186 320385
rect 270130 320311 270186 320320
rect 270040 318504 270092 318510
rect 270040 318446 270092 318452
rect 269948 318436 270000 318442
rect 269948 318378 270000 318384
rect 269854 318200 269910 318209
rect 269854 318135 269910 318144
rect 269764 292188 269816 292194
rect 269764 292130 269816 292136
rect 269764 283620 269816 283626
rect 269764 283562 269816 283568
rect 269776 246673 269804 283562
rect 269762 246664 269818 246673
rect 269762 246599 269818 246608
rect 269764 246424 269816 246430
rect 269764 246366 269816 246372
rect 269776 238134 269804 246366
rect 269868 239154 269896 318135
rect 269946 245168 270002 245177
rect 269946 245103 270002 245112
rect 269960 239358 269988 245103
rect 269948 239352 270000 239358
rect 269948 239294 270000 239300
rect 270052 239222 270080 318446
rect 270144 311438 270172 320311
rect 270236 318578 270264 325666
rect 270316 321632 270368 321638
rect 270316 321574 270368 321580
rect 270224 318572 270276 318578
rect 270224 318514 270276 318520
rect 270132 311432 270184 311438
rect 270132 311374 270184 311380
rect 270130 241768 270186 241777
rect 270130 241703 270186 241712
rect 270144 240514 270172 241703
rect 270132 240508 270184 240514
rect 270132 240450 270184 240456
rect 270132 240236 270184 240242
rect 270132 240178 270184 240184
rect 270040 239216 270092 239222
rect 270040 239158 270092 239164
rect 269856 239148 269908 239154
rect 269856 239090 269908 239096
rect 269764 238128 269816 238134
rect 269764 238070 269816 238076
rect 269856 238128 269908 238134
rect 269856 238070 269908 238076
rect 269868 236570 269896 238070
rect 270144 237289 270172 240178
rect 270236 239329 270264 318514
rect 270328 318442 270356 321574
rect 270316 318436 270368 318442
rect 270316 318378 270368 318384
rect 270420 315858 270448 395247
rect 271144 385212 271196 385218
rect 271144 385154 271196 385160
rect 271052 358760 271104 358766
rect 271052 358702 271104 358708
rect 271064 357474 271092 358702
rect 271052 357468 271104 357474
rect 271052 357410 271104 357416
rect 270960 317008 271012 317014
rect 270960 316950 271012 316956
rect 270408 315852 270460 315858
rect 270408 315794 270460 315800
rect 270420 315450 270448 315794
rect 270408 315444 270460 315450
rect 270408 315386 270460 315392
rect 270408 309120 270460 309126
rect 270408 309062 270460 309068
rect 270420 308514 270448 309062
rect 270408 308508 270460 308514
rect 270408 308450 270460 308456
rect 270316 303680 270368 303686
rect 270316 303622 270368 303628
rect 270222 239320 270278 239329
rect 270222 239255 270278 239264
rect 270130 237280 270186 237289
rect 270130 237215 270186 237224
rect 269856 236564 269908 236570
rect 269856 236506 269908 236512
rect 270132 235476 270184 235482
rect 270132 235418 270184 235424
rect 269764 235204 269816 235210
rect 269764 235146 269816 235152
rect 269672 233232 269724 233238
rect 269672 233174 269724 233180
rect 269028 230988 269080 230994
rect 269028 230930 269080 230936
rect 268948 230540 269068 230568
rect 268764 229066 268976 229094
rect 268212 219406 268332 219434
rect 267922 155680 267978 155689
rect 267922 155615 267978 155624
rect 267830 155544 267886 155553
rect 267830 155479 267886 155488
rect 267922 141808 267978 141817
rect 267922 141743 267978 141752
rect 265348 141704 265400 141710
rect 265348 141646 265400 141652
rect 267004 141500 267056 141506
rect 267004 141442 267056 141448
rect 265622 97336 265678 97345
rect 265622 97271 265678 97280
rect 265348 4004 265400 4010
rect 265348 3946 265400 3952
rect 264244 3392 264296 3398
rect 264244 3334 264296 3340
rect 265360 480 265388 3946
rect 265636 3330 265664 97271
rect 267016 4146 267044 141442
rect 267936 141438 267964 141743
rect 267924 141432 267976 141438
rect 267924 141374 267976 141380
rect 268212 129742 268240 219406
rect 268948 144702 268976 229066
rect 268936 144696 268988 144702
rect 268936 144638 268988 144644
rect 268948 144226 268976 144638
rect 268936 144220 268988 144226
rect 268936 144162 268988 144168
rect 269040 139262 269068 230540
rect 269304 229900 269356 229906
rect 269304 229842 269356 229848
rect 269396 229900 269448 229906
rect 269396 229842 269448 229848
rect 269316 229702 269344 229842
rect 269304 229696 269356 229702
rect 269304 229638 269356 229644
rect 269408 229094 269436 229842
rect 269316 229066 269436 229094
rect 269316 228206 269344 229066
rect 269304 228200 269356 228206
rect 269304 228142 269356 228148
rect 269120 154148 269172 154154
rect 269120 154090 269172 154096
rect 269132 148918 269160 154090
rect 269120 148912 269172 148918
rect 269120 148854 269172 148860
rect 269316 143546 269344 228142
rect 269776 151609 269804 235146
rect 270144 233832 270172 235418
rect 270328 234433 270356 303622
rect 270500 291372 270552 291378
rect 270500 291314 270552 291320
rect 270408 253360 270460 253366
rect 270408 253302 270460 253308
rect 270420 237726 270448 253302
rect 270408 237720 270460 237726
rect 270408 237662 270460 237668
rect 270408 235408 270460 235414
rect 270408 235350 270460 235356
rect 270314 234424 270370 234433
rect 270314 234359 270370 234368
rect 270144 233804 270264 233832
rect 270132 233708 270184 233714
rect 270132 233650 270184 233656
rect 270040 232484 270092 232490
rect 270040 232426 270092 232432
rect 270052 232150 270080 232426
rect 270040 232144 270092 232150
rect 270040 232086 270092 232092
rect 270144 154154 270172 233650
rect 270132 154148 270184 154154
rect 270132 154090 270184 154096
rect 270144 153270 270172 154090
rect 270132 153264 270184 153270
rect 270132 153206 270184 153212
rect 270236 151814 270264 233804
rect 270316 233232 270368 233238
rect 270316 233174 270368 233180
rect 270052 151786 270264 151814
rect 269762 151600 269818 151609
rect 269762 151535 269818 151544
rect 269776 151201 269804 151535
rect 269762 151192 269818 151201
rect 269762 151127 269818 151136
rect 270052 148986 270080 151786
rect 270328 149138 270356 233174
rect 270236 149110 270356 149138
rect 270040 148980 270092 148986
rect 270040 148922 270092 148928
rect 270236 148186 270264 149110
rect 270316 148980 270368 148986
rect 270316 148922 270368 148928
rect 270328 148374 270356 148922
rect 270316 148368 270368 148374
rect 270316 148310 270368 148316
rect 270236 148158 270356 148186
rect 270328 146130 270356 148158
rect 270316 146124 270368 146130
rect 270316 146066 270368 146072
rect 270328 145722 270356 146066
rect 270316 145716 270368 145722
rect 270316 145658 270368 145664
rect 269212 143540 269264 143546
rect 269212 143482 269264 143488
rect 269304 143540 269356 143546
rect 269304 143482 269356 143488
rect 269764 143540 269816 143546
rect 269764 143482 269816 143488
rect 269224 142934 269252 143482
rect 269212 142928 269264 142934
rect 269212 142870 269264 142876
rect 269028 139256 269080 139262
rect 269028 139198 269080 139204
rect 269040 138718 269068 139198
rect 269028 138712 269080 138718
rect 269028 138654 269080 138660
rect 268200 129736 268252 129742
rect 268200 129678 268252 129684
rect 269028 129736 269080 129742
rect 269028 129678 269080 129684
rect 269040 129130 269068 129678
rect 269028 129124 269080 129130
rect 269028 129066 269080 129072
rect 269118 32464 269174 32473
rect 269118 32399 269174 32408
rect 269132 16574 269160 32399
rect 269132 16546 269712 16574
rect 267004 4140 267056 4146
rect 267004 4082 267056 4088
rect 267648 4072 267700 4078
rect 267700 4020 267780 4026
rect 267648 4014 267780 4020
rect 267660 3998 267780 4014
rect 265624 3324 265676 3330
rect 265624 3266 265676 3272
rect 266544 3324 266596 3330
rect 266544 3266 266596 3272
rect 266556 480 266584 3266
rect 267752 480 267780 3998
rect 268844 3936 268896 3942
rect 268844 3878 268896 3884
rect 268856 480 268884 3878
rect 269684 3482 269712 16546
rect 269776 3942 269804 143482
rect 270420 129674 270448 235350
rect 270512 228682 270540 291314
rect 270776 291304 270828 291310
rect 270776 291246 270828 291252
rect 270592 241324 270644 241330
rect 270592 241266 270644 241272
rect 270604 238649 270632 241266
rect 270684 240984 270736 240990
rect 270684 240926 270736 240932
rect 270696 240242 270724 240926
rect 270684 240236 270736 240242
rect 270684 240178 270736 240184
rect 270684 239352 270736 239358
rect 270684 239294 270736 239300
rect 270696 238678 270724 239294
rect 270684 238672 270736 238678
rect 270590 238640 270646 238649
rect 270684 238614 270736 238620
rect 270590 238575 270646 238584
rect 270604 233238 270632 238575
rect 270592 233232 270644 233238
rect 270592 233174 270644 233180
rect 270684 232484 270736 232490
rect 270684 232426 270736 232432
rect 270592 232212 270644 232218
rect 270592 232154 270644 232160
rect 270500 228676 270552 228682
rect 270500 228618 270552 228624
rect 270604 157321 270632 232154
rect 270590 157312 270646 157321
rect 270590 157247 270646 157256
rect 270696 155281 270724 232426
rect 270788 228614 270816 291246
rect 270868 245744 270920 245750
rect 270868 245686 270920 245692
rect 270880 239630 270908 245686
rect 270972 241330 271000 316950
rect 271064 291854 271092 357410
rect 271052 291848 271104 291854
rect 271052 291790 271104 291796
rect 271156 291310 271184 385154
rect 271236 382424 271288 382430
rect 271236 382366 271288 382372
rect 271248 291378 271276 382366
rect 271340 370802 271368 450774
rect 274456 400308 274508 400314
rect 274456 400250 274508 400256
rect 273168 399696 273220 399702
rect 273168 399638 273220 399644
rect 271418 395720 271474 395729
rect 271418 395655 271474 395664
rect 271328 370796 271380 370802
rect 271328 370738 271380 370744
rect 271340 370598 271368 370738
rect 271328 370592 271380 370598
rect 271328 370534 271380 370540
rect 271328 321156 271380 321162
rect 271328 321098 271380 321104
rect 271340 318102 271368 321098
rect 271432 320929 271460 395655
rect 272984 395548 273036 395554
rect 272984 395490 273036 395496
rect 271604 395480 271656 395486
rect 271604 395422 271656 395428
rect 271512 388680 271564 388686
rect 271512 388622 271564 388628
rect 271418 320920 271474 320929
rect 271418 320855 271474 320864
rect 271328 318096 271380 318102
rect 271328 318038 271380 318044
rect 271328 316124 271380 316130
rect 271328 316066 271380 316072
rect 271236 291372 271288 291378
rect 271236 291314 271288 291320
rect 271144 291304 271196 291310
rect 271144 291246 271196 291252
rect 271144 280832 271196 280838
rect 271144 280774 271196 280780
rect 271052 247920 271104 247926
rect 271052 247862 271104 247868
rect 270960 241324 271012 241330
rect 270960 241266 271012 241272
rect 270868 239624 270920 239630
rect 270868 239566 270920 239572
rect 270776 228608 270828 228614
rect 270776 228550 270828 228556
rect 270776 226364 270828 226370
rect 270776 226306 270828 226312
rect 270788 157282 270816 226306
rect 270776 157276 270828 157282
rect 270776 157218 270828 157224
rect 270682 155272 270738 155281
rect 270682 155207 270738 155216
rect 270880 136542 270908 239566
rect 271064 238513 271092 247862
rect 271156 241670 271184 280774
rect 271236 279472 271288 279478
rect 271236 279414 271288 279420
rect 271248 245002 271276 279414
rect 271236 244996 271288 245002
rect 271236 244938 271288 244944
rect 271144 241664 271196 241670
rect 271144 241606 271196 241612
rect 271144 241392 271196 241398
rect 271144 241334 271196 241340
rect 271156 240854 271184 241334
rect 271144 240848 271196 240854
rect 271144 240790 271196 240796
rect 271236 239760 271288 239766
rect 271236 239702 271288 239708
rect 271050 238504 271106 238513
rect 271050 238439 271106 238448
rect 271248 238105 271276 239702
rect 271234 238096 271290 238105
rect 271234 238031 271290 238040
rect 270958 235376 271014 235385
rect 270958 235311 271014 235320
rect 270972 232490 271000 235311
rect 270960 232484 271012 232490
rect 270960 232426 271012 232432
rect 271144 230444 271196 230450
rect 271144 230386 271196 230392
rect 271156 155106 271184 230386
rect 271340 227730 271368 316066
rect 271524 314634 271552 388622
rect 271616 321162 271644 395422
rect 271694 393952 271750 393961
rect 271694 393887 271750 393896
rect 271604 321156 271656 321162
rect 271604 321098 271656 321104
rect 271604 321020 271656 321026
rect 271604 320962 271656 320968
rect 271616 316034 271644 320962
rect 271708 320906 271736 393887
rect 271786 392592 271842 392601
rect 271786 392527 271842 392536
rect 271800 321026 271828 392527
rect 272522 388512 272578 388521
rect 272522 388447 272578 388456
rect 272340 374468 272392 374474
rect 272340 374410 272392 374416
rect 272248 322312 272300 322318
rect 272248 322254 272300 322260
rect 271788 321020 271840 321026
rect 271788 320962 271840 320968
rect 271708 320878 271828 320906
rect 271696 318368 271748 318374
rect 271696 318310 271748 318316
rect 271708 318102 271736 318310
rect 271696 318096 271748 318102
rect 271696 318038 271748 318044
rect 271616 316006 271736 316034
rect 271800 316033 271828 320878
rect 272260 316713 272288 322254
rect 272246 316704 272302 316713
rect 272246 316639 272302 316648
rect 271512 314628 271564 314634
rect 271512 314570 271564 314576
rect 271420 314084 271472 314090
rect 271420 314026 271472 314032
rect 271432 230518 271460 314026
rect 271708 313721 271736 316006
rect 271786 316024 271842 316033
rect 271786 315959 271842 315968
rect 271800 315081 271828 315959
rect 271786 315072 271842 315081
rect 271786 315007 271842 315016
rect 271694 313712 271750 313721
rect 271694 313647 271750 313656
rect 271708 313449 271736 313647
rect 271694 313440 271750 313449
rect 271694 313375 271750 313384
rect 271880 311364 271932 311370
rect 271880 311306 271932 311312
rect 271602 309632 271658 309641
rect 271602 309567 271658 309576
rect 271616 248414 271644 309567
rect 271696 297424 271748 297430
rect 271696 297366 271748 297372
rect 271524 248386 271644 248414
rect 271524 245750 271552 248386
rect 271512 245744 271564 245750
rect 271512 245686 271564 245692
rect 271604 240916 271656 240922
rect 271604 240858 271656 240864
rect 271512 239624 271564 239630
rect 271512 239566 271564 239572
rect 271524 238746 271552 239566
rect 271616 239494 271644 240858
rect 271604 239488 271656 239494
rect 271604 239430 271656 239436
rect 271512 238740 271564 238746
rect 271512 238682 271564 238688
rect 271616 232218 271644 239430
rect 271604 232212 271656 232218
rect 271604 232154 271656 232160
rect 271708 231441 271736 297366
rect 271788 243568 271840 243574
rect 271788 243510 271840 243516
rect 271800 237425 271828 243510
rect 271786 237416 271842 237425
rect 271786 237351 271842 237360
rect 271694 231432 271750 231441
rect 271694 231367 271750 231376
rect 271420 230512 271472 230518
rect 271420 230454 271472 230460
rect 271328 227724 271380 227730
rect 271328 227666 271380 227672
rect 271340 226370 271368 227666
rect 271328 226364 271380 226370
rect 271328 226306 271380 226312
rect 271892 221610 271920 311306
rect 272352 296002 272380 374410
rect 272432 372768 272484 372774
rect 272432 372710 272484 372716
rect 272340 295996 272392 296002
rect 272340 295938 272392 295944
rect 272444 294846 272472 372710
rect 272536 322182 272564 388447
rect 272798 383072 272854 383081
rect 272798 383007 272854 383016
rect 272616 381064 272668 381070
rect 272616 381006 272668 381012
rect 272524 322176 272576 322182
rect 272524 322118 272576 322124
rect 272536 321706 272564 322118
rect 272524 321700 272576 321706
rect 272524 321642 272576 321648
rect 272522 319832 272578 319841
rect 272522 319767 272578 319776
rect 272432 294840 272484 294846
rect 272432 294782 272484 294788
rect 272156 291848 272208 291854
rect 272156 291790 272208 291796
rect 272340 291848 272392 291854
rect 272340 291790 272392 291796
rect 271972 291576 272024 291582
rect 271972 291518 272024 291524
rect 271984 291242 272012 291518
rect 272064 291440 272116 291446
rect 272064 291382 272116 291388
rect 271972 291236 272024 291242
rect 271972 291178 272024 291184
rect 271984 229430 272012 291178
rect 271972 229424 272024 229430
rect 271972 229366 272024 229372
rect 271972 222828 272024 222834
rect 271972 222770 272024 222776
rect 271880 221604 271932 221610
rect 271880 221546 271932 221552
rect 271788 157276 271840 157282
rect 271788 157218 271840 157224
rect 271800 156738 271828 157218
rect 271788 156732 271840 156738
rect 271788 156674 271840 156680
rect 271144 155100 271196 155106
rect 271144 155042 271196 155048
rect 270868 136536 270920 136542
rect 270868 136478 270920 136484
rect 270408 129668 270460 129674
rect 270408 129610 270460 129616
rect 270420 129062 270448 129610
rect 270408 129056 270460 129062
rect 270408 128998 270460 129004
rect 269764 3936 269816 3942
rect 269764 3878 269816 3884
rect 269684 3454 270080 3482
rect 270052 480 270080 3454
rect 271156 3330 271184 155042
rect 271984 139330 272012 222770
rect 272076 211818 272104 291382
rect 272168 228546 272196 291790
rect 272352 291446 272380 291790
rect 272340 291440 272392 291446
rect 272340 291382 272392 291388
rect 272248 247784 272300 247790
rect 272248 247726 272300 247732
rect 272260 241058 272288 247726
rect 272248 241052 272300 241058
rect 272248 240994 272300 241000
rect 272156 228540 272208 228546
rect 272156 228482 272208 228488
rect 272064 211812 272116 211818
rect 272064 211754 272116 211760
rect 272260 158098 272288 240994
rect 272536 222834 272564 319767
rect 272628 291582 272656 381006
rect 272708 379908 272760 379914
rect 272708 379850 272760 379856
rect 272720 291650 272748 379850
rect 272812 325694 272840 383007
rect 272812 325666 272932 325694
rect 272798 321464 272854 321473
rect 272798 321399 272854 321408
rect 272812 321065 272840 321399
rect 272798 321056 272854 321065
rect 272798 320991 272854 321000
rect 272904 319530 272932 325666
rect 272996 321473 273024 395490
rect 273076 374400 273128 374406
rect 273076 374342 273128 374348
rect 272982 321464 273038 321473
rect 272982 321399 273038 321408
rect 272984 320952 273036 320958
rect 272984 320894 273036 320900
rect 272892 319524 272944 319530
rect 272892 319466 272944 319472
rect 272996 319410 273024 320894
rect 272904 319382 273024 319410
rect 272798 317112 272854 317121
rect 272798 317047 272854 317056
rect 272708 291644 272760 291650
rect 272708 291586 272760 291592
rect 272616 291576 272668 291582
rect 272616 291518 272668 291524
rect 272708 237584 272760 237590
rect 272708 237526 272760 237532
rect 272720 234598 272748 237526
rect 272708 234592 272760 234598
rect 272708 234534 272760 234540
rect 272614 231160 272670 231169
rect 272614 231095 272670 231104
rect 272524 222828 272576 222834
rect 272524 222770 272576 222776
rect 272248 158092 272300 158098
rect 272248 158034 272300 158040
rect 272628 140690 272656 231095
rect 272812 230489 272840 317047
rect 272904 233782 272932 319382
rect 272982 317248 273038 317257
rect 272982 317183 273038 317192
rect 272996 316713 273024 317183
rect 272982 316704 273038 316713
rect 272982 316639 273038 316648
rect 272982 316296 273038 316305
rect 272982 316231 273038 316240
rect 272892 233776 272944 233782
rect 272892 233718 272944 233724
rect 272798 230480 272854 230489
rect 272798 230415 272854 230424
rect 272996 229702 273024 316231
rect 273088 292058 273116 374342
rect 273180 322318 273208 399638
rect 273994 395856 274050 395865
rect 273994 395791 274050 395800
rect 273812 385688 273864 385694
rect 273812 385630 273864 385636
rect 273168 322312 273220 322318
rect 273168 322254 273220 322260
rect 273168 322176 273220 322182
rect 273168 322118 273220 322124
rect 273180 319297 273208 322118
rect 273718 321056 273774 321065
rect 273718 320991 273774 321000
rect 273166 319288 273222 319297
rect 273166 319223 273222 319232
rect 273352 310072 273404 310078
rect 273352 310014 273404 310020
rect 273076 292052 273128 292058
rect 273076 291994 273128 292000
rect 273260 239556 273312 239562
rect 273260 239498 273312 239504
rect 273272 238882 273300 239498
rect 273260 238876 273312 238882
rect 273260 238818 273312 238824
rect 273168 234592 273220 234598
rect 273168 234534 273220 234540
rect 272984 229696 273036 229702
rect 272984 229638 273036 229644
rect 273180 151745 273208 234534
rect 273166 151736 273222 151745
rect 273166 151671 273222 151680
rect 273180 151065 273208 151671
rect 273166 151056 273222 151065
rect 273166 150991 273222 151000
rect 273272 147422 273300 238818
rect 273364 219094 273392 310014
rect 273444 241052 273496 241058
rect 273444 240994 273496 241000
rect 273456 238241 273484 240994
rect 273536 238468 273588 238474
rect 273536 238410 273588 238416
rect 273442 238232 273498 238241
rect 273442 238167 273498 238176
rect 273456 230450 273484 238167
rect 273548 237998 273576 238410
rect 273536 237992 273588 237998
rect 273536 237934 273588 237940
rect 273444 230444 273496 230450
rect 273444 230386 273496 230392
rect 273444 224936 273496 224942
rect 273444 224878 273496 224884
rect 273352 219088 273404 219094
rect 273352 219030 273404 219036
rect 273260 147416 273312 147422
rect 273260 147358 273312 147364
rect 273456 142934 273484 224878
rect 273548 158953 273576 237934
rect 273732 232694 273760 320991
rect 273824 319462 273852 385630
rect 273904 372088 273956 372094
rect 273904 372030 273956 372036
rect 273916 319734 273944 372030
rect 273904 319728 273956 319734
rect 274008 319705 274036 395791
rect 274364 395344 274416 395350
rect 274364 395286 274416 395292
rect 274088 383240 274140 383246
rect 274088 383182 274140 383188
rect 273904 319670 273956 319676
rect 273994 319696 274050 319705
rect 273994 319631 274050 319640
rect 273812 319456 273864 319462
rect 273812 319398 273864 319404
rect 273824 317642 273852 319398
rect 274100 318714 274128 383182
rect 274180 376032 274232 376038
rect 274180 375974 274232 375980
rect 274088 318708 274140 318714
rect 274088 318650 274140 318656
rect 273824 317614 273944 317642
rect 273810 316160 273866 316169
rect 273810 316095 273866 316104
rect 273824 256766 273852 316095
rect 273812 256760 273864 256766
rect 273812 256702 273864 256708
rect 273720 232688 273772 232694
rect 273720 232630 273772 232636
rect 273628 232212 273680 232218
rect 273628 232154 273680 232160
rect 273640 160857 273668 232154
rect 273916 224942 273944 317614
rect 273996 315444 274048 315450
rect 273996 315386 274048 315392
rect 273904 224936 273956 224942
rect 273904 224878 273956 224884
rect 274008 224330 274036 315386
rect 274192 288425 274220 375974
rect 274272 375896 274324 375902
rect 274272 375838 274324 375844
rect 274284 288454 274312 375838
rect 274376 315994 274404 395286
rect 274468 318510 274496 400250
rect 274560 372706 274588 463694
rect 275284 461644 275336 461650
rect 275284 461586 275336 461592
rect 275296 460970 275324 461586
rect 275284 460964 275336 460970
rect 275284 460906 275336 460912
rect 275296 374746 275324 460906
rect 275926 403064 275982 403073
rect 275926 402999 275982 403008
rect 275836 400240 275888 400246
rect 275836 400182 275888 400188
rect 275558 391368 275614 391377
rect 275558 391303 275614 391312
rect 275466 382936 275522 382945
rect 275466 382871 275522 382880
rect 275376 376100 275428 376106
rect 275376 376042 275428 376048
rect 275284 374740 275336 374746
rect 275284 374682 275336 374688
rect 275192 373108 275244 373114
rect 275192 373050 275244 373056
rect 275100 372972 275152 372978
rect 275100 372914 275152 372920
rect 274548 372700 274600 372706
rect 274548 372642 274600 372648
rect 274560 365090 274588 372642
rect 274548 365084 274600 365090
rect 274548 365026 274600 365032
rect 274546 319696 274602 319705
rect 274546 319631 274602 319640
rect 274560 319161 274588 319631
rect 274546 319152 274602 319161
rect 274546 319087 274602 319096
rect 274456 318504 274508 318510
rect 274456 318446 274508 318452
rect 274548 317484 274600 317490
rect 274548 317426 274600 317432
rect 274456 317076 274508 317082
rect 274456 317018 274508 317024
rect 274364 315988 274416 315994
rect 274364 315930 274416 315936
rect 274364 307420 274416 307426
rect 274364 307362 274416 307368
rect 274272 288448 274324 288454
rect 274178 288416 274234 288425
rect 274272 288390 274324 288396
rect 274178 288351 274234 288360
rect 274272 239420 274324 239426
rect 274272 239362 274324 239368
rect 274284 237930 274312 239362
rect 274272 237924 274324 237930
rect 274272 237866 274324 237872
rect 274284 232218 274312 237866
rect 274376 235929 274404 307362
rect 274468 241058 274496 317018
rect 274560 241369 274588 317426
rect 275008 301572 275060 301578
rect 275008 301514 275060 301520
rect 274640 256760 274692 256766
rect 274640 256702 274692 256708
rect 274546 241360 274602 241369
rect 274546 241295 274602 241304
rect 274456 241052 274508 241058
rect 274456 240994 274508 241000
rect 274652 236910 274680 256702
rect 274732 240712 274784 240718
rect 274732 240654 274784 240660
rect 274640 236904 274692 236910
rect 274640 236846 274692 236852
rect 274546 236464 274602 236473
rect 274546 236399 274602 236408
rect 274560 235958 274588 236399
rect 274548 235952 274600 235958
rect 274362 235920 274418 235929
rect 274548 235894 274600 235900
rect 274362 235855 274418 235864
rect 274272 232212 274324 232218
rect 274272 232154 274324 232160
rect 274456 230444 274508 230450
rect 274456 230386 274508 230392
rect 273996 224324 274048 224330
rect 273996 224266 274048 224272
rect 273626 160848 273682 160857
rect 273626 160783 273682 160792
rect 273534 158944 273590 158953
rect 273534 158879 273590 158888
rect 274468 150278 274496 230386
rect 274456 150272 274508 150278
rect 274456 150214 274508 150220
rect 274468 149122 274496 150214
rect 274456 149116 274508 149122
rect 274456 149058 274508 149064
rect 273444 142928 273496 142934
rect 273444 142870 273496 142876
rect 272616 140684 272668 140690
rect 272616 140626 272668 140632
rect 272628 140078 272656 140626
rect 272616 140072 272668 140078
rect 272616 140014 272668 140020
rect 271972 139324 272024 139330
rect 271972 139266 272024 139272
rect 271984 138786 272012 139266
rect 271972 138780 272024 138786
rect 271972 138722 272024 138728
rect 272246 138000 272302 138009
rect 272246 137935 272302 137944
rect 272260 137902 272288 137935
rect 272248 137896 272300 137902
rect 272248 137838 272300 137844
rect 272260 136678 272288 137838
rect 272248 136672 272300 136678
rect 272248 136614 272300 136620
rect 271788 136536 271840 136542
rect 271788 136478 271840 136484
rect 271800 135930 271828 136478
rect 271788 135924 271840 135930
rect 271788 135866 271840 135872
rect 274560 128314 274588 235894
rect 274640 150136 274692 150142
rect 274640 150078 274692 150084
rect 274652 149530 274680 150078
rect 274640 149524 274692 149530
rect 274640 149466 274692 149472
rect 274088 128308 274140 128314
rect 274088 128250 274140 128256
rect 274548 128308 274600 128314
rect 274548 128250 274600 128256
rect 274100 127634 274128 128250
rect 274088 127628 274140 127634
rect 274088 127570 274140 127576
rect 273260 119400 273312 119406
rect 273260 119342 273312 119348
rect 272432 3868 272484 3874
rect 272432 3810 272484 3816
rect 271236 3392 271288 3398
rect 271236 3334 271288 3340
rect 271144 3324 271196 3330
rect 271144 3266 271196 3272
rect 271248 480 271276 3334
rect 272444 480 272472 3810
rect 262926 354 263038 480
rect 262508 326 263038 354
rect 262926 -960 263038 326
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273272 354 273300 119342
rect 274652 4010 274680 149466
rect 274744 125594 274772 240654
rect 274824 237040 274876 237046
rect 274824 236982 274876 236988
rect 274836 139398 274864 236982
rect 274916 231804 274968 231810
rect 274916 231746 274968 231752
rect 274928 150142 274956 231746
rect 275020 220454 275048 301514
rect 275112 294642 275140 372914
rect 275100 294636 275152 294642
rect 275100 294578 275152 294584
rect 275204 293418 275232 373050
rect 275282 320240 275338 320249
rect 275282 320175 275338 320184
rect 275192 293412 275244 293418
rect 275192 293354 275244 293360
rect 275296 232150 275324 320175
rect 275388 291718 275416 376042
rect 275480 320657 275508 382871
rect 275572 320793 275600 391303
rect 275652 375964 275704 375970
rect 275652 375906 275704 375912
rect 275558 320784 275614 320793
rect 275558 320719 275614 320728
rect 275466 320648 275522 320657
rect 275466 320583 275522 320592
rect 275480 320249 275508 320583
rect 275572 320521 275600 320719
rect 275558 320512 275614 320521
rect 275558 320447 275614 320456
rect 275466 320240 275522 320249
rect 275466 320175 275522 320184
rect 275560 318844 275612 318850
rect 275560 318786 275612 318792
rect 275468 317756 275520 317762
rect 275468 317698 275520 317704
rect 275376 291712 275428 291718
rect 275376 291654 275428 291660
rect 275376 261520 275428 261526
rect 275376 261462 275428 261468
rect 275388 237046 275416 261462
rect 275376 237040 275428 237046
rect 275376 236982 275428 236988
rect 275374 235920 275430 235929
rect 275374 235855 275430 235864
rect 275284 232144 275336 232150
rect 275284 232086 275336 232092
rect 275008 220448 275060 220454
rect 275008 220390 275060 220396
rect 275296 219434 275324 232086
rect 275112 219406 275324 219434
rect 275112 171134 275140 219406
rect 275112 171106 275232 171134
rect 275204 150210 275232 171106
rect 275192 150204 275244 150210
rect 275192 150146 275244 150152
rect 274916 150136 274968 150142
rect 274916 150078 274968 150084
rect 275204 149802 275232 150146
rect 275192 149796 275244 149802
rect 275192 149738 275244 149744
rect 275100 149116 275152 149122
rect 275100 149058 275152 149064
rect 275112 142154 275140 149058
rect 275190 149016 275246 149025
rect 275388 149002 275416 235855
rect 275480 231470 275508 317698
rect 275572 234190 275600 318786
rect 275664 291922 275692 375906
rect 275744 372904 275796 372910
rect 275744 372846 275796 372852
rect 275756 292466 275784 372846
rect 275848 318034 275876 400182
rect 275940 319122 275968 402999
rect 276848 399016 276900 399022
rect 276848 398958 276900 398964
rect 276756 398948 276808 398954
rect 276756 398890 276808 398896
rect 276664 385824 276716 385830
rect 276664 385766 276716 385772
rect 276572 370592 276624 370598
rect 276572 370534 276624 370540
rect 276018 369472 276074 369481
rect 276018 369407 276074 369416
rect 276032 368665 276060 369407
rect 276018 368656 276074 368665
rect 276018 368591 276074 368600
rect 276386 368656 276442 368665
rect 276386 368591 276442 368600
rect 275928 319116 275980 319122
rect 275928 319058 275980 319064
rect 275836 318028 275888 318034
rect 275836 317970 275888 317976
rect 275848 317506 275876 317970
rect 275848 317478 276060 317506
rect 275836 313472 275888 313478
rect 275836 313414 275888 313420
rect 275848 301345 275876 313414
rect 275928 307352 275980 307358
rect 275928 307294 275980 307300
rect 275834 301336 275890 301345
rect 275834 301271 275890 301280
rect 275744 292460 275796 292466
rect 275744 292402 275796 292408
rect 275652 291916 275704 291922
rect 275652 291858 275704 291864
rect 275744 247852 275796 247858
rect 275744 247794 275796 247800
rect 275652 236904 275704 236910
rect 275652 236846 275704 236852
rect 275560 234184 275612 234190
rect 275560 234126 275612 234132
rect 275468 231464 275520 231470
rect 275468 231406 275520 231412
rect 275480 230450 275508 231406
rect 275468 230444 275520 230450
rect 275468 230386 275520 230392
rect 275664 154630 275692 236846
rect 275756 231810 275784 247794
rect 275940 237386 275968 307294
rect 275928 237380 275980 237386
rect 275928 237322 275980 237328
rect 275940 237182 275968 237322
rect 275928 237176 275980 237182
rect 275928 237118 275980 237124
rect 276032 235822 276060 317478
rect 276204 242344 276256 242350
rect 276204 242286 276256 242292
rect 276216 236162 276244 242286
rect 276296 237380 276348 237386
rect 276296 237322 276348 237328
rect 276204 236156 276256 236162
rect 276204 236098 276256 236104
rect 276020 235816 276072 235822
rect 276020 235758 276072 235764
rect 276020 232756 276072 232762
rect 276020 232698 276072 232704
rect 276032 232558 276060 232698
rect 276020 232552 276072 232558
rect 276020 232494 276072 232500
rect 275744 231804 275796 231810
rect 275744 231746 275796 231752
rect 276112 231804 276164 231810
rect 276112 231746 276164 231752
rect 276124 231266 276152 231746
rect 276112 231260 276164 231266
rect 276112 231202 276164 231208
rect 275652 154624 275704 154630
rect 275652 154566 275704 154572
rect 275664 150249 275692 154566
rect 275650 150240 275706 150249
rect 275650 150175 275706 150184
rect 275246 148974 275416 149002
rect 275190 148951 275246 148960
rect 275204 148345 275232 148951
rect 275190 148336 275246 148345
rect 275190 148271 275246 148280
rect 276124 147558 276152 231202
rect 276216 158817 276244 236098
rect 276202 158808 276258 158817
rect 276202 158743 276258 158752
rect 276308 153678 276336 237322
rect 276400 233238 276428 368591
rect 276584 319598 276612 370534
rect 276572 319592 276624 319598
rect 276572 319534 276624 319540
rect 276480 319252 276532 319258
rect 276480 319194 276532 319200
rect 276492 234258 276520 319194
rect 276584 317642 276612 319534
rect 276676 317762 276704 385766
rect 276768 321094 276796 398890
rect 276756 321088 276808 321094
rect 276756 321030 276808 321036
rect 276860 320482 276888 398958
rect 276940 398200 276992 398206
rect 276940 398142 276992 398148
rect 276848 320476 276900 320482
rect 276848 320418 276900 320424
rect 276860 318850 276888 320418
rect 276848 318844 276900 318850
rect 276848 318786 276900 318792
rect 276952 318646 276980 398142
rect 277122 395584 277178 395593
rect 277122 395519 277178 395528
rect 277032 392012 277084 392018
rect 277032 391954 277084 391960
rect 276940 318640 276992 318646
rect 276940 318582 276992 318588
rect 276664 317756 276716 317762
rect 276664 317698 276716 317704
rect 276584 317614 276888 317642
rect 276756 316192 276808 316198
rect 276756 316134 276808 316140
rect 276664 315512 276716 315518
rect 276664 315454 276716 315460
rect 276480 234252 276532 234258
rect 276480 234194 276532 234200
rect 276388 233232 276440 233238
rect 276388 233174 276440 233180
rect 276676 222970 276704 315454
rect 276768 229906 276796 316134
rect 276860 232694 276888 317614
rect 276952 317490 276980 318582
rect 276940 317484 276992 317490
rect 276940 317426 276992 317432
rect 276938 316432 276994 316441
rect 276938 316367 276994 316376
rect 276848 232688 276900 232694
rect 276848 232630 276900 232636
rect 276952 231810 276980 316367
rect 277044 313206 277072 391954
rect 277136 314498 277164 395519
rect 277320 374542 277348 465054
rect 278596 454980 278648 454986
rect 278596 454922 278648 454928
rect 278504 397656 278556 397662
rect 278504 397598 278556 397604
rect 278412 387252 278464 387258
rect 278412 387194 278464 387200
rect 277768 383172 277820 383178
rect 277768 383114 277820 383120
rect 277308 374536 277360 374542
rect 277308 374478 277360 374484
rect 277216 372836 277268 372842
rect 277216 372778 277268 372784
rect 277124 314492 277176 314498
rect 277124 314434 277176 314440
rect 277032 313200 277084 313206
rect 277032 313142 277084 313148
rect 277124 308848 277176 308854
rect 277124 308790 277176 308796
rect 277032 232756 277084 232762
rect 277032 232698 277084 232704
rect 276940 231804 276992 231810
rect 276940 231746 276992 231752
rect 276756 229900 276808 229906
rect 276756 229842 276808 229848
rect 276664 222964 276716 222970
rect 276664 222906 276716 222912
rect 277044 155145 277072 232698
rect 277136 224126 277164 308790
rect 277228 290698 277256 372778
rect 277320 363662 277348 374478
rect 277308 363656 277360 363662
rect 277308 363598 277360 363604
rect 277674 358864 277730 358873
rect 277674 358799 277676 358808
rect 277728 358799 277730 358808
rect 277676 358770 277728 358776
rect 277676 318844 277728 318850
rect 277676 318786 277728 318792
rect 277216 290692 277268 290698
rect 277216 290634 277268 290640
rect 277400 241528 277452 241534
rect 277400 241470 277452 241476
rect 277412 235346 277440 241470
rect 277490 240272 277546 240281
rect 277490 240207 277546 240216
rect 277400 235340 277452 235346
rect 277400 235282 277452 235288
rect 277124 224120 277176 224126
rect 277124 224062 277176 224068
rect 277030 155136 277086 155145
rect 277030 155071 277086 155080
rect 277412 154426 277440 235282
rect 277504 160721 277532 240207
rect 277688 232898 277716 318786
rect 277780 314401 277808 383114
rect 277860 374264 277912 374270
rect 277860 374206 277912 374212
rect 277872 358766 277900 374206
rect 278136 373176 278188 373182
rect 278136 373118 278188 373124
rect 278044 372292 278096 372298
rect 278044 372234 278096 372240
rect 277952 371476 278004 371482
rect 277952 371418 278004 371424
rect 277860 358760 277912 358766
rect 277860 358702 277912 358708
rect 277964 327758 277992 371418
rect 277952 327752 278004 327758
rect 277952 327694 278004 327700
rect 278056 322250 278084 372234
rect 278044 322244 278096 322250
rect 278044 322186 278096 322192
rect 278042 321464 278098 321473
rect 278042 321399 278098 321408
rect 278056 320657 278084 321399
rect 278042 320648 278098 320657
rect 278042 320583 278098 320592
rect 278044 319932 278096 319938
rect 278044 319874 278096 319880
rect 278056 318918 278084 319874
rect 278044 318912 278096 318918
rect 278044 318854 278096 318860
rect 278044 318572 278096 318578
rect 278044 318514 278096 318520
rect 278056 318306 278084 318514
rect 278044 318300 278096 318306
rect 278044 318242 278096 318248
rect 278042 315208 278098 315217
rect 278042 315143 278098 315152
rect 277766 314392 277822 314401
rect 277766 314327 277822 314336
rect 277952 312724 278004 312730
rect 277952 312666 278004 312672
rect 277860 242208 277912 242214
rect 277860 242150 277912 242156
rect 277872 240281 277900 242150
rect 277858 240272 277914 240281
rect 277858 240207 277914 240216
rect 277964 236337 277992 312666
rect 277950 236328 278006 236337
rect 277950 236263 278006 236272
rect 277676 232892 277728 232898
rect 277676 232834 277728 232840
rect 278056 222873 278084 315143
rect 278148 293282 278176 373118
rect 278228 372632 278280 372638
rect 278228 372574 278280 372580
rect 278240 293350 278268 372574
rect 278320 370456 278372 370462
rect 278320 370398 278372 370404
rect 278332 321065 278360 370398
rect 278318 321056 278374 321065
rect 278318 320991 278374 321000
rect 278320 319184 278372 319190
rect 278320 319126 278372 319132
rect 278228 293344 278280 293350
rect 278228 293286 278280 293292
rect 278136 293276 278188 293282
rect 278136 293218 278188 293224
rect 278136 240916 278188 240922
rect 278136 240858 278188 240864
rect 278148 240242 278176 240858
rect 278136 240236 278188 240242
rect 278136 240178 278188 240184
rect 278148 238762 278176 240178
rect 278148 238734 278268 238762
rect 278136 238604 278188 238610
rect 278136 238546 278188 238552
rect 278042 222864 278098 222873
rect 278042 222799 278098 222808
rect 277490 160712 277546 160721
rect 277490 160647 277546 160656
rect 277400 154420 277452 154426
rect 277400 154362 277452 154368
rect 276296 153672 276348 153678
rect 276296 153614 276348 153620
rect 276112 147552 276164 147558
rect 276112 147494 276164 147500
rect 276308 142154 276336 153614
rect 278044 148708 278096 148714
rect 278044 148650 278096 148656
rect 276388 147552 276440 147558
rect 276388 147494 276440 147500
rect 276400 147082 276428 147494
rect 276388 147076 276440 147082
rect 276388 147018 276440 147024
rect 275112 142126 275324 142154
rect 274824 139392 274876 139398
rect 274824 139334 274876 139340
rect 274732 125588 274784 125594
rect 274732 125530 274784 125536
rect 274640 4004 274692 4010
rect 274640 3946 274692 3952
rect 275296 3398 275324 142126
rect 276032 142126 276336 142154
rect 275376 139392 275428 139398
rect 275376 139334 275428 139340
rect 275388 138854 275416 139334
rect 275376 138848 275428 138854
rect 275376 138790 275428 138796
rect 275376 125588 275428 125594
rect 275376 125530 275428 125536
rect 275388 124914 275416 125530
rect 275376 124908 275428 124914
rect 275376 124850 275428 124856
rect 275284 3392 275336 3398
rect 275284 3334 275336 3340
rect 274824 3324 274876 3330
rect 274824 3266 274876 3272
rect 274836 480 274864 3266
rect 276032 480 276060 142126
rect 276110 109712 276166 109721
rect 276110 109647 276166 109656
rect 276124 16574 276152 109647
rect 276124 16546 276704 16574
rect 273598 354 273710 480
rect 273272 326 273710 354
rect 273598 -960 273710 326
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 276676 354 276704 16546
rect 278056 3058 278084 148650
rect 278148 141982 278176 238546
rect 278240 144838 278268 238734
rect 278332 229838 278360 319126
rect 278424 314634 278452 387194
rect 278516 320142 278544 397598
rect 278608 371142 278636 454922
rect 278688 454844 278740 454850
rect 278688 454786 278740 454792
rect 278596 371136 278648 371142
rect 278596 371078 278648 371084
rect 278608 370666 278636 371078
rect 278700 371074 278728 454786
rect 281264 452192 281316 452198
rect 281264 452134 281316 452140
rect 279884 451988 279936 451994
rect 279884 451930 279936 451936
rect 279608 388748 279660 388754
rect 279608 388690 279660 388696
rect 279146 384296 279202 384305
rect 279146 384231 279202 384240
rect 279056 373040 279108 373046
rect 279056 372982 279108 372988
rect 278688 371068 278740 371074
rect 278688 371010 278740 371016
rect 278596 370660 278648 370666
rect 278596 370602 278648 370608
rect 278504 320136 278556 320142
rect 278504 320078 278556 320084
rect 278516 318850 278544 320078
rect 278504 318844 278556 318850
rect 278504 318786 278556 318792
rect 278688 317280 278740 317286
rect 278688 317222 278740 317228
rect 278504 315240 278556 315246
rect 278504 315182 278556 315188
rect 278412 314628 278464 314634
rect 278412 314570 278464 314576
rect 278516 233714 278544 315182
rect 278596 311908 278648 311914
rect 278596 311850 278648 311856
rect 278608 235210 278636 311850
rect 278700 239698 278728 317222
rect 278780 315920 278832 315926
rect 278780 315862 278832 315868
rect 278792 315314 278820 315862
rect 278780 315308 278832 315314
rect 278780 315250 278832 315256
rect 278872 313200 278924 313206
rect 278872 313142 278924 313148
rect 278884 312050 278912 313142
rect 278872 312044 278924 312050
rect 278872 311986 278924 311992
rect 278780 242276 278832 242282
rect 278780 242218 278832 242224
rect 278792 240582 278820 242218
rect 278780 240576 278832 240582
rect 278780 240518 278832 240524
rect 278688 239692 278740 239698
rect 278688 239634 278740 239640
rect 278596 235204 278648 235210
rect 278596 235146 278648 235152
rect 278780 233912 278832 233918
rect 278780 233854 278832 233860
rect 278504 233708 278556 233714
rect 278504 233650 278556 233656
rect 278320 229832 278372 229838
rect 278320 229774 278372 229780
rect 278228 144832 278280 144838
rect 278228 144774 278280 144780
rect 278136 141976 278188 141982
rect 278136 141918 278188 141924
rect 278148 141438 278176 141918
rect 278136 141432 278188 141438
rect 278136 141374 278188 141380
rect 278792 16574 278820 233854
rect 278884 228313 278912 311986
rect 279068 291174 279096 372982
rect 279160 315926 279188 384231
rect 279240 371408 279292 371414
rect 279240 371350 279292 371356
rect 279252 355366 279280 371350
rect 279516 371340 279568 371346
rect 279516 371282 279568 371288
rect 279332 371272 279384 371278
rect 279332 371214 279384 371220
rect 279240 355360 279292 355366
rect 279240 355302 279292 355308
rect 279344 351218 279372 371214
rect 279424 358828 279476 358834
rect 279424 358770 279476 358776
rect 279332 351212 279384 351218
rect 279332 351154 279384 351160
rect 279148 315920 279200 315926
rect 279148 315862 279200 315868
rect 279332 303136 279384 303142
rect 279332 303078 279384 303084
rect 279056 291168 279108 291174
rect 279056 291110 279108 291116
rect 278964 240576 279016 240582
rect 278964 240518 279016 240524
rect 278870 228304 278926 228313
rect 278870 228239 278926 228248
rect 278976 159089 279004 240518
rect 279344 234122 279372 303078
rect 279332 234116 279384 234122
rect 279332 234058 279384 234064
rect 278962 159080 279018 159089
rect 278962 159015 279018 159024
rect 279436 113150 279464 358770
rect 279528 324970 279556 371282
rect 279516 324964 279568 324970
rect 279516 324906 279568 324912
rect 279620 320113 279648 388690
rect 279700 375828 279752 375834
rect 279700 375770 279752 375776
rect 279606 320104 279662 320113
rect 279606 320039 279662 320048
rect 279516 318912 279568 318918
rect 279516 318854 279568 318860
rect 279528 232286 279556 318854
rect 279606 317928 279662 317937
rect 279606 317863 279662 317872
rect 279620 232762 279648 317863
rect 279712 292126 279740 375770
rect 279896 372026 279924 451930
rect 280710 451480 280766 451489
rect 280710 451415 280766 451424
rect 280066 401840 280122 401849
rect 280066 401775 280122 401784
rect 279976 400376 280028 400382
rect 279976 400318 280028 400324
rect 279884 372020 279936 372026
rect 279884 371962 279936 371968
rect 279896 371482 279924 371962
rect 279884 371476 279936 371482
rect 279884 371418 279936 371424
rect 279884 370252 279936 370258
rect 279884 370194 279936 370200
rect 279896 367062 279924 370194
rect 279884 367056 279936 367062
rect 279884 366998 279936 367004
rect 279988 320006 280016 400318
rect 279976 320000 280028 320006
rect 279976 319942 280028 319948
rect 279988 319258 280016 319942
rect 280080 319666 280108 401775
rect 280160 373992 280212 373998
rect 280160 373934 280212 373940
rect 280172 372162 280200 373934
rect 280160 372156 280212 372162
rect 280160 372098 280212 372104
rect 280172 365022 280200 372098
rect 280724 371686 280752 451415
rect 281078 449168 281134 449177
rect 281078 449103 281134 449112
rect 280988 392692 281040 392698
rect 280988 392634 281040 392640
rect 280896 385756 280948 385762
rect 280896 385698 280948 385704
rect 280804 382968 280856 382974
rect 280804 382910 280856 382916
rect 280712 371680 280764 371686
rect 280710 371648 280712 371657
rect 280764 371648 280766 371657
rect 280710 371583 280766 371592
rect 280620 371544 280672 371550
rect 280620 371486 280672 371492
rect 280434 369744 280490 369753
rect 280434 369679 280490 369688
rect 280448 369345 280476 369679
rect 280434 369336 280490 369345
rect 280434 369271 280490 369280
rect 280160 365016 280212 365022
rect 280160 364958 280212 364964
rect 280068 319660 280120 319666
rect 280068 319602 280120 319608
rect 279976 319252 280028 319258
rect 279976 319194 280028 319200
rect 280080 319190 280108 319602
rect 280068 319184 280120 319190
rect 280068 319126 280120 319132
rect 279792 318844 279844 318850
rect 279792 318786 279844 318792
rect 279700 292120 279752 292126
rect 279700 292062 279752 292068
rect 279804 237017 279832 318786
rect 280160 317416 280212 317422
rect 280160 317358 280212 317364
rect 280172 316946 280200 317358
rect 280160 316940 280212 316946
rect 280160 316882 280212 316888
rect 280160 314492 280212 314498
rect 280160 314434 280212 314440
rect 280172 314226 280200 314434
rect 280160 314220 280212 314226
rect 280160 314162 280212 314168
rect 279976 310072 280028 310078
rect 279976 310014 280028 310020
rect 279790 237008 279846 237017
rect 279790 236943 279846 236952
rect 279988 235686 280016 310014
rect 280068 306400 280120 306406
rect 280068 306342 280120 306348
rect 279976 235680 280028 235686
rect 279976 235622 280028 235628
rect 280080 233918 280108 306342
rect 280068 233912 280120 233918
rect 280068 233854 280120 233860
rect 279608 232756 279660 232762
rect 279608 232698 279660 232704
rect 279700 232620 279752 232626
rect 279700 232562 279752 232568
rect 279516 232280 279568 232286
rect 279516 232222 279568 232228
rect 279712 151094 279740 232562
rect 280172 221921 280200 314162
rect 280252 232552 280304 232558
rect 280252 232494 280304 232500
rect 280264 231402 280292 232494
rect 280252 231396 280304 231402
rect 280252 231338 280304 231344
rect 280158 221912 280214 221921
rect 280158 221847 280214 221856
rect 279700 151088 279752 151094
rect 279700 151030 279752 151036
rect 279712 150890 279740 151030
rect 279700 150884 279752 150890
rect 279700 150826 279752 150832
rect 280264 144770 280292 231338
rect 280448 153202 280476 369271
rect 280632 360874 280660 371486
rect 280712 371476 280764 371482
rect 280712 371418 280764 371424
rect 280620 360868 280672 360874
rect 280620 360810 280672 360816
rect 280724 359514 280752 371418
rect 280712 359508 280764 359514
rect 280712 359450 280764 359456
rect 280710 356824 280766 356833
rect 280710 356759 280766 356768
rect 280724 356726 280752 356759
rect 280712 356720 280764 356726
rect 280712 356662 280764 356668
rect 280710 345808 280766 345817
rect 280710 345743 280766 345752
rect 280724 345710 280752 345743
rect 280712 345704 280764 345710
rect 280712 345646 280764 345652
rect 280816 328454 280844 382910
rect 280724 328426 280844 328454
rect 280724 319841 280752 328426
rect 280710 319832 280766 319841
rect 280710 319767 280766 319776
rect 280908 318794 280936 385698
rect 280724 318766 280936 318794
rect 280724 317937 280752 318766
rect 280710 317928 280766 317937
rect 280710 317863 280766 317872
rect 281000 317422 281028 392634
rect 281092 371958 281120 449103
rect 281172 448588 281224 448594
rect 281172 448530 281224 448536
rect 281184 372201 281212 448530
rect 281276 373318 281304 452134
rect 281540 448656 281592 448662
rect 281540 448598 281592 448604
rect 282828 448656 282880 448662
rect 282828 448598 282880 448604
rect 281552 404326 281580 448598
rect 281540 404320 281592 404326
rect 281540 404262 281592 404268
rect 282000 404320 282052 404326
rect 282000 404262 282052 404268
rect 282012 403646 282040 404262
rect 282000 403640 282052 403646
rect 282000 403582 282052 403588
rect 282092 400444 282144 400450
rect 282092 400386 282144 400392
rect 281448 399492 281500 399498
rect 281448 399434 281500 399440
rect 281356 399084 281408 399090
rect 281356 399026 281408 399032
rect 281264 373312 281316 373318
rect 281264 373254 281316 373260
rect 281170 372192 281226 372201
rect 281170 372127 281226 372136
rect 281080 371952 281132 371958
rect 281080 371894 281132 371900
rect 281184 371890 281212 372127
rect 281172 371884 281224 371890
rect 281172 371826 281224 371832
rect 281264 371612 281316 371618
rect 281264 371554 281316 371560
rect 281080 370116 281132 370122
rect 281080 370058 281132 370064
rect 281092 345817 281120 370058
rect 281276 356833 281304 371554
rect 281262 356824 281318 356833
rect 281262 356759 281318 356768
rect 281078 345808 281134 345817
rect 281078 345743 281134 345752
rect 281368 345014 281396 399026
rect 281460 372065 281488 399434
rect 281540 396840 281592 396846
rect 281540 396782 281592 396788
rect 281446 372056 281502 372065
rect 281446 371991 281502 372000
rect 281460 369170 281488 371991
rect 281448 369164 281500 369170
rect 281448 369106 281500 369112
rect 281368 344986 281488 345014
rect 281460 318850 281488 344986
rect 281448 318844 281500 318850
rect 281448 318786 281500 318792
rect 281552 318238 281580 396782
rect 281632 395140 281684 395146
rect 281632 395082 281684 395088
rect 281644 320618 281672 395082
rect 281724 389904 281776 389910
rect 281724 389846 281776 389852
rect 281632 320612 281684 320618
rect 281632 320554 281684 320560
rect 281630 320512 281686 320521
rect 281630 320447 281686 320456
rect 281540 318232 281592 318238
rect 281540 318174 281592 318180
rect 281644 318170 281672 320447
rect 281736 320249 281764 389846
rect 281816 380248 281868 380254
rect 281816 380190 281868 380196
rect 281722 320240 281778 320249
rect 281722 320175 281778 320184
rect 281736 319433 281764 320175
rect 281828 319569 281856 380190
rect 281908 377460 281960 377466
rect 281908 377402 281960 377408
rect 281920 319802 281948 377402
rect 281998 319832 282054 319841
rect 281908 319796 281960 319802
rect 281998 319767 282054 319776
rect 281908 319738 281960 319744
rect 281814 319560 281870 319569
rect 281814 319495 281870 319504
rect 281722 319424 281778 319433
rect 281722 319359 281778 319368
rect 281906 319424 281962 319433
rect 281906 319359 281962 319368
rect 281920 318850 281948 319359
rect 282012 319025 282040 319767
rect 281998 319016 282054 319025
rect 281998 318951 282054 318960
rect 281908 318844 281960 318850
rect 281908 318786 281960 318792
rect 282104 318782 282132 400386
rect 282736 385960 282788 385966
rect 282736 385902 282788 385908
rect 282276 373924 282328 373930
rect 282276 373866 282328 373872
rect 282288 371929 282316 373866
rect 282748 372094 282776 385902
rect 282840 374678 282868 448598
rect 282932 409222 282960 702406
rect 298744 501016 298796 501022
rect 298744 500958 298796 500964
rect 289820 454572 289872 454578
rect 289820 454514 289872 454520
rect 286322 449032 286378 449041
rect 286322 448967 286378 448976
rect 284482 444952 284538 444961
rect 284482 444887 284538 444896
rect 282920 409216 282972 409222
rect 282920 409158 282972 409164
rect 282920 398268 282972 398274
rect 282920 398210 282972 398216
rect 282932 395146 282960 398210
rect 282920 395140 282972 395146
rect 282920 395082 282972 395088
rect 282828 374672 282880 374678
rect 282828 374614 282880 374620
rect 282840 373994 282868 374614
rect 282840 373966 282960 373994
rect 282932 372094 282960 373966
rect 282736 372088 282788 372094
rect 282736 372030 282788 372036
rect 282920 372088 282972 372094
rect 282920 372030 282972 372036
rect 282274 371920 282330 371929
rect 282748 371890 282776 372030
rect 282274 371855 282330 371864
rect 282736 371884 282788 371890
rect 282736 371826 282788 371832
rect 283656 371884 283708 371890
rect 283656 371826 283708 371832
rect 282276 371816 282328 371822
rect 282276 371758 282328 371764
rect 282184 371748 282236 371754
rect 282184 371690 282236 371696
rect 282196 353977 282224 371690
rect 282288 360913 282316 371758
rect 283668 369866 283696 371826
rect 284496 370025 284524 444887
rect 284944 428460 284996 428466
rect 284944 428402 284996 428408
rect 284956 383654 284984 428402
rect 285034 401976 285090 401985
rect 285034 401911 285090 401920
rect 284588 383626 284984 383654
rect 284588 372881 284616 383626
rect 285048 379514 285076 401911
rect 285126 392728 285182 392737
rect 285126 392663 285182 392672
rect 284956 379486 285076 379514
rect 284574 372872 284630 372881
rect 284574 372807 284630 372816
rect 284482 370016 284538 370025
rect 284482 369951 284538 369960
rect 284588 369866 284616 372807
rect 284956 370161 284984 379486
rect 285140 370462 285168 392663
rect 286336 383654 286364 448967
rect 289728 438184 289780 438190
rect 289728 438126 289780 438132
rect 288348 424380 288400 424386
rect 288348 424322 288400 424328
rect 286336 383626 286732 383654
rect 286704 373017 286732 383626
rect 288360 379514 288388 424322
rect 289740 379514 289768 438126
rect 289832 383654 289860 454514
rect 294604 453552 294656 453558
rect 294604 453494 294656 453500
rect 291844 451920 291896 451926
rect 291844 451862 291896 451868
rect 289832 383626 290136 383654
rect 288268 379486 288388 379514
rect 289648 379486 289768 379514
rect 287428 373312 287480 373318
rect 287428 373254 287480 373260
rect 286690 373008 286746 373017
rect 286690 372943 286746 372952
rect 286046 372736 286102 372745
rect 286046 372671 286102 372680
rect 285220 371680 285272 371686
rect 285220 371622 285272 371628
rect 285128 370456 285180 370462
rect 285128 370398 285180 370404
rect 284942 370152 284998 370161
rect 284942 370087 284998 370096
rect 284850 370016 284906 370025
rect 284850 369951 284906 369960
rect 283668 369838 284004 369866
rect 284372 369838 284616 369866
rect 284864 369730 284892 369951
rect 284740 369702 284892 369730
rect 284956 369594 284984 370087
rect 285232 369866 285260 371622
rect 286060 370161 286088 372671
rect 286324 371952 286376 371958
rect 286324 371894 286376 371900
rect 286046 370152 286102 370161
rect 286046 370087 286102 370096
rect 285232 369838 285476 369866
rect 286060 369854 286088 370087
rect 286336 369866 286364 371894
rect 286704 369866 286732 372943
rect 287152 371272 287204 371278
rect 287152 371214 287204 371220
rect 286060 369826 286226 369854
rect 286336 369838 286580 369866
rect 286704 369838 286948 369866
rect 285080 369608 285136 369617
rect 284956 369566 285080 369594
rect 287164 369594 287192 371214
rect 287440 369866 287468 373254
rect 288268 372298 288296 379486
rect 288256 372292 288308 372298
rect 288256 372234 288308 372240
rect 288268 372162 288296 372234
rect 287704 372156 287756 372162
rect 287704 372098 287756 372104
rect 288256 372156 288308 372162
rect 288256 372098 288308 372104
rect 287612 371884 287664 371890
rect 287612 371826 287664 371832
rect 287624 371346 287652 371826
rect 287716 371686 287744 372098
rect 287704 371680 287756 371686
rect 287704 371622 287756 371628
rect 287612 371340 287664 371346
rect 287612 371282 287664 371288
rect 288268 369866 288296 372098
rect 288532 372088 288584 372094
rect 288532 372030 288584 372036
rect 288348 371340 288400 371346
rect 288348 371282 288400 371288
rect 288360 371074 288388 371282
rect 288348 371068 288400 371074
rect 288348 371010 288400 371016
rect 288544 369866 288572 372030
rect 289648 371521 289676 379486
rect 290002 372192 290058 372201
rect 290002 372127 290058 372136
rect 289634 371512 289690 371521
rect 289634 371447 289690 371456
rect 289358 370696 289414 370705
rect 289358 370631 289414 370640
rect 289372 369866 289400 370631
rect 289648 369866 289676 371447
rect 289728 371272 289780 371278
rect 289728 371214 289780 371220
rect 289740 371142 289768 371214
rect 289728 371136 289780 371142
rect 289728 371078 289780 371084
rect 287440 369838 287684 369866
rect 288268 369838 288420 369866
rect 288544 369838 288788 369866
rect 289004 369838 289400 369866
rect 289524 369838 289676 369866
rect 288024 369744 288080 369753
rect 288024 369679 288080 369688
rect 287288 369608 287344 369617
rect 287164 369566 287288 369594
rect 285080 369543 285136 369552
rect 287288 369543 287344 369552
rect 289004 369442 289032 369838
rect 290016 369730 290044 372127
rect 289892 369702 290044 369730
rect 290108 369866 290136 383626
rect 291292 376168 291344 376174
rect 291292 376110 291344 376116
rect 291304 375630 291332 376110
rect 291292 375624 291344 375630
rect 291292 375566 291344 375572
rect 291856 372337 291884 451862
rect 291934 439512 291990 439521
rect 291934 439447 291990 439456
rect 291948 376174 291976 439447
rect 293224 409148 293276 409154
rect 293224 409090 293276 409096
rect 292028 406428 292080 406434
rect 292028 406370 292080 406376
rect 292040 383654 292068 406370
rect 292040 383626 292252 383654
rect 291936 376168 291988 376174
rect 291936 376110 291988 376116
rect 292224 376038 292252 383626
rect 293236 376754 293264 409090
rect 293314 400888 293370 400897
rect 293314 400823 293370 400832
rect 293052 376726 293264 376754
rect 292304 376168 292356 376174
rect 292304 376110 292356 376116
rect 292212 376032 292264 376038
rect 292212 375974 292264 375980
rect 290646 372328 290702 372337
rect 290646 372263 290702 372272
rect 291842 372328 291898 372337
rect 291842 372263 291898 372272
rect 290660 371385 290688 372263
rect 290646 371376 290702 371385
rect 290646 371311 290702 371320
rect 291844 371340 291896 371346
rect 290660 370138 290688 371311
rect 291844 371282 291896 371288
rect 290740 371272 290792 371278
rect 290740 371214 290792 371220
rect 290614 370110 290688 370138
rect 290108 369838 290260 369866
rect 290614 369852 290642 370110
rect 290752 369866 290780 371214
rect 291856 369866 291884 371282
rect 290752 369838 290996 369866
rect 291568 369844 291620 369850
rect 290108 369481 290136 369838
rect 291856 369838 292100 369866
rect 291568 369786 291620 369792
rect 291580 369730 291608 369786
rect 291364 369702 291608 369730
rect 290094 369472 290150 369481
rect 288992 369436 289044 369442
rect 291488 369442 291516 369702
rect 292224 369646 292252 375974
rect 292316 369866 292344 376110
rect 293052 376106 293080 376726
rect 293040 376100 293092 376106
rect 293040 376042 293092 376048
rect 293052 369986 293080 376042
rect 293328 374814 293356 400823
rect 293316 374808 293368 374814
rect 293316 374750 293368 374756
rect 294328 374808 294380 374814
rect 294328 374750 294380 374756
rect 293328 373674 293356 374750
rect 294340 374066 294368 374750
rect 294328 374060 294380 374066
rect 294328 374002 294380 374008
rect 293236 373646 293356 373674
rect 293236 370138 293264 373646
rect 293868 372156 293920 372162
rect 293868 372098 293920 372104
rect 293314 372056 293370 372065
rect 293314 371991 293370 372000
rect 293190 370110 293264 370138
rect 293040 369980 293092 369986
rect 293040 369922 293092 369928
rect 292580 369912 292632 369918
rect 292316 369860 292580 369866
rect 292316 369854 292632 369860
rect 292316 369838 292620 369854
rect 293052 369730 293080 369922
rect 293190 369852 293218 370110
rect 293328 369866 293356 371991
rect 293880 371890 293908 372098
rect 293868 371884 293920 371890
rect 293868 371826 293920 371832
rect 293880 370138 293908 371826
rect 294340 370138 294368 374002
rect 294512 373380 294564 373386
rect 294512 373322 294564 373328
rect 294524 373250 294552 373322
rect 294512 373244 294564 373250
rect 294512 373186 294564 373192
rect 293880 370110 293954 370138
rect 293328 369838 293572 369866
rect 293926 369852 293954 370110
rect 294294 370110 294368 370138
rect 294294 369852 294322 370110
rect 294524 369866 294552 373186
rect 294616 373182 294644 453494
rect 294696 452124 294748 452130
rect 294696 452066 294748 452072
rect 294708 373538 294736 452066
rect 297364 450900 297416 450906
rect 297364 450842 297416 450848
rect 294788 450696 294840 450702
rect 294788 450638 294840 450644
rect 294800 374814 294828 450638
rect 295984 450424 296036 450430
rect 295984 450366 296036 450372
rect 295338 398168 295394 398177
rect 295338 398103 295394 398112
rect 295352 396846 295380 398103
rect 295340 396840 295392 396846
rect 295340 396782 295392 396788
rect 295996 376754 296024 450366
rect 297376 383654 297404 450842
rect 298756 402966 298784 500958
rect 298836 455456 298888 455462
rect 298836 455398 298888 455404
rect 298744 402960 298796 402966
rect 298744 402902 298796 402908
rect 298742 399800 298798 399809
rect 298742 399735 298798 399744
rect 295812 376726 296024 376754
rect 297100 383626 297404 383654
rect 294788 374808 294840 374814
rect 294788 374750 294840 374756
rect 295812 374610 295840 376726
rect 295800 374604 295852 374610
rect 295800 374546 295852 374552
rect 294708 373510 294828 373538
rect 294604 373176 294656 373182
rect 294604 373118 294656 373124
rect 294800 372162 294828 373510
rect 295340 373176 295392 373182
rect 295340 373118 295392 373124
rect 294788 372156 294840 372162
rect 294788 372098 294840 372104
rect 294788 372020 294840 372026
rect 294788 371962 294840 371968
rect 294800 369866 294828 371962
rect 295352 370138 295380 373118
rect 295812 370138 295840 374546
rect 297100 374202 297128 383626
rect 298560 375964 298612 375970
rect 298560 375906 298612 375912
rect 298572 375630 298600 375906
rect 298560 375624 298612 375630
rect 298560 375566 298612 375572
rect 297456 375556 297508 375562
rect 297456 375498 297508 375504
rect 297088 374196 297140 374202
rect 297088 374138 297140 374144
rect 296628 373312 296680 373318
rect 296628 373254 296680 373260
rect 296640 372638 296668 373254
rect 296628 372632 296680 372638
rect 296628 372574 296680 372580
rect 295892 370388 295944 370394
rect 295892 370330 295944 370336
rect 295352 370110 295426 370138
rect 294524 369838 294676 369866
rect 294800 369838 295044 369866
rect 295398 369852 295426 370110
rect 295766 370110 295840 370138
rect 295766 369852 295794 370110
rect 295904 369866 295932 370330
rect 296640 369866 296668 372574
rect 297100 369866 297128 374138
rect 297364 373924 297416 373930
rect 297364 373866 297416 373872
rect 297376 371929 297404 373866
rect 297362 371920 297418 371929
rect 297362 371855 297418 371864
rect 295904 369838 296392 369866
rect 296516 369838 296668 369866
rect 296884 369838 297128 369866
rect 292836 369702 293080 369730
rect 291936 369640 291988 369646
rect 291936 369582 291988 369588
rect 292212 369640 292264 369646
rect 292212 369582 292264 369588
rect 291948 369458 291976 369582
rect 296364 369510 296392 369838
rect 297468 369594 297496 375498
rect 297824 373108 297876 373114
rect 297824 373050 297876 373056
rect 297836 369594 297864 373050
rect 298100 370660 298152 370666
rect 298100 370602 298152 370608
rect 298112 370054 298140 370602
rect 298100 370048 298152 370054
rect 298100 369990 298152 369996
rect 298112 369866 298140 369990
rect 298572 369866 298600 375566
rect 298756 372978 298784 399735
rect 298848 375494 298876 455398
rect 299492 453422 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 412652 703582 413508 703610
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 332520 700330 332548 703520
rect 348804 700398 348832 703520
rect 348792 700392 348844 700398
rect 348792 700334 348844 700340
rect 364340 700392 364392 700398
rect 364340 700334 364392 700340
rect 332508 700324 332560 700330
rect 332508 700266 332560 700272
rect 363604 698692 363656 698698
rect 363604 698634 363656 698640
rect 359464 670744 359516 670750
rect 359464 670686 359516 670692
rect 358452 576904 358504 576910
rect 358452 576846 358504 576852
rect 355324 484424 355376 484430
rect 355324 484366 355376 484372
rect 334716 457156 334768 457162
rect 334716 457098 334768 457104
rect 333520 457020 333572 457026
rect 333520 456962 333572 456968
rect 332048 456952 332100 456958
rect 332048 456894 332100 456900
rect 320824 456884 320876 456890
rect 320824 456826 320876 456832
rect 301504 455592 301556 455598
rect 301504 455534 301556 455540
rect 299480 453416 299532 453422
rect 299480 453358 299532 453364
rect 300122 451616 300178 451625
rect 300122 451551 300178 451560
rect 298926 401024 298982 401033
rect 298926 400959 298982 400968
rect 298940 375630 298968 400959
rect 298928 375624 298980 375630
rect 298928 375566 298980 375572
rect 298836 375488 298888 375494
rect 298836 375430 298888 375436
rect 298848 374898 298876 375430
rect 298848 374870 299244 374898
rect 298836 374128 298888 374134
rect 298836 374070 298888 374076
rect 298744 372972 298796 372978
rect 298744 372914 298796 372920
rect 298756 370138 298784 372914
rect 298848 372502 298876 374070
rect 298836 372496 298888 372502
rect 298836 372438 298888 372444
rect 297988 369838 298140 369866
rect 298356 369838 298600 369866
rect 298710 370110 298784 370138
rect 298710 369852 298738 370110
rect 298848 369866 298876 372438
rect 299216 369866 299244 374870
rect 299388 374672 299440 374678
rect 299388 374614 299440 374620
rect 299400 373114 299428 374614
rect 299388 373108 299440 373114
rect 299388 373050 299440 373056
rect 299940 373040 299992 373046
rect 299940 372982 299992 372988
rect 298848 369838 299092 369866
rect 299216 369838 299460 369866
rect 299952 369594 299980 372982
rect 300136 370161 300164 451551
rect 300214 449984 300270 449993
rect 300214 449919 300270 449928
rect 300228 375766 300256 449919
rect 300306 400072 300362 400081
rect 300306 400007 300362 400016
rect 300216 375760 300268 375766
rect 300216 375702 300268 375708
rect 300122 370152 300178 370161
rect 300122 370087 300178 370096
rect 300228 370002 300256 375702
rect 300320 373046 300348 400007
rect 300400 398676 300452 398682
rect 300400 398618 300452 398624
rect 300412 381857 300440 398618
rect 300398 381848 300454 381857
rect 300398 381783 300454 381792
rect 301516 375562 301544 455534
rect 304264 455524 304316 455530
rect 304264 455466 304316 455472
rect 302884 450764 302936 450770
rect 302884 450706 302936 450712
rect 301594 446448 301650 446457
rect 301594 446383 301650 446392
rect 301608 376922 301636 446383
rect 302148 392828 302200 392834
rect 302148 392770 302200 392776
rect 301596 376916 301648 376922
rect 301596 376858 301648 376864
rect 301504 375556 301556 375562
rect 301504 375498 301556 375504
rect 300860 373448 300912 373454
rect 300860 373390 300912 373396
rect 300308 373040 300360 373046
rect 300308 372982 300360 372988
rect 300872 372910 300900 373390
rect 300860 372904 300912 372910
rect 300860 372846 300912 372852
rect 300308 370932 300360 370938
rect 300308 370874 300360 370880
rect 300320 370326 300348 370874
rect 300308 370320 300360 370326
rect 300308 370262 300360 370268
rect 300182 369974 300256 370002
rect 300182 369852 300210 369974
rect 300320 369866 300348 370262
rect 300872 370138 300900 372846
rect 301044 372768 301096 372774
rect 301044 372710 301096 372716
rect 300872 370110 300946 370138
rect 300320 369838 300564 369866
rect 300918 369852 300946 370110
rect 301056 370054 301084 372710
rect 301504 370728 301556 370734
rect 301504 370670 301556 370676
rect 301044 370048 301096 370054
rect 301044 369990 301096 369996
rect 301516 369866 301544 370670
rect 301608 370138 301636 376858
rect 301608 370110 301682 370138
rect 301300 369838 301544 369866
rect 301654 369852 301682 370110
rect 301872 370048 301924 370054
rect 301872 369990 301924 369996
rect 301884 369866 301912 369990
rect 301884 369838 302036 369866
rect 297252 369566 297496 369594
rect 297620 369566 297864 369594
rect 299828 369566 299980 369594
rect 301424 369578 301452 369838
rect 301412 369572 301464 369578
rect 301412 369514 301464 369520
rect 290094 369407 290150 369416
rect 291476 369436 291528 369442
rect 288992 369378 289044 369384
rect 291732 369430 291976 369458
rect 296352 369504 296404 369510
rect 302160 369481 302188 392770
rect 302896 376754 302924 450706
rect 302974 398304 303030 398313
rect 302974 398239 303030 398248
rect 302988 385801 303016 398239
rect 303344 392760 303396 392766
rect 303344 392702 303396 392708
rect 302974 385792 303030 385801
rect 302974 385727 303030 385736
rect 302620 376726 302924 376754
rect 302620 375902 302648 376726
rect 302608 375896 302660 375902
rect 302608 375838 302660 375844
rect 302620 369730 302648 375838
rect 303252 374468 303304 374474
rect 303252 374410 303304 374416
rect 303264 372434 303292 374410
rect 303252 372428 303304 372434
rect 303252 372370 303304 372376
rect 302974 370832 303030 370841
rect 302974 370767 303030 370776
rect 302744 369880 302800 369889
rect 302988 369866 303016 370767
rect 303264 369866 303292 372370
rect 302800 369838 303016 369866
rect 303140 369838 303292 369866
rect 302744 369815 302800 369824
rect 302404 369702 302648 369730
rect 303356 369481 303384 392702
rect 304276 379846 304304 455466
rect 307024 454912 307076 454918
rect 307024 454854 307076 454860
rect 304356 449336 304408 449342
rect 304356 449278 304408 449284
rect 303620 379840 303672 379846
rect 303620 379782 303672 379788
rect 304264 379840 304316 379846
rect 304264 379782 304316 379788
rect 303632 379514 303660 379782
rect 303632 379486 304304 379514
rect 304172 373516 304224 373522
rect 304172 373458 304224 373464
rect 303528 372836 303580 372842
rect 303528 372778 303580 372784
rect 303540 372366 303568 372778
rect 303528 372360 303580 372366
rect 303528 372302 303580 372308
rect 303540 370138 303568 372302
rect 304080 371884 304132 371890
rect 304080 371826 304132 371832
rect 303494 370110 303568 370138
rect 303494 369852 303522 370110
rect 304092 369730 304120 371826
rect 304184 370138 304212 373458
rect 304276 370818 304304 379486
rect 304368 374406 304396 449278
rect 305644 449268 305696 449274
rect 305644 449210 305696 449216
rect 305000 409216 305052 409222
rect 305000 409158 305052 409164
rect 305012 405686 305040 409158
rect 305000 405680 305052 405686
rect 305000 405622 305052 405628
rect 305092 398472 305144 398478
rect 305092 398414 305144 398420
rect 305000 398404 305052 398410
rect 305000 398346 305052 398352
rect 305012 396001 305040 398346
rect 304998 395992 305054 396001
rect 304998 395927 305054 395936
rect 305104 395185 305132 398414
rect 305090 395176 305146 395185
rect 305090 395111 305146 395120
rect 305656 376754 305684 449210
rect 305736 405680 305788 405686
rect 305736 405622 305788 405628
rect 305748 383654 305776 405622
rect 307036 383654 307064 454854
rect 317604 454504 317656 454510
rect 317604 454446 317656 454452
rect 316868 454368 316920 454374
rect 316868 454310 316920 454316
rect 309048 453416 309100 453422
rect 309048 453358 309100 453364
rect 308402 452840 308458 452849
rect 308402 452775 308458 452784
rect 307760 450492 307812 450498
rect 307760 450434 307812 450440
rect 307668 397520 307720 397526
rect 307668 397462 307720 397468
rect 307680 394670 307708 397462
rect 307668 394664 307720 394670
rect 307668 394606 307720 394612
rect 305748 383626 305868 383654
rect 307036 383626 307156 383654
rect 305380 376726 305684 376754
rect 304356 374400 304408 374406
rect 304356 374342 304408 374348
rect 304368 373522 304396 374342
rect 305380 374338 305408 376726
rect 305368 374332 305420 374338
rect 305368 374274 305420 374280
rect 304356 373516 304408 373522
rect 304356 373458 304408 373464
rect 305092 370864 305144 370870
rect 304276 370790 304764 370818
rect 305092 370806 305144 370812
rect 304184 370110 304258 370138
rect 304230 369852 304258 370110
rect 304736 369866 304764 370790
rect 305104 370190 305132 370806
rect 305092 370184 305144 370190
rect 305380 370138 305408 374274
rect 305840 371754 305868 383626
rect 306196 374740 306248 374746
rect 306196 374682 306248 374688
rect 305828 371748 305880 371754
rect 305828 371690 305880 371696
rect 305460 370796 305512 370802
rect 305460 370738 305512 370744
rect 305092 370126 305144 370132
rect 304736 369838 304980 369866
rect 305104 369782 305132 370126
rect 305334 370110 305408 370138
rect 305334 369852 305362 370110
rect 305472 369866 305500 370738
rect 305840 369866 305868 371690
rect 305472 369838 305716 369866
rect 305840 369838 306084 369866
rect 303876 369702 304120 369730
rect 304724 369776 304776 369782
rect 304724 369718 304776 369724
rect 305092 369776 305144 369782
rect 305092 369718 305144 369724
rect 306208 369730 306236 374682
rect 307128 373930 307156 383626
rect 307772 379514 307800 450434
rect 308128 411936 308180 411942
rect 308128 411878 308180 411884
rect 308140 411262 308168 411878
rect 308128 411256 308180 411262
rect 308128 411198 308180 411204
rect 307944 391944 307996 391950
rect 307944 391886 307996 391892
rect 307956 390697 307984 391886
rect 307942 390688 307998 390697
rect 307942 390623 307998 390632
rect 308416 383654 308444 452775
rect 309060 449274 309088 453358
rect 315304 453144 315356 453150
rect 315304 453086 315356 453092
rect 313924 450152 313976 450158
rect 313924 450094 313976 450100
rect 314014 450120 314070 450129
rect 309048 449268 309100 449274
rect 309048 449210 309100 449216
rect 309140 449200 309192 449206
rect 309140 449142 309192 449148
rect 309048 411256 309100 411262
rect 309048 411198 309100 411204
rect 308324 383626 308444 383654
rect 307772 379486 307892 379514
rect 307864 376786 307892 379486
rect 307852 376780 307904 376786
rect 307852 376722 307904 376728
rect 307116 373924 307168 373930
rect 307116 373866 307168 373872
rect 306564 370252 306616 370258
rect 306564 370194 306616 370200
rect 306576 369866 306604 370194
rect 307128 370138 307156 373866
rect 307300 372564 307352 372570
rect 307300 372506 307352 372512
rect 307128 370110 307202 370138
rect 306576 369852 306820 369866
rect 307174 369852 307202 370110
rect 307312 369866 307340 372506
rect 307760 371680 307812 371686
rect 307760 371622 307812 371628
rect 307772 371210 307800 371622
rect 307760 371204 307812 371210
rect 307760 371146 307812 371152
rect 307864 370138 307892 376722
rect 308324 371754 308352 383626
rect 308404 374536 308456 374542
rect 308404 374478 308456 374484
rect 308312 371748 308364 371754
rect 308312 371690 308364 371696
rect 308324 370138 308352 371690
rect 307864 370110 307938 370138
rect 306576 369838 306834 369852
rect 307312 369838 307556 369866
rect 307910 369852 307938 370110
rect 308278 370110 308352 370138
rect 308278 369852 308306 370110
rect 308416 369866 308444 374478
rect 309060 370138 309088 411198
rect 309152 379778 309180 449142
rect 312542 448896 312598 448905
rect 312542 448831 312598 448840
rect 309782 447808 309838 447817
rect 309782 447743 309838 447752
rect 309140 379772 309192 379778
rect 309140 379714 309192 379720
rect 309014 370110 309088 370138
rect 308416 369838 308660 369866
rect 309014 369852 309042 370110
rect 309152 369866 309180 379714
rect 309796 375465 309824 447743
rect 311164 443692 311216 443698
rect 311164 443634 311216 443640
rect 311176 419490 311204 443634
rect 311900 420232 311952 420238
rect 311900 420174 311952 420180
rect 311912 419490 311940 420174
rect 311164 419484 311216 419490
rect 311164 419426 311216 419432
rect 311900 419484 311952 419490
rect 311900 419426 311952 419432
rect 311176 418198 311204 419426
rect 310704 418192 310756 418198
rect 310704 418134 310756 418140
rect 311164 418192 311216 418198
rect 311164 418134 311216 418140
rect 310520 414724 310572 414730
rect 310520 414666 310572 414672
rect 310532 413982 310560 414666
rect 310520 413976 310572 413982
rect 310520 413918 310572 413924
rect 310428 407788 310480 407794
rect 310428 407730 310480 407736
rect 310440 407046 310468 407730
rect 309876 407040 309928 407046
rect 309876 406982 309928 406988
rect 310428 407040 310480 407046
rect 310428 406982 310480 406988
rect 309888 383654 309916 406982
rect 309968 398540 310020 398546
rect 309968 398482 310020 398488
rect 309980 391921 310008 398482
rect 309966 391912 310022 391921
rect 309966 391847 310022 391856
rect 309888 383626 310284 383654
rect 309782 375456 309838 375465
rect 309782 375391 309838 375400
rect 309796 370138 309824 375391
rect 310256 371793 310284 383626
rect 310532 376754 310560 413918
rect 310532 376726 310652 376754
rect 310242 371784 310298 371793
rect 310242 371719 310298 371728
rect 309750 370110 309824 370138
rect 309152 369838 309396 369866
rect 309750 369852 309778 370110
rect 310256 369866 310284 371719
rect 310624 370297 310652 376726
rect 310716 371657 310744 418134
rect 311164 399560 311216 399566
rect 311164 399502 311216 399508
rect 311176 379514 311204 399502
rect 311808 391400 311860 391406
rect 311808 391342 311860 391348
rect 311716 391264 311768 391270
rect 311716 391206 311768 391212
rect 311728 379514 311756 391206
rect 311084 379486 311204 379514
rect 311452 379486 311756 379514
rect 311084 375698 311112 379486
rect 311072 375692 311124 375698
rect 311072 375634 311124 375640
rect 310702 371648 310758 371657
rect 310702 371583 310758 371592
rect 310610 370288 310666 370297
rect 310610 370223 310666 370232
rect 310256 369838 310500 369866
rect 306806 369730 306834 369838
rect 304736 369594 304764 369718
rect 306208 369702 306452 369730
rect 306806 369716 306972 369730
rect 306820 369702 306972 369716
rect 304612 369566 304764 369594
rect 296352 369446 296404 369452
rect 302146 369472 302202 369481
rect 302146 369407 302202 369416
rect 303342 369472 303398 369481
rect 306944 369442 306972 369702
rect 310624 369646 310652 370223
rect 310716 369889 310744 371583
rect 310702 369880 310758 369889
rect 311084 369866 311112 375634
rect 310868 369838 311112 369866
rect 310702 369815 310758 369824
rect 310612 369640 310664 369646
rect 310612 369582 310664 369588
rect 310980 369640 311032 369646
rect 311032 369588 311236 369594
rect 310980 369582 311236 369588
rect 310992 369566 311236 369582
rect 311452 369481 311480 379486
rect 311576 369880 311632 369889
rect 311576 369815 311632 369824
rect 311820 369617 311848 391342
rect 312556 376990 312584 448831
rect 312636 419484 312688 419490
rect 312636 419426 312688 419432
rect 311992 376984 312044 376990
rect 311992 376926 312044 376932
rect 312544 376984 312596 376990
rect 312544 376926 312596 376932
rect 312004 370138 312032 376926
rect 312648 371618 312676 419426
rect 313556 418124 313608 418130
rect 313556 418066 313608 418072
rect 313568 417722 313596 418066
rect 313556 417716 313608 417722
rect 313556 417658 313608 417664
rect 312728 416084 312780 416090
rect 312728 416026 312780 416032
rect 312740 387705 312768 416026
rect 313372 402280 313424 402286
rect 313372 402222 313424 402228
rect 312818 399528 312874 399537
rect 312818 399463 312874 399472
rect 312726 387696 312782 387705
rect 312726 387631 312782 387640
rect 312636 371612 312688 371618
rect 312636 371554 312688 371560
rect 312740 370138 312768 387631
rect 312832 379514 312860 399463
rect 313188 391468 313240 391474
rect 313188 391410 313240 391416
rect 312832 379486 312952 379514
rect 312924 375834 312952 379486
rect 312912 375828 312964 375834
rect 312912 375770 312964 375776
rect 312820 371612 312872 371618
rect 312820 371554 312872 371560
rect 311958 370110 312032 370138
rect 312556 370110 312768 370138
rect 311958 369852 311986 370110
rect 312082 369744 312138 369753
rect 312556 369730 312584 370110
rect 312832 369866 312860 371554
rect 312708 369838 312860 369866
rect 312924 369866 312952 375770
rect 312924 369838 313076 369866
rect 312138 369702 312584 369730
rect 312082 369679 312138 369688
rect 311806 369608 311862 369617
rect 311806 369543 311862 369552
rect 313200 369481 313228 391410
rect 313384 381002 313412 402222
rect 313372 380996 313424 381002
rect 313372 380938 313424 380944
rect 313384 373046 313412 380938
rect 313372 373040 313424 373046
rect 313372 372982 313424 372988
rect 313568 370433 313596 417658
rect 313936 402966 313964 450094
rect 314014 450055 314070 450064
rect 314028 417722 314056 450055
rect 314660 421592 314712 421598
rect 314660 421534 314712 421540
rect 314672 420918 314700 421534
rect 314660 420912 314712 420918
rect 314660 420854 314712 420860
rect 314016 417716 314068 417722
rect 314016 417658 314068 417664
rect 314016 405000 314068 405006
rect 314016 404942 314068 404948
rect 314028 404258 314056 404942
rect 315316 404326 315344 453086
rect 316776 452940 316828 452946
rect 316776 452882 316828 452888
rect 316684 452736 316736 452742
rect 316684 452678 316736 452684
rect 315580 422340 315632 422346
rect 315580 422282 315632 422288
rect 315396 420912 315448 420918
rect 315396 420854 315448 420860
rect 315304 404320 315356 404326
rect 315304 404262 315356 404268
rect 314016 404252 314068 404258
rect 314016 404194 314068 404200
rect 313924 402960 313976 402966
rect 313924 402902 313976 402908
rect 313936 402286 313964 402902
rect 313924 402280 313976 402286
rect 313924 402222 313976 402228
rect 313922 401296 313978 401305
rect 313922 401231 313978 401240
rect 313936 378486 313964 401231
rect 313924 378480 313976 378486
rect 313924 378422 313976 378428
rect 313936 378282 313964 378422
rect 313924 378276 313976 378282
rect 313924 378218 313976 378224
rect 314028 371550 314056 404194
rect 315316 402974 315344 404262
rect 314948 402946 315344 402974
rect 314292 392148 314344 392154
rect 314292 392090 314344 392096
rect 314200 378276 314252 378282
rect 314200 378218 314252 378224
rect 314016 371544 314068 371550
rect 314016 371486 314068 371492
rect 313554 370424 313610 370433
rect 313554 370359 313610 370368
rect 313568 369866 313596 370359
rect 314028 369866 314056 371486
rect 314212 370138 314240 378218
rect 313444 369838 313596 369866
rect 313812 369838 314056 369866
rect 314166 370110 314240 370138
rect 314166 369852 314194 370110
rect 314304 369481 314332 392090
rect 314384 391536 314436 391542
rect 314384 391478 314436 391484
rect 314396 369617 314424 391478
rect 314948 383654 314976 402946
rect 315302 399664 315358 399673
rect 315302 399599 315358 399608
rect 314948 383626 315252 383654
rect 314844 380384 314896 380390
rect 314844 380326 314896 380332
rect 314856 379914 314884 380326
rect 314844 379908 314896 379914
rect 314844 379850 314896 379856
rect 314856 379514 314884 379850
rect 315224 379514 315252 383626
rect 315316 380390 315344 399599
rect 315304 380384 315356 380390
rect 315304 380326 315356 380332
rect 314856 379486 315068 379514
rect 315224 379486 315344 379514
rect 314936 373652 314988 373658
rect 314936 373594 314988 373600
rect 314660 373040 314712 373046
rect 314660 372982 314712 372988
rect 314382 369608 314438 369617
rect 314672 369594 314700 372982
rect 314948 372570 314976 373594
rect 314936 372564 314988 372570
rect 314936 372506 314988 372512
rect 314948 370138 314976 372506
rect 314902 370110 314976 370138
rect 314902 369852 314930 370110
rect 315040 369866 315068 379486
rect 315316 370138 315344 379486
rect 315408 373538 315436 420854
rect 315488 403028 315540 403034
rect 315488 402970 315540 402976
rect 315500 373658 315528 402970
rect 315592 402898 315620 422282
rect 316224 407108 316276 407114
rect 316224 407050 316276 407056
rect 315580 402892 315632 402898
rect 315580 402834 315632 402840
rect 316132 402892 316184 402898
rect 316132 402834 316184 402840
rect 315856 391332 315908 391338
rect 315856 391274 315908 391280
rect 315488 373652 315540 373658
rect 315488 373594 315540 373600
rect 315408 373510 315804 373538
rect 315776 371414 315804 373510
rect 315764 371408 315816 371414
rect 315764 371350 315816 371356
rect 315316 370110 315436 370138
rect 315408 369866 315436 370110
rect 315040 369838 315284 369866
rect 315408 369838 315652 369866
rect 315776 369730 315804 371350
rect 315868 369889 315896 391274
rect 316144 376854 316172 402834
rect 316132 376848 316184 376854
rect 316132 376790 316184 376796
rect 315854 369880 315910 369889
rect 316144 369866 316172 376790
rect 316236 371618 316264 407050
rect 316696 394670 316724 452678
rect 316788 422346 316816 452882
rect 316776 422340 316828 422346
rect 316776 422282 316828 422288
rect 316880 407114 316908 454310
rect 316868 407108 316920 407114
rect 316868 407050 316920 407056
rect 316316 394664 316368 394670
rect 316316 394606 316368 394612
rect 316684 394664 316736 394670
rect 316684 394606 316736 394612
rect 316328 383654 316356 394606
rect 316328 383626 316540 383654
rect 316224 371612 316276 371618
rect 316224 371554 316276 371560
rect 316512 369866 316540 383626
rect 316868 371612 316920 371618
rect 316868 371554 316920 371560
rect 316880 369866 316908 371554
rect 317616 370122 317644 454446
rect 319444 454300 319496 454306
rect 319444 454242 319496 454248
rect 318064 452872 318116 452878
rect 318064 452814 318116 452820
rect 317972 374264 318024 374270
rect 317972 374206 318024 374212
rect 317604 370116 317656 370122
rect 317604 370058 317656 370064
rect 317616 369866 317644 370058
rect 316144 369838 316388 369866
rect 316512 369838 316756 369866
rect 316880 369838 317124 369866
rect 317616 369838 317860 369866
rect 315854 369815 315910 369824
rect 317604 369776 317656 369782
rect 315776 369702 316020 369730
rect 317492 369724 317604 369730
rect 317492 369718 317656 369724
rect 317492 369702 317644 369718
rect 314548 369566 314700 369594
rect 317984 369594 318012 374206
rect 318076 371686 318104 452814
rect 318156 450288 318208 450294
rect 318156 450230 318208 450236
rect 318168 383654 318196 450230
rect 318708 389972 318760 389978
rect 318708 389914 318760 389920
rect 318168 383626 318380 383654
rect 318064 371680 318116 371686
rect 318064 371622 318116 371628
rect 318076 369782 318104 371622
rect 318352 370530 318380 383626
rect 318432 374808 318484 374814
rect 318432 374750 318484 374756
rect 318444 374270 318472 374750
rect 318432 374264 318484 374270
rect 318432 374206 318484 374212
rect 318340 370524 318392 370530
rect 318340 370466 318392 370472
rect 318352 369866 318380 370466
rect 318352 369838 318596 369866
rect 318064 369776 318116 369782
rect 318064 369718 318116 369724
rect 317984 369566 318228 369594
rect 314382 369543 314438 369552
rect 318720 369481 318748 389914
rect 319076 385008 319128 385014
rect 319076 384950 319128 384956
rect 319088 383722 319116 384950
rect 319076 383716 319128 383722
rect 319076 383658 319128 383664
rect 318892 382424 318944 382430
rect 318892 382366 318944 382372
rect 318904 382294 318932 382366
rect 318892 382288 318944 382294
rect 318892 382230 318944 382236
rect 318984 382288 319036 382294
rect 318984 382230 319036 382236
rect 318904 374746 318932 382230
rect 318892 374740 318944 374746
rect 318892 374682 318944 374688
rect 318996 370122 319024 382230
rect 318984 370116 319036 370122
rect 318984 370058 319036 370064
rect 319088 369866 319116 383658
rect 319456 382294 319484 454242
rect 319536 450220 319588 450226
rect 319536 450162 319588 450168
rect 319444 382288 319496 382294
rect 319444 382230 319496 382236
rect 319548 378418 319576 450162
rect 319628 436756 319680 436762
rect 319628 436698 319680 436704
rect 319640 382430 319668 436698
rect 319718 401160 319774 401169
rect 319718 401095 319774 401104
rect 319732 385014 319760 401095
rect 319812 390108 319864 390114
rect 319812 390050 319864 390056
rect 319720 385008 319772 385014
rect 319720 384950 319772 384956
rect 319628 382424 319680 382430
rect 319628 382366 319680 382372
rect 319536 378412 319588 378418
rect 319536 378354 319588 378360
rect 319168 374740 319220 374746
rect 319168 374682 319220 374688
rect 318964 369838 319116 369866
rect 319180 369866 319208 374682
rect 319548 369866 319576 378354
rect 319180 369838 319332 369866
rect 319548 369838 319700 369866
rect 319824 369481 319852 390050
rect 319904 390040 319956 390046
rect 319904 389982 319956 389988
rect 319916 369617 319944 389982
rect 320180 386368 320232 386374
rect 320180 386310 320232 386316
rect 320192 385218 320220 386310
rect 320180 385212 320232 385218
rect 320180 385154 320232 385160
rect 320192 374746 320220 385154
rect 320836 381342 320864 456826
rect 327816 455796 327868 455802
rect 327816 455738 327868 455744
rect 324964 455728 325016 455734
rect 324964 455670 325016 455676
rect 322204 455660 322256 455666
rect 322204 455602 322256 455608
rect 320916 450628 320968 450634
rect 320916 450570 320968 450576
rect 320272 381336 320324 381342
rect 320272 381278 320324 381284
rect 320824 381336 320876 381342
rect 320824 381278 320876 381284
rect 320284 381070 320312 381278
rect 320272 381064 320324 381070
rect 320272 381006 320324 381012
rect 320180 374740 320232 374746
rect 320180 374682 320232 374688
rect 320284 370122 320312 381006
rect 320928 379574 320956 450570
rect 321008 450356 321060 450362
rect 321008 450298 321060 450304
rect 321020 386374 321048 450298
rect 321376 394188 321428 394194
rect 321376 394130 321428 394136
rect 321284 393440 321336 393446
rect 321284 393382 321336 393388
rect 321008 386368 321060 386374
rect 321008 386310 321060 386316
rect 320916 379568 320968 379574
rect 320916 379510 320968 379516
rect 320640 371408 320692 371414
rect 320640 371350 320692 371356
rect 320042 370116 320094 370122
rect 320042 370058 320094 370064
rect 320272 370116 320324 370122
rect 320272 370058 320324 370064
rect 320054 369852 320082 370058
rect 320652 369730 320680 371350
rect 320928 369866 320956 379510
rect 321008 374740 321060 374746
rect 321008 374682 321060 374688
rect 320804 369838 320956 369866
rect 321020 369866 321048 374682
rect 321020 369838 321172 369866
rect 320436 369702 320680 369730
rect 319902 369608 319958 369617
rect 319902 369543 319958 369552
rect 321296 369481 321324 393382
rect 321388 369617 321416 394130
rect 321744 385008 321796 385014
rect 321744 384950 321796 384956
rect 321756 383790 321784 384950
rect 321744 383784 321796 383790
rect 321744 383726 321796 383732
rect 321756 383654 321784 383726
rect 321756 383626 322060 383654
rect 321652 382696 321704 382702
rect 321652 382638 321704 382644
rect 321664 382498 321692 382638
rect 321652 382492 321704 382498
rect 321652 382434 321704 382440
rect 321664 374610 321692 382434
rect 321836 375420 321888 375426
rect 321836 375362 321888 375368
rect 321652 374604 321704 374610
rect 321652 374546 321704 374552
rect 321848 370138 321876 375362
rect 321514 370116 321566 370122
rect 321848 370110 321922 370138
rect 321514 370058 321566 370064
rect 321526 369852 321554 370058
rect 321894 369852 321922 370110
rect 322032 369866 322060 383626
rect 322216 371890 322244 455602
rect 322388 454436 322440 454442
rect 322388 454378 322440 454384
rect 322296 453008 322348 453014
rect 322296 452950 322348 452956
rect 322308 375426 322336 452950
rect 322400 385014 322428 454378
rect 323676 453076 323728 453082
rect 323676 453018 323728 453024
rect 323584 452804 323636 452810
rect 323584 452746 323636 452752
rect 322480 445052 322532 445058
rect 322480 444994 322532 445000
rect 322388 385008 322440 385014
rect 322388 384950 322440 384956
rect 322492 382702 322520 444994
rect 322940 386368 322992 386374
rect 322940 386310 322992 386316
rect 322952 385150 322980 386310
rect 322940 385144 322992 385150
rect 322940 385086 322992 385092
rect 322480 382696 322532 382702
rect 322480 382638 322532 382644
rect 322296 375420 322348 375426
rect 322296 375362 322348 375368
rect 322388 374604 322440 374610
rect 322388 374546 322440 374552
rect 322204 371884 322256 371890
rect 322204 371826 322256 371832
rect 322400 369866 322428 374546
rect 322848 373040 322900 373046
rect 322848 372982 322900 372988
rect 322860 369866 322888 372982
rect 322952 371396 322980 385086
rect 323032 381744 323084 381750
rect 323032 381686 323084 381692
rect 323044 380934 323072 381686
rect 323032 380928 323084 380934
rect 323032 380870 323084 380876
rect 323044 373046 323072 380870
rect 323596 379514 323624 452746
rect 323688 381750 323716 453018
rect 323766 399936 323822 399945
rect 323766 399871 323822 399880
rect 323780 386374 323808 399871
rect 324228 397996 324280 398002
rect 324228 397938 324280 397944
rect 324240 390017 324268 397938
rect 324226 390008 324282 390017
rect 324226 389943 324282 389952
rect 324596 388816 324648 388822
rect 324596 388758 324648 388764
rect 323768 386368 323820 386374
rect 323768 386310 323820 386316
rect 324318 385792 324374 385801
rect 324318 385727 324374 385736
rect 324332 383858 324360 385727
rect 324608 385082 324636 388758
rect 324596 385076 324648 385082
rect 324596 385018 324648 385024
rect 324320 383852 324372 383858
rect 324320 383794 324372 383800
rect 324332 383654 324360 383794
rect 324332 383626 324452 383654
rect 323676 381744 323728 381750
rect 323676 381686 323728 381692
rect 324320 379568 324372 379574
rect 323596 379486 323900 379514
rect 324320 379510 324372 379516
rect 323872 378214 323900 379486
rect 323860 378208 323912 378214
rect 323860 378150 323912 378156
rect 323032 373040 323084 373046
rect 323032 372982 323084 372988
rect 322952 371368 323164 371396
rect 323136 369866 323164 371368
rect 323584 371340 323636 371346
rect 323584 371282 323636 371288
rect 322032 369838 322276 369866
rect 322400 369838 322644 369866
rect 322860 369838 323012 369866
rect 323136 369838 323380 369866
rect 321374 369608 321430 369617
rect 323596 369594 323624 371282
rect 323872 369866 323900 378150
rect 324332 374814 324360 379510
rect 324320 374808 324372 374814
rect 324320 374750 324372 374756
rect 324424 374542 324452 383626
rect 324504 379636 324556 379642
rect 324504 379578 324556 379584
rect 324516 374610 324544 379578
rect 324504 374604 324556 374610
rect 324504 374546 324556 374552
rect 324412 374536 324464 374542
rect 324412 374478 324464 374484
rect 324608 369866 324636 385018
rect 324976 379514 325004 455670
rect 325056 453212 325108 453218
rect 325056 453154 325108 453160
rect 325068 379574 325096 453154
rect 325148 407788 325200 407794
rect 325148 407730 325200 407736
rect 325160 379642 325188 407730
rect 327540 399900 327592 399906
rect 327540 399842 327592 399848
rect 327552 398274 327580 399842
rect 327724 398812 327776 398818
rect 327724 398754 327776 398760
rect 327540 398268 327592 398274
rect 327540 398210 327592 398216
rect 325148 379636 325200 379642
rect 325148 379578 325200 379584
rect 324884 379486 325004 379514
rect 325056 379568 325108 379574
rect 325056 379510 325108 379516
rect 324688 374604 324740 374610
rect 324688 374546 324740 374552
rect 323872 369838 324116 369866
rect 324484 369838 324636 369866
rect 324700 369866 324728 374546
rect 324884 370841 324912 379486
rect 324964 374808 325016 374814
rect 324964 374750 325016 374756
rect 324870 370832 324926 370841
rect 324870 370767 324926 370776
rect 324976 369866 325004 374750
rect 325332 374536 325384 374542
rect 325332 374478 325384 374484
rect 325344 369866 325372 374478
rect 326252 371272 326304 371278
rect 326252 371214 326304 371220
rect 326264 369866 326292 371214
rect 324700 369838 324852 369866
rect 324976 369838 325220 369866
rect 325344 369838 325588 369866
rect 325956 369838 326292 369866
rect 323596 369566 323748 369594
rect 321374 369543 321430 369552
rect 311438 369472 311494 369481
rect 303342 369407 303398 369416
rect 306932 369436 306984 369442
rect 291476 369378 291528 369384
rect 311438 369407 311494 369416
rect 313186 369472 313242 369481
rect 313186 369407 313242 369416
rect 314290 369472 314346 369481
rect 314290 369407 314346 369416
rect 318706 369472 318762 369481
rect 318706 369407 318762 369416
rect 319810 369472 319866 369481
rect 319810 369407 319866 369416
rect 321282 369472 321338 369481
rect 321282 369407 321338 369416
rect 306932 369378 306984 369384
rect 285816 369336 285872 369345
rect 285816 369271 285872 369280
rect 287288 369336 287344 369345
rect 287288 369271 287344 369280
rect 309000 369336 309056 369345
rect 309000 369271 309056 369280
rect 310104 369336 310160 369345
rect 310104 369271 310160 369280
rect 282274 360904 282330 360913
rect 282274 360839 282330 360848
rect 282182 353968 282238 353977
rect 282182 353903 282238 353912
rect 327446 333296 327502 333305
rect 327446 333231 327502 333240
rect 327460 321609 327488 333231
rect 327538 330440 327594 330449
rect 327538 330375 327594 330384
rect 327446 321600 327502 321609
rect 327446 321535 327502 321544
rect 282274 321328 282330 321337
rect 282274 321263 282330 321272
rect 282288 320793 282316 321263
rect 282274 320784 282330 320793
rect 282274 320719 282330 320728
rect 283240 320784 283296 320793
rect 283240 320719 283296 320728
rect 284252 320784 284308 320793
rect 284252 320719 284308 320728
rect 287472 320784 287528 320793
rect 287472 320719 287528 320728
rect 288208 320784 288264 320793
rect 288208 320719 288264 320728
rect 290600 320784 290656 320793
rect 290600 320719 290656 320728
rect 291152 320784 291208 320793
rect 291152 320719 291208 320728
rect 291888 320784 291944 320793
rect 291888 320719 291944 320728
rect 292624 320784 292680 320793
rect 292624 320719 292680 320728
rect 296488 320784 296544 320793
rect 296488 320719 296544 320728
rect 297316 320784 297372 320793
rect 297316 320719 297372 320728
rect 298144 320784 298200 320793
rect 298144 320719 298200 320728
rect 299064 320784 299120 320793
rect 303388 320784 303444 320793
rect 299906 320754 299934 320756
rect 299064 320719 299120 320728
rect 299894 320748 299946 320754
rect 303388 320719 303444 320728
rect 306700 320784 306756 320793
rect 306700 320719 306756 320728
rect 308816 320784 308872 320793
rect 308816 320719 308872 320728
rect 323536 320784 323592 320793
rect 323536 320719 323592 320728
rect 324088 320784 324144 320793
rect 324088 320719 324144 320728
rect 324364 320784 324420 320793
rect 324364 320719 324420 320728
rect 325192 320784 325248 320793
rect 325192 320719 325248 320728
rect 325744 320784 325800 320793
rect 325744 320719 325800 320728
rect 327032 320784 327088 320793
rect 327032 320719 327088 320728
rect 299894 320690 299946 320696
rect 283332 320648 283388 320657
rect 282276 320612 282328 320618
rect 283332 320583 283388 320592
rect 283608 320648 283664 320657
rect 283608 320583 283664 320592
rect 286184 320648 286240 320657
rect 286184 320583 286240 320592
rect 313048 320648 313104 320657
rect 313048 320583 313104 320592
rect 315808 320648 315864 320657
rect 315808 320583 315864 320592
rect 317096 320648 317152 320657
rect 317096 320583 317152 320592
rect 317648 320648 317704 320657
rect 317648 320583 317704 320592
rect 318016 320648 318072 320657
rect 318016 320583 318072 320592
rect 318200 320648 318256 320657
rect 318200 320583 318256 320592
rect 318936 320648 318992 320657
rect 318936 320583 318992 320592
rect 319212 320648 319268 320657
rect 319212 320583 319268 320592
rect 282276 320554 282328 320560
rect 282288 320521 282316 320554
rect 282274 320512 282330 320521
rect 282184 320476 282236 320482
rect 282274 320447 282330 320456
rect 282872 320512 282928 320521
rect 282872 320447 282928 320456
rect 283976 320512 284032 320521
rect 283976 320447 284032 320456
rect 286552 320512 286608 320521
rect 286552 320447 286608 320456
rect 288668 320512 288724 320521
rect 288668 320447 288724 320456
rect 292348 320512 292404 320521
rect 292348 320447 292404 320456
rect 293728 320512 293784 320521
rect 293728 320447 293784 320456
rect 294004 320512 294060 320521
rect 294004 320447 294060 320456
rect 294832 320512 294888 320521
rect 294832 320447 294888 320456
rect 297868 320512 297924 320521
rect 297868 320447 297924 320456
rect 298604 320512 298660 320521
rect 298604 320447 298660 320456
rect 305596 320512 305652 320521
rect 305596 320447 305652 320456
rect 308356 320512 308412 320521
rect 308356 320447 308412 320456
rect 310380 320512 310436 320521
rect 310380 320447 310436 320456
rect 322064 320512 322120 320521
rect 322064 320447 322120 320456
rect 322248 320512 322304 320521
rect 322248 320447 322304 320456
rect 323352 320512 323408 320521
rect 323352 320447 323408 320456
rect 323812 320512 323868 320521
rect 323812 320447 323868 320456
rect 324640 320512 324696 320521
rect 324640 320447 324696 320456
rect 326112 320512 326168 320521
rect 326112 320447 326168 320456
rect 282184 320418 282236 320424
rect 282196 320210 282224 320418
rect 282184 320204 282236 320210
rect 282184 320146 282236 320152
rect 282184 320000 282236 320006
rect 282184 319942 282236 319948
rect 282196 318850 282224 319942
rect 282184 318844 282236 318850
rect 282184 318786 282236 318792
rect 282092 318776 282144 318782
rect 282092 318718 282144 318724
rect 281632 318164 281684 318170
rect 281632 318106 281684 318112
rect 282288 318102 282316 320447
rect 284344 320376 284400 320385
rect 284344 320311 284400 320320
rect 285448 320376 285504 320385
rect 285448 320311 285504 320320
rect 285724 320376 285780 320385
rect 285724 320311 285780 320320
rect 287748 320376 287804 320385
rect 287748 320311 287804 320320
rect 289496 320376 289552 320385
rect 289496 320311 289552 320320
rect 290048 320376 290104 320385
rect 290048 320311 290104 320320
rect 291704 320376 291760 320385
rect 291704 320311 291760 320320
rect 307896 320376 307952 320385
rect 307896 320311 307952 320320
rect 309552 320376 309608 320385
rect 309552 320311 309608 320320
rect 310104 320376 310160 320385
rect 310104 320311 310160 320320
rect 310288 320376 310344 320385
rect 310288 320311 310344 320320
rect 310656 320376 310712 320385
rect 310656 320311 310712 320320
rect 311392 320376 311448 320385
rect 311392 320311 311448 320320
rect 316452 320376 316508 320385
rect 316452 320311 316508 320320
rect 320132 320376 320188 320385
rect 320132 320311 320188 320320
rect 320316 320376 320372 320385
rect 320316 320311 320372 320320
rect 320776 320376 320832 320385
rect 320776 320311 320832 320320
rect 321604 320376 321660 320385
rect 321604 320311 321660 320320
rect 323260 320376 323316 320385
rect 323260 320311 323316 320320
rect 324272 320376 324328 320385
rect 324272 320311 324328 320320
rect 325468 320376 325524 320385
rect 325468 320311 325524 320320
rect 326388 320376 326444 320385
rect 326388 320311 326444 320320
rect 327400 320376 327456 320385
rect 327400 320311 327456 320320
rect 282504 320240 282560 320249
rect 282504 320175 282560 320184
rect 292808 320240 292864 320249
rect 292808 320175 292864 320184
rect 293176 320240 293232 320249
rect 293176 320175 293232 320184
rect 294188 320240 294244 320249
rect 294188 320175 294244 320184
rect 294556 320240 294612 320249
rect 294556 320175 294612 320184
rect 295936 320240 295992 320249
rect 295936 320175 295992 320184
rect 297040 320240 297096 320249
rect 297040 320175 297096 320184
rect 297408 320240 297464 320249
rect 297408 320175 297464 320184
rect 298420 320240 298476 320249
rect 298420 320175 298476 320184
rect 302008 320240 302064 320249
rect 302008 320175 302064 320184
rect 307988 320240 308044 320249
rect 307988 320175 308044 320184
rect 312036 320240 312092 320249
rect 312036 320175 312092 320184
rect 312680 320240 312736 320249
rect 312680 320175 312736 320184
rect 313600 320240 313656 320249
rect 313600 320175 313656 320184
rect 314152 320240 314208 320249
rect 314152 320175 314208 320184
rect 316636 320240 316692 320249
rect 316636 320175 316692 320184
rect 317740 320240 317796 320249
rect 317740 320175 317796 320184
rect 283148 320104 283204 320113
rect 282610 319954 282638 320076
rect 282564 319926 282638 319954
rect 282368 319796 282420 319802
rect 282368 319738 282420 319744
rect 282380 319410 282408 319738
rect 282564 319569 282592 319926
rect 282702 319818 282730 320076
rect 282794 319954 282822 320076
rect 282794 319926 282868 319954
rect 282656 319790 282730 319818
rect 282550 319560 282606 319569
rect 282550 319495 282606 319504
rect 282656 319410 282684 319790
rect 282840 319716 282868 319926
rect 282380 319382 282684 319410
rect 282748 319688 282868 319716
rect 282978 319716 283006 320076
rect 283070 319784 283098 320076
rect 283792 320104 283848 320113
rect 283148 320039 283204 320048
rect 283162 319852 283190 320039
rect 283438 319852 283466 320076
rect 283530 319954 283558 320076
rect 283530 319926 283650 319954
rect 283622 319852 283650 319926
rect 283162 319824 283236 319852
rect 283438 319824 283512 319852
rect 283070 319756 283144 319784
rect 282978 319688 283052 319716
rect 282276 318096 282328 318102
rect 282276 318038 282328 318044
rect 282380 317880 282408 319382
rect 282460 318776 282512 318782
rect 282460 318718 282512 318724
rect 282104 317852 282408 317880
rect 280988 317416 281040 317422
rect 280988 317358 281040 317364
rect 280804 317348 280856 317354
rect 280804 317290 280856 317296
rect 280816 234054 280844 317290
rect 280896 315104 280948 315110
rect 280896 315046 280948 315052
rect 280908 235414 280936 315046
rect 282104 311894 282132 317852
rect 282276 316260 282328 316266
rect 282276 316202 282328 316208
rect 282184 314152 282236 314158
rect 282184 314094 282236 314100
rect 281644 311866 282132 311894
rect 281644 311302 281672 311866
rect 281632 311296 281684 311302
rect 281632 311238 281684 311244
rect 280988 307692 281040 307698
rect 280988 307634 281040 307640
rect 280896 235408 280948 235414
rect 280896 235350 280948 235356
rect 280804 234048 280856 234054
rect 280804 233990 280856 233996
rect 281000 230042 281028 307634
rect 282090 306912 282146 306921
rect 282090 306847 282146 306856
rect 281080 304904 281132 304910
rect 281080 304846 281132 304852
rect 281092 231713 281120 304846
rect 282104 235113 282132 306847
rect 282090 235104 282146 235113
rect 282090 235039 282146 235048
rect 281540 232756 281592 232762
rect 281540 232698 281592 232704
rect 281078 231704 281134 231713
rect 281078 231639 281134 231648
rect 281552 231062 281580 232698
rect 281540 231056 281592 231062
rect 281540 230998 281592 231004
rect 280988 230036 281040 230042
rect 280988 229978 281040 229984
rect 280802 218648 280858 218657
rect 280802 218583 280858 218592
rect 280436 153196 280488 153202
rect 280436 153138 280488 153144
rect 280252 144764 280304 144770
rect 280252 144706 280304 144712
rect 280816 126954 280844 218583
rect 281552 148442 281580 230998
rect 282196 219026 282224 314094
rect 282288 229974 282316 316202
rect 282368 310276 282420 310282
rect 282368 310218 282420 310224
rect 282276 229968 282328 229974
rect 282276 229910 282328 229916
rect 282380 224398 282408 310218
rect 282472 239057 282500 318718
rect 282748 318238 282776 319688
rect 282920 319388 282972 319394
rect 282920 319330 282972 319336
rect 282826 318744 282882 318753
rect 282826 318679 282882 318688
rect 282736 318232 282788 318238
rect 282736 318174 282788 318180
rect 282840 315330 282868 318679
rect 282932 317898 282960 319330
rect 283024 319161 283052 319688
rect 283116 319394 283144 319756
rect 283104 319388 283156 319394
rect 283104 319330 283156 319336
rect 283010 319152 283066 319161
rect 283010 319087 283066 319096
rect 283104 319116 283156 319122
rect 283104 319058 283156 319064
rect 283116 318889 283144 319058
rect 283102 318880 283158 318889
rect 283102 318815 283158 318824
rect 282920 317892 282972 317898
rect 282920 317834 282972 317840
rect 283116 317762 283144 318815
rect 282920 317756 282972 317762
rect 282920 317698 282972 317704
rect 283104 317756 283156 317762
rect 283104 317698 283156 317704
rect 282656 315302 282868 315330
rect 282656 310010 282684 315302
rect 282736 311976 282788 311982
rect 282736 311918 282788 311924
rect 282644 310004 282696 310010
rect 282644 309946 282696 309952
rect 282644 304496 282696 304502
rect 282644 304438 282696 304444
rect 282458 239048 282514 239057
rect 282458 238983 282514 238992
rect 282552 235272 282604 235278
rect 282552 235214 282604 235220
rect 282458 234016 282514 234025
rect 282458 233951 282514 233960
rect 282368 224392 282420 224398
rect 282368 224334 282420 224340
rect 282184 219020 282236 219026
rect 282184 218962 282236 218968
rect 282276 155848 282328 155854
rect 282276 155790 282328 155796
rect 282288 155242 282316 155790
rect 282276 155236 282328 155242
rect 282276 155178 282328 155184
rect 282472 155122 282500 233951
rect 282564 155854 282592 235214
rect 282656 227458 282684 304438
rect 282748 235482 282776 311918
rect 282828 310208 282880 310214
rect 282828 310150 282880 310156
rect 282736 235476 282788 235482
rect 282736 235418 282788 235424
rect 282840 234394 282868 310150
rect 282932 238921 282960 317698
rect 283208 317642 283236 319824
rect 283286 319424 283342 319433
rect 283286 319359 283342 319368
rect 283380 319388 283432 319394
rect 283300 317665 283328 319359
rect 283380 319330 283432 319336
rect 283024 317614 283236 317642
rect 283286 317656 283342 317665
rect 283024 294710 283052 317614
rect 283286 317591 283342 317600
rect 283392 316010 283420 319330
rect 283116 315982 283420 316010
rect 283116 300490 283144 315982
rect 283484 311894 283512 319824
rect 283576 319824 283650 319852
rect 283576 319394 283604 319824
rect 283714 319716 283742 320076
rect 284712 320104 284768 320113
rect 283792 320039 283848 320048
rect 283898 319818 283926 320076
rect 284082 319954 284110 320076
rect 284036 319926 284110 319954
rect 284174 319954 284202 320076
rect 284174 319926 284248 319954
rect 283898 319790 283972 319818
rect 283668 319688 283742 319716
rect 283564 319388 283616 319394
rect 283564 319330 283616 319336
rect 283668 317529 283696 319688
rect 283746 319424 283802 319433
rect 283746 319359 283802 319368
rect 283654 317520 283710 317529
rect 283654 317455 283710 317464
rect 283760 311894 283788 319359
rect 283944 318794 283972 319790
rect 283852 318766 283972 318794
rect 283852 317150 283880 318766
rect 284036 317801 284064 319926
rect 284220 318646 284248 319926
rect 284298 319832 284354 319841
rect 284450 319784 284478 320076
rect 284298 319767 284354 319776
rect 284208 318640 284260 318646
rect 284208 318582 284260 318588
rect 284022 317792 284078 317801
rect 284022 317727 284078 317736
rect 284116 317688 284168 317694
rect 284116 317630 284168 317636
rect 283840 317144 283892 317150
rect 283840 317086 283892 317092
rect 283208 311866 283512 311894
rect 283576 311866 283788 311894
rect 284128 311894 284156 317630
rect 284312 317506 284340 319767
rect 284404 319756 284478 319784
rect 284542 319784 284570 320076
rect 284634 319920 284662 320076
rect 285172 320104 285228 320113
rect 284712 320039 284768 320048
rect 284818 319954 284846 320076
rect 284772 319926 284846 319954
rect 284634 319892 284708 319920
rect 284542 319756 284616 319784
rect 284404 319716 284432 319756
rect 284404 319688 284524 319716
rect 284496 319258 284524 319688
rect 284484 319252 284536 319258
rect 284484 319194 284536 319200
rect 284390 317792 284446 317801
rect 284390 317727 284446 317736
rect 284220 317478 284340 317506
rect 284220 317257 284248 317478
rect 284206 317248 284262 317257
rect 284206 317183 284262 317192
rect 284300 317144 284352 317150
rect 284300 317086 284352 317092
rect 284128 311866 284248 311894
rect 283208 307630 283236 311866
rect 283196 307624 283248 307630
rect 283196 307566 283248 307572
rect 283104 300484 283156 300490
rect 283104 300426 283156 300432
rect 283116 296714 283144 300426
rect 283116 296686 283512 296714
rect 283484 296177 283512 296686
rect 283470 296168 283526 296177
rect 283470 296103 283526 296112
rect 283012 294704 283064 294710
rect 283012 294646 283064 294652
rect 283472 244928 283524 244934
rect 283472 244870 283524 244876
rect 283012 240984 283064 240990
rect 283012 240926 283064 240932
rect 283024 240378 283052 240926
rect 283012 240372 283064 240378
rect 283012 240314 283064 240320
rect 282918 238912 282974 238921
rect 282918 238847 282974 238856
rect 282918 236056 282974 236065
rect 282918 235991 282974 236000
rect 282828 234388 282880 234394
rect 282828 234330 282880 234336
rect 282644 227452 282696 227458
rect 282644 227394 282696 227400
rect 282552 155848 282604 155854
rect 282552 155790 282604 155796
rect 282288 155094 282500 155122
rect 282288 154494 282316 155094
rect 282276 154488 282328 154494
rect 282276 154430 282328 154436
rect 282288 153882 282316 154430
rect 282276 153876 282328 153882
rect 282276 153818 282328 153824
rect 281540 148436 281592 148442
rect 281540 148378 281592 148384
rect 281552 148170 281580 148378
rect 281540 148164 281592 148170
rect 281540 148106 281592 148112
rect 282184 145852 282236 145858
rect 282184 145794 282236 145800
rect 281448 144764 281500 144770
rect 281448 144706 281500 144712
rect 281460 144362 281488 144706
rect 281448 144356 281500 144362
rect 281448 144298 281500 144304
rect 280804 126948 280856 126954
rect 280804 126890 280856 126896
rect 281448 126948 281500 126954
rect 281448 126890 281500 126896
rect 281460 126410 281488 126890
rect 281448 126404 281500 126410
rect 281448 126346 281500 126352
rect 279424 113144 279476 113150
rect 279424 113086 279476 113092
rect 280158 108352 280214 108361
rect 280158 108287 280214 108296
rect 280172 16574 280200 108287
rect 278792 16546 279096 16574
rect 280172 16546 280752 16574
rect 278320 3392 278372 3398
rect 278320 3334 278372 3340
rect 278044 3052 278096 3058
rect 278044 2994 278096 3000
rect 278332 480 278360 3334
rect 277094 354 277206 480
rect 276676 326 277206 354
rect 277094 -960 277206 326
rect 278290 -960 278402 480
rect 279068 354 279096 16546
rect 280724 480 280752 16546
rect 282196 3058 282224 145794
rect 282932 16574 282960 235991
rect 283024 142118 283052 240314
rect 283484 236881 283512 244870
rect 283470 236872 283526 236881
rect 283470 236807 283526 236816
rect 283484 236065 283512 236807
rect 283470 236056 283526 236065
rect 283470 235991 283526 236000
rect 283576 235550 283604 311866
rect 283748 311296 283800 311302
rect 283748 311238 283800 311244
rect 283656 310004 283708 310010
rect 283656 309946 283708 309952
rect 283564 235544 283616 235550
rect 283564 235486 283616 235492
rect 283564 232688 283616 232694
rect 283564 232630 283616 232636
rect 283576 232422 283604 232630
rect 283564 232416 283616 232422
rect 283564 232358 283616 232364
rect 283576 143410 283604 232358
rect 283668 224262 283696 309946
rect 283760 231334 283788 311238
rect 284024 307896 284076 307902
rect 284024 307838 284076 307844
rect 283932 301572 283984 301578
rect 283932 301514 283984 301520
rect 283840 298104 283892 298110
rect 283840 298046 283892 298052
rect 283852 297566 283880 298046
rect 283840 297560 283892 297566
rect 283840 297502 283892 297508
rect 283748 231328 283800 231334
rect 283748 231270 283800 231276
rect 283656 224256 283708 224262
rect 283656 224198 283708 224204
rect 283852 220522 283880 297502
rect 283944 225865 283972 301514
rect 284036 233850 284064 307838
rect 284116 299056 284168 299062
rect 284116 298998 284168 299004
rect 284128 241233 284156 298998
rect 284220 298110 284248 311866
rect 284208 298104 284260 298110
rect 284208 298046 284260 298052
rect 284208 254584 284260 254590
rect 284208 254526 284260 254532
rect 284114 241224 284170 241233
rect 284114 241159 284170 241168
rect 284220 233986 284248 254526
rect 284208 233980 284260 233986
rect 284208 233922 284260 233928
rect 284024 233844 284076 233850
rect 284024 233786 284076 233792
rect 283930 225856 283986 225865
rect 283930 225791 283986 225800
rect 283840 220516 283892 220522
rect 283840 220458 283892 220464
rect 284220 219434 284248 233922
rect 284312 220658 284340 317086
rect 284404 311166 284432 317727
rect 284496 317150 284524 319194
rect 284588 318753 284616 319756
rect 284574 318744 284630 318753
rect 284574 318679 284630 318688
rect 284484 317144 284536 317150
rect 284484 317086 284536 317092
rect 284484 314560 284536 314566
rect 284484 314502 284536 314508
rect 284392 311160 284444 311166
rect 284392 311102 284444 311108
rect 284496 310978 284524 314502
rect 284404 310950 284524 310978
rect 284404 242049 284432 310950
rect 284588 296714 284616 318679
rect 284680 316470 284708 319892
rect 284772 318442 284800 319926
rect 284910 319818 284938 320076
rect 284864 319790 284938 319818
rect 284760 318436 284812 318442
rect 284760 318378 284812 318384
rect 284668 316464 284720 316470
rect 284668 316406 284720 316412
rect 284668 316328 284720 316334
rect 284668 316270 284720 316276
rect 284496 296686 284616 296714
rect 284390 242040 284446 242049
rect 284390 241975 284446 241984
rect 284392 236972 284444 236978
rect 284392 236914 284444 236920
rect 284300 220652 284352 220658
rect 284300 220594 284352 220600
rect 284128 219406 284248 219434
rect 284128 167074 284156 219406
rect 283656 167068 283708 167074
rect 283656 167010 283708 167016
rect 284116 167068 284168 167074
rect 284116 167010 284168 167016
rect 283668 158030 283696 167010
rect 283656 158024 283708 158030
rect 283656 157966 283708 157972
rect 284404 152454 284432 236914
rect 284496 220726 284524 296686
rect 284680 295089 284708 316270
rect 284864 315654 284892 319790
rect 285002 319716 285030 320076
rect 285094 319784 285122 320076
rect 286276 320104 286332 320113
rect 285172 320039 285228 320048
rect 285278 319920 285306 320076
rect 285232 319892 285306 319920
rect 285094 319756 285168 319784
rect 284956 319688 285030 319716
rect 284956 317422 284984 319688
rect 285036 319320 285088 319326
rect 285036 319262 285088 319268
rect 284944 317416 284996 317422
rect 284944 317358 284996 317364
rect 284852 315648 284904 315654
rect 284852 315590 284904 315596
rect 284760 314628 284812 314634
rect 284760 314570 284812 314576
rect 284666 295080 284722 295089
rect 284666 295015 284722 295024
rect 284680 294001 284708 295015
rect 284666 293992 284722 294001
rect 284666 293927 284722 293936
rect 284772 240961 284800 314570
rect 285048 311894 285076 319262
rect 285140 316334 285168 319756
rect 285232 319546 285260 319892
rect 285370 319784 285398 320076
rect 285554 319954 285582 320076
rect 285508 319926 285582 319954
rect 285646 319954 285674 320076
rect 285646 319926 285720 319954
rect 285508 319818 285536 319926
rect 285508 319790 285628 319818
rect 285370 319756 285444 319784
rect 285232 319518 285352 319546
rect 285220 319388 285272 319394
rect 285220 319330 285272 319336
rect 285128 316328 285180 316334
rect 285128 316270 285180 316276
rect 285232 314566 285260 319330
rect 285324 318782 285352 319518
rect 285312 318776 285364 318782
rect 285312 318718 285364 318724
rect 285416 318617 285444 319756
rect 285600 319705 285628 319790
rect 285586 319696 285642 319705
rect 285586 319631 285642 319640
rect 285600 319326 285628 319631
rect 285692 319394 285720 319926
rect 285830 319920 285858 320076
rect 285784 319892 285858 319920
rect 285680 319388 285732 319394
rect 285680 319330 285732 319336
rect 285588 319320 285640 319326
rect 285588 319262 285640 319268
rect 285402 318608 285458 318617
rect 285402 318543 285458 318552
rect 285416 317801 285444 318543
rect 285402 317792 285458 317801
rect 285402 317727 285458 317736
rect 285784 317506 285812 319892
rect 285922 319818 285950 320076
rect 285876 319790 285950 319818
rect 285876 319297 285904 319790
rect 286014 319682 286042 320076
rect 286106 319818 286134 320076
rect 287104 320104 287160 320113
rect 286276 320039 286332 320048
rect 286382 319920 286410 320076
rect 286336 319892 286410 319920
rect 286106 319790 286180 319818
rect 286014 319654 286088 319682
rect 285862 319288 285918 319297
rect 285862 319223 285918 319232
rect 286060 317898 286088 319654
rect 286152 318374 286180 319790
rect 286140 318368 286192 318374
rect 286140 318310 286192 318316
rect 286048 317892 286100 317898
rect 286048 317834 286100 317840
rect 286060 317762 286088 317834
rect 286048 317756 286100 317762
rect 286048 317698 286100 317704
rect 286336 317642 286364 319892
rect 286474 319784 286502 320076
rect 286658 319954 286686 320076
rect 285600 317478 285812 317506
rect 286060 317614 286364 317642
rect 286428 319756 286502 319784
rect 286612 319926 286686 319954
rect 285312 316464 285364 316470
rect 285312 316406 285364 316412
rect 285220 314560 285272 314566
rect 285220 314502 285272 314508
rect 284864 311866 285076 311894
rect 284864 311234 284892 311866
rect 284852 311228 284904 311234
rect 284852 311170 284904 311176
rect 285324 306374 285352 316406
rect 285600 314634 285628 317478
rect 286060 316146 286088 317614
rect 286324 317552 286376 317558
rect 286324 317494 286376 317500
rect 285876 316118 286088 316146
rect 285772 315784 285824 315790
rect 285772 315726 285824 315732
rect 285784 315382 285812 315726
rect 285772 315376 285824 315382
rect 285772 315318 285824 315324
rect 285588 314628 285640 314634
rect 285588 314570 285640 314576
rect 285048 306346 285352 306374
rect 285048 305590 285076 306346
rect 285036 305584 285088 305590
rect 285036 305526 285088 305532
rect 285048 243574 285076 305526
rect 285876 304978 285904 316118
rect 286140 315784 286192 315790
rect 286140 315726 286192 315732
rect 286048 315716 286100 315722
rect 286048 315658 286100 315664
rect 285956 314356 286008 314362
rect 285956 314298 286008 314304
rect 285968 306338 285996 314298
rect 286060 310321 286088 315658
rect 286046 310312 286102 310321
rect 286046 310247 286102 310256
rect 285956 306332 286008 306338
rect 285956 306274 286008 306280
rect 285864 304972 285916 304978
rect 285864 304914 285916 304920
rect 285310 302968 285366 302977
rect 285310 302903 285366 302912
rect 285218 302016 285274 302025
rect 285218 301951 285274 301960
rect 285126 293992 285182 294001
rect 285126 293927 285182 293936
rect 285036 243568 285088 243574
rect 285036 243510 285088 243516
rect 284758 240952 284814 240961
rect 284758 240887 284814 240896
rect 285140 239601 285168 293927
rect 285126 239592 285182 239601
rect 285126 239527 285182 239536
rect 284758 237416 284814 237425
rect 284758 237351 284814 237360
rect 284772 236978 284800 237351
rect 284760 236972 284812 236978
rect 284760 236914 284812 236920
rect 285126 233880 285182 233889
rect 285126 233815 285182 233824
rect 285036 229764 285088 229770
rect 285036 229706 285088 229712
rect 284484 220720 284536 220726
rect 284484 220662 284536 220668
rect 284392 152448 284444 152454
rect 284392 152390 284444 152396
rect 284300 147484 284352 147490
rect 284300 147426 284352 147432
rect 284312 146946 284340 147426
rect 284300 146940 284352 146946
rect 284300 146882 284352 146888
rect 284944 144832 284996 144838
rect 284944 144774 284996 144780
rect 283104 143404 283156 143410
rect 283104 143346 283156 143352
rect 283564 143404 283616 143410
rect 283564 143346 283616 143352
rect 283116 142866 283144 143346
rect 283104 142860 283156 142866
rect 283104 142802 283156 142808
rect 283012 142112 283064 142118
rect 283012 142054 283064 142060
rect 283024 137358 283052 142054
rect 283012 137352 283064 137358
rect 283012 137294 283064 137300
rect 284390 94480 284446 94489
rect 284390 94415 284446 94424
rect 282932 16546 283144 16574
rect 281908 3052 281960 3058
rect 281908 2994 281960 3000
rect 282184 3052 282236 3058
rect 282184 2994 282236 3000
rect 281920 480 281948 2994
rect 283116 480 283144 16546
rect 284404 6914 284432 94415
rect 284312 6886 284432 6914
rect 284312 480 284340 6886
rect 284956 4078 284984 144774
rect 285048 140758 285076 229706
rect 285140 146946 285168 233815
rect 285232 223009 285260 301951
rect 285324 227089 285352 302903
rect 286152 300830 286180 315726
rect 286336 311370 286364 317494
rect 286428 317218 286456 319756
rect 286612 319716 286640 319926
rect 286750 319784 286778 320076
rect 286520 319688 286640 319716
rect 286704 319756 286778 319784
rect 286416 317212 286468 317218
rect 286416 317154 286468 317160
rect 286520 314362 286548 319688
rect 286704 315790 286732 319756
rect 286842 319716 286870 320076
rect 286934 319818 286962 320076
rect 287026 319920 287054 320076
rect 288300 320104 288356 320113
rect 287104 320039 287160 320048
rect 287210 319954 287238 320076
rect 287164 319926 287238 319954
rect 287026 319892 287100 319920
rect 286934 319790 287008 319818
rect 286796 319688 286870 319716
rect 286692 315784 286744 315790
rect 286692 315726 286744 315732
rect 286796 315722 286824 319688
rect 286980 318986 287008 319790
rect 286968 318980 287020 318986
rect 286968 318922 287020 318928
rect 287072 318866 287100 319892
rect 287164 319802 287192 319926
rect 287152 319796 287204 319802
rect 287302 319784 287330 320076
rect 287152 319738 287204 319744
rect 287256 319756 287330 319784
rect 287394 319784 287422 320076
rect 287394 319756 287468 319784
rect 287164 319190 287192 319738
rect 287152 319184 287204 319190
rect 287152 319126 287204 319132
rect 286888 318838 287100 318866
rect 286784 315716 286836 315722
rect 286784 315658 286836 315664
rect 286508 314356 286560 314362
rect 286508 314298 286560 314304
rect 286888 311894 286916 318838
rect 287256 317642 287284 319756
rect 287334 319696 287390 319705
rect 287334 319631 287390 319640
rect 287348 317762 287376 319631
rect 287336 317756 287388 317762
rect 287336 317698 287388 317704
rect 286612 311866 286916 311894
rect 286980 317614 287284 317642
rect 286324 311364 286376 311370
rect 286324 311306 286376 311312
rect 286416 311364 286468 311370
rect 286416 311306 286468 311312
rect 286324 303476 286376 303482
rect 286324 303418 286376 303424
rect 286140 300824 286192 300830
rect 286140 300766 286192 300772
rect 285772 240100 285824 240106
rect 285772 240042 285824 240048
rect 285784 239358 285812 240042
rect 285772 239352 285824 239358
rect 285772 239294 285824 239300
rect 285588 236020 285640 236026
rect 285588 235962 285640 235968
rect 285600 235498 285628 235962
rect 285680 235884 285732 235890
rect 285680 235826 285732 235832
rect 285692 235618 285720 235826
rect 285680 235612 285732 235618
rect 285680 235554 285732 235560
rect 285600 235470 285720 235498
rect 285310 227080 285366 227089
rect 285310 227015 285366 227024
rect 285218 223000 285274 223009
rect 285218 222935 285274 222944
rect 285128 146940 285180 146946
rect 285128 146882 285180 146888
rect 285036 140752 285088 140758
rect 285036 140694 285088 140700
rect 285048 140146 285076 140694
rect 285036 140140 285088 140146
rect 285036 140082 285088 140088
rect 285692 133890 285720 235470
rect 285784 137970 285812 239294
rect 286336 224194 286364 303418
rect 286428 232830 286456 311306
rect 286506 309768 286562 309777
rect 286506 309703 286562 309712
rect 286520 234598 286548 309703
rect 286612 301646 286640 311866
rect 286784 308372 286836 308378
rect 286784 308314 286836 308320
rect 286692 304292 286744 304298
rect 286692 304234 286744 304240
rect 286600 301640 286652 301646
rect 286600 301582 286652 301588
rect 286598 295216 286654 295225
rect 286598 295151 286654 295160
rect 286508 234592 286560 234598
rect 286508 234534 286560 234540
rect 286416 232824 286468 232830
rect 286416 232766 286468 232772
rect 286324 224188 286376 224194
rect 286324 224130 286376 224136
rect 286612 220590 286640 295151
rect 286704 231169 286732 304234
rect 286796 240106 286824 308314
rect 286980 306374 287008 317614
rect 287152 317484 287204 317490
rect 287152 317426 287204 317432
rect 287060 316328 287112 316334
rect 287060 316270 287112 316276
rect 287072 313274 287100 316270
rect 287060 313268 287112 313274
rect 287060 313210 287112 313216
rect 287164 311894 287192 317426
rect 287440 316010 287468 319756
rect 287578 319716 287606 320076
rect 287670 319784 287698 320076
rect 287854 319852 287882 320076
rect 287808 319824 287882 319852
rect 287670 319756 287744 319784
rect 287578 319688 287652 319716
rect 287520 319388 287572 319394
rect 287520 319330 287572 319336
rect 287532 316334 287560 319330
rect 287520 316328 287572 316334
rect 287520 316270 287572 316276
rect 287440 315982 287560 316010
rect 287336 315784 287388 315790
rect 287336 315726 287388 315732
rect 287244 315716 287296 315722
rect 287244 315658 287296 315664
rect 287072 311866 287192 311894
rect 287072 310146 287100 311866
rect 287060 310140 287112 310146
rect 287060 310082 287112 310088
rect 286888 306346 287008 306374
rect 286888 295225 286916 306346
rect 286968 300144 287020 300150
rect 286968 300086 287020 300092
rect 286874 295216 286930 295225
rect 286874 295151 286930 295160
rect 286876 253224 286928 253230
rect 286876 253166 286928 253172
rect 286784 240100 286836 240106
rect 286784 240042 286836 240048
rect 286888 237250 286916 253166
rect 286876 237244 286928 237250
rect 286876 237186 286928 237192
rect 286888 236026 286916 237186
rect 286876 236020 286928 236026
rect 286876 235962 286928 235968
rect 286980 235890 287008 300086
rect 287256 299033 287284 315658
rect 287348 302190 287376 315726
rect 287428 315648 287480 315654
rect 287428 315590 287480 315596
rect 287440 303618 287468 315590
rect 287532 305522 287560 315982
rect 287520 305516 287572 305522
rect 287520 305458 287572 305464
rect 287532 305046 287560 305458
rect 287520 305040 287572 305046
rect 287520 304982 287572 304988
rect 287428 303612 287480 303618
rect 287428 303554 287480 303560
rect 287336 302184 287388 302190
rect 287336 302126 287388 302132
rect 287242 299024 287298 299033
rect 287242 298959 287298 298968
rect 287624 295186 287652 319688
rect 287716 319410 287744 319756
rect 287808 319705 287836 319824
rect 287946 319784 287974 320076
rect 287900 319756 287974 319784
rect 288038 319784 288066 320076
rect 288130 319920 288158 320076
rect 288576 320104 288632 320113
rect 288300 320039 288356 320048
rect 288130 319892 288204 319920
rect 288038 319756 288112 319784
rect 287794 319696 287850 319705
rect 287794 319631 287850 319640
rect 287716 319382 287836 319410
rect 287702 319288 287758 319297
rect 287702 319223 287758 319232
rect 287716 315790 287744 319223
rect 287808 316334 287836 319382
rect 287796 316328 287848 316334
rect 287796 316270 287848 316276
rect 287704 315784 287756 315790
rect 287704 315726 287756 315732
rect 287796 315784 287848 315790
rect 287796 315726 287848 315732
rect 287808 307766 287836 315726
rect 287900 315722 287928 319756
rect 287978 319696 288034 319705
rect 287978 319631 288034 319640
rect 287992 319394 288020 319631
rect 287980 319388 288032 319394
rect 287980 319330 288032 319336
rect 288084 318306 288112 319756
rect 288176 318714 288204 319892
rect 288406 319852 288434 320076
rect 288254 319832 288310 319841
rect 288254 319767 288310 319776
rect 288360 319824 288434 319852
rect 288498 319852 288526 320076
rect 288944 320104 289000 320113
rect 288576 320039 288632 320048
rect 288774 319920 288802 320076
rect 288728 319892 288802 319920
rect 288866 319920 288894 320076
rect 289312 320104 289368 320113
rect 288944 320039 289000 320048
rect 289050 319938 289078 320076
rect 289038 319932 289090 319938
rect 288866 319892 288940 319920
rect 288498 319824 288572 319852
rect 288164 318708 288216 318714
rect 288164 318650 288216 318656
rect 288072 318300 288124 318306
rect 288072 318242 288124 318248
rect 288268 317914 288296 319767
rect 288084 317886 288296 317914
rect 287980 316328 288032 316334
rect 287980 316270 288032 316276
rect 287888 315716 287940 315722
rect 287888 315658 287940 315664
rect 287888 310412 287940 310418
rect 287888 310354 287940 310360
rect 287796 307760 287848 307766
rect 287796 307702 287848 307708
rect 287796 305040 287848 305046
rect 287796 304982 287848 304988
rect 287704 299124 287756 299130
rect 287704 299066 287756 299072
rect 287612 295180 287664 295186
rect 287612 295122 287664 295128
rect 287624 294370 287652 295122
rect 287612 294364 287664 294370
rect 287612 294306 287664 294312
rect 287716 240854 287744 299066
rect 287808 296041 287836 304982
rect 287794 296032 287850 296041
rect 287794 295967 287850 295976
rect 287704 240848 287756 240854
rect 287704 240790 287756 240796
rect 287796 240508 287848 240514
rect 287796 240450 287848 240456
rect 286968 235884 287020 235890
rect 286968 235826 287020 235832
rect 287704 235884 287756 235890
rect 287704 235826 287756 235832
rect 286690 231160 286746 231169
rect 286690 231095 286746 231104
rect 286600 220584 286652 220590
rect 286600 220526 286652 220532
rect 285772 137964 285824 137970
rect 285772 137906 285824 137912
rect 285784 137290 285812 137906
rect 285772 137284 285824 137290
rect 285772 137226 285824 137232
rect 285680 133884 285732 133890
rect 285680 133826 285732 133832
rect 285692 133278 285720 133826
rect 285680 133272 285732 133278
rect 285680 133214 285732 133220
rect 287058 26888 287114 26897
rect 287058 26823 287114 26832
rect 287072 16574 287100 26823
rect 287072 16546 287376 16574
rect 284944 4072 284996 4078
rect 284944 4014 284996 4020
rect 286600 3800 286652 3806
rect 286600 3742 286652 3748
rect 285404 3052 285456 3058
rect 285404 2994 285456 3000
rect 285416 480 285444 2994
rect 286612 480 286640 3742
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287348 354 287376 16546
rect 287716 3126 287744 235826
rect 287808 132462 287836 240450
rect 287900 221678 287928 310354
rect 287992 296682 288020 316270
rect 288084 315654 288112 317886
rect 288256 317756 288308 317762
rect 288256 317698 288308 317704
rect 288162 315752 288218 315761
rect 288162 315687 288218 315696
rect 288072 315648 288124 315654
rect 288072 315590 288124 315596
rect 288176 314945 288204 315687
rect 288162 314936 288218 314945
rect 288162 314871 288218 314880
rect 288268 312662 288296 317698
rect 288360 315790 288388 319824
rect 288544 319546 288572 319824
rect 288728 319682 288756 319892
rect 288912 319818 288940 319892
rect 289038 319874 289090 319880
rect 288912 319790 289032 319818
rect 288452 319518 288572 319546
rect 288636 319654 288756 319682
rect 288808 319728 288860 319734
rect 288808 319670 288860 319676
rect 288348 315784 288400 315790
rect 288348 315726 288400 315732
rect 288256 312656 288308 312662
rect 288256 312598 288308 312604
rect 288452 310457 288480 319518
rect 288636 319410 288664 319654
rect 288544 319382 288664 319410
rect 288544 317966 288572 319382
rect 288622 319288 288678 319297
rect 288622 319223 288678 319232
rect 288532 317960 288584 317966
rect 288532 317902 288584 317908
rect 288636 316010 288664 319223
rect 288714 319152 288770 319161
rect 288714 319087 288770 319096
rect 288544 315982 288664 316010
rect 288544 311846 288572 315982
rect 288728 315874 288756 319087
rect 288636 315846 288756 315874
rect 288532 311840 288584 311846
rect 288532 311782 288584 311788
rect 288636 311778 288664 315846
rect 288716 314288 288768 314294
rect 288716 314230 288768 314236
rect 288624 311772 288676 311778
rect 288624 311714 288676 311720
rect 288438 310448 288494 310457
rect 288438 310383 288494 310392
rect 288164 304428 288216 304434
rect 288164 304370 288216 304376
rect 288072 303340 288124 303346
rect 288072 303282 288124 303288
rect 287980 296676 288032 296682
rect 287980 296618 288032 296624
rect 287992 296313 288020 296618
rect 287978 296304 288034 296313
rect 287978 296239 288034 296248
rect 287980 240848 288032 240854
rect 287980 240790 288032 240796
rect 287992 240514 288020 240790
rect 287980 240508 288032 240514
rect 287980 240450 288032 240456
rect 287980 236700 288032 236706
rect 287980 236642 288032 236648
rect 287888 221672 287940 221678
rect 287888 221614 287940 221620
rect 287992 153134 288020 236642
rect 288084 224466 288112 303282
rect 288176 228274 288204 304370
rect 288348 303272 288400 303278
rect 288348 303214 288400 303220
rect 288256 299396 288308 299402
rect 288256 299338 288308 299344
rect 288268 299033 288296 299338
rect 288254 299024 288310 299033
rect 288254 298959 288310 298968
rect 288256 294364 288308 294370
rect 288256 294306 288308 294312
rect 288164 228268 288216 228274
rect 288164 228210 288216 228216
rect 288072 224460 288124 224466
rect 288072 224402 288124 224408
rect 288268 220794 288296 294306
rect 288360 230110 288388 303214
rect 288728 299470 288756 314230
rect 288820 301646 288848 319670
rect 288900 319388 288952 319394
rect 288900 319330 288952 319336
rect 288808 301640 288860 301646
rect 288808 301582 288860 301588
rect 288716 299464 288768 299470
rect 288716 299406 288768 299412
rect 288624 298104 288676 298110
rect 288624 298046 288676 298052
rect 288636 296750 288664 298046
rect 288624 296744 288676 296750
rect 288624 296686 288676 296692
rect 288636 295254 288664 296686
rect 288912 295322 288940 319330
rect 289004 319122 289032 319790
rect 289142 319716 289170 320076
rect 289234 319784 289262 320076
rect 289680 320104 289736 320113
rect 289312 320039 289368 320048
rect 289418 319818 289446 320076
rect 289372 319790 289446 319818
rect 289602 319818 289630 320076
rect 289864 320104 289920 320113
rect 289680 320039 289736 320048
rect 289786 319920 289814 320076
rect 290416 320104 290472 320113
rect 289864 320039 289920 320048
rect 289786 319892 289860 319920
rect 289726 319832 289782 319841
rect 289602 319790 289676 319818
rect 289234 319756 289308 319784
rect 289096 319688 289170 319716
rect 288992 319116 289044 319122
rect 288992 319058 289044 319064
rect 289096 314294 289124 319688
rect 289174 317520 289230 317529
rect 289174 317455 289230 317464
rect 289084 314288 289136 314294
rect 289084 314230 289136 314236
rect 289188 311894 289216 317455
rect 289280 315790 289308 319756
rect 289372 317393 289400 319790
rect 289450 319696 289506 319705
rect 289450 319631 289506 319640
rect 289358 317384 289414 317393
rect 289358 317319 289414 317328
rect 289268 315784 289320 315790
rect 289268 315726 289320 315732
rect 289096 311866 289216 311894
rect 288900 295316 288952 295322
rect 288900 295258 288952 295264
rect 288624 295248 288676 295254
rect 288624 295190 288676 295196
rect 288912 294953 288940 295258
rect 288898 294944 288954 294953
rect 288898 294879 288954 294888
rect 288992 246356 289044 246362
rect 288992 246298 289044 246304
rect 288440 241460 288492 241466
rect 288440 241402 288492 241408
rect 288452 240310 288480 241402
rect 288440 240304 288492 240310
rect 288440 240246 288492 240252
rect 288348 230104 288400 230110
rect 288348 230046 288400 230052
rect 288256 220788 288308 220794
rect 288256 220730 288308 220736
rect 287980 153128 288032 153134
rect 287980 153070 288032 153076
rect 288348 153128 288400 153134
rect 288348 153070 288400 153076
rect 288360 152522 288388 153070
rect 288348 152516 288400 152522
rect 288348 152458 288400 152464
rect 287796 132456 287848 132462
rect 287796 132398 287848 132404
rect 287808 131850 287836 132398
rect 287796 131844 287848 131850
rect 287796 131786 287848 131792
rect 288452 126886 288480 240246
rect 289004 237454 289032 246298
rect 288532 237448 288584 237454
rect 288532 237390 288584 237396
rect 288992 237448 289044 237454
rect 288992 237390 289044 237396
rect 288544 156670 288572 237390
rect 289096 223038 289124 311866
rect 289268 311500 289320 311506
rect 289268 311442 289320 311448
rect 289174 310856 289230 310865
rect 289174 310791 289230 310800
rect 289188 239465 289216 310791
rect 289174 239456 289230 239465
rect 289174 239391 289230 239400
rect 289176 230988 289228 230994
rect 289176 230930 289228 230936
rect 289084 223032 289136 223038
rect 289084 222974 289136 222980
rect 289084 156732 289136 156738
rect 289084 156674 289136 156680
rect 288532 156664 288584 156670
rect 288532 156606 288584 156612
rect 288440 126880 288492 126886
rect 288440 126822 288492 126828
rect 288992 4004 289044 4010
rect 288992 3946 289044 3952
rect 287704 3120 287756 3126
rect 287704 3062 287756 3068
rect 289004 480 289032 3946
rect 289096 3058 289124 156674
rect 289188 142050 289216 230930
rect 289280 225486 289308 311442
rect 289360 299464 289412 299470
rect 289360 299406 289412 299412
rect 289372 299198 289400 299406
rect 289464 299266 289492 319631
rect 289648 318345 289676 319790
rect 289726 319767 289782 319776
rect 289634 318336 289690 318345
rect 289634 318271 289690 318280
rect 289740 317422 289768 319767
rect 289832 319394 289860 319892
rect 289970 319784 289998 320076
rect 290154 319954 290182 320076
rect 289924 319756 289998 319784
rect 290108 319926 290182 319954
rect 289820 319388 289872 319394
rect 289820 319330 289872 319336
rect 289924 318238 289952 319756
rect 290004 319320 290056 319326
rect 290004 319262 290056 319268
rect 289912 318232 289964 318238
rect 289912 318174 289964 318180
rect 289728 317416 289780 317422
rect 289728 317358 289780 317364
rect 289728 315784 289780 315790
rect 289728 315726 289780 315732
rect 289636 301640 289688 301646
rect 289636 301582 289688 301588
rect 289452 299260 289504 299266
rect 289452 299202 289504 299208
rect 289360 299192 289412 299198
rect 289360 299134 289412 299140
rect 289372 238950 289400 299134
rect 289360 238944 289412 238950
rect 289360 238886 289412 238892
rect 289360 236020 289412 236026
rect 289360 235962 289412 235968
rect 289268 225480 289320 225486
rect 289268 225422 289320 225428
rect 289372 155990 289400 235962
rect 289464 219434 289492 299202
rect 289544 297696 289596 297702
rect 289544 297638 289596 297644
rect 289452 219428 289504 219434
rect 289452 219370 289504 219376
rect 289556 219162 289584 297638
rect 289648 294545 289676 301582
rect 289740 298110 289768 315726
rect 290016 311545 290044 319262
rect 290108 318345 290136 319926
rect 290246 319784 290274 320076
rect 290338 319818 290366 320076
rect 290876 320104 290932 320113
rect 290416 320039 290472 320048
rect 290522 319920 290550 320076
rect 290706 319954 290734 320076
rect 290660 319926 290734 319954
rect 290522 319892 290596 319920
rect 290462 319832 290518 319841
rect 290338 319790 290412 319818
rect 290200 319756 290274 319784
rect 290094 318336 290150 318345
rect 290094 318271 290150 318280
rect 290108 317529 290136 318271
rect 290200 317694 290228 319756
rect 290278 319696 290334 319705
rect 290278 319631 290334 319640
rect 290292 317694 290320 319631
rect 290384 319326 290412 319790
rect 290462 319767 290518 319776
rect 290372 319320 290424 319326
rect 290372 319262 290424 319268
rect 290476 318714 290504 319767
rect 290464 318708 290516 318714
rect 290464 318650 290516 318656
rect 290372 318504 290424 318510
rect 290372 318446 290424 318452
rect 290188 317688 290240 317694
rect 290188 317630 290240 317636
rect 290280 317688 290332 317694
rect 290280 317630 290332 317636
rect 290094 317520 290150 317529
rect 290094 317455 290150 317464
rect 290096 317416 290148 317422
rect 290096 317358 290148 317364
rect 290002 311536 290058 311545
rect 290002 311471 290058 311480
rect 290108 299062 290136 317358
rect 290292 315790 290320 317630
rect 290280 315784 290332 315790
rect 290280 315726 290332 315732
rect 290384 311894 290412 318446
rect 290476 315738 290504 318650
rect 290568 318322 290596 319892
rect 290660 318646 290688 319926
rect 290798 319784 290826 320076
rect 291428 320104 291484 320113
rect 290876 320039 290932 320048
rect 290982 319784 291010 320076
rect 291074 319852 291102 320076
rect 291074 319824 291148 319852
rect 290798 319756 290872 319784
rect 290982 319756 291056 319784
rect 290844 319410 290872 319756
rect 291028 319512 291056 319756
rect 291120 319705 291148 319824
rect 291258 319784 291286 320076
rect 291212 319756 291286 319784
rect 291350 319784 291378 320076
rect 292164 320104 292220 320113
rect 291428 320039 291484 320048
rect 291534 319852 291562 320076
rect 291488 319824 291562 319852
rect 291350 319756 291424 319784
rect 291106 319696 291162 319705
rect 291106 319631 291162 319640
rect 291028 319484 291148 319512
rect 290844 319382 290964 319410
rect 290936 319376 290964 319382
rect 290936 319348 291010 319376
rect 290982 319274 291010 319348
rect 290936 319246 291010 319274
rect 290738 319152 290794 319161
rect 290738 319087 290794 319096
rect 290648 318640 290700 318646
rect 290648 318582 290700 318588
rect 290660 318510 290688 318582
rect 290648 318504 290700 318510
rect 290648 318446 290700 318452
rect 290568 318294 290688 318322
rect 290556 318164 290608 318170
rect 290556 318106 290608 318112
rect 290568 315874 290596 318106
rect 290660 316010 290688 318294
rect 290752 316849 290780 319087
rect 290830 318880 290886 318889
rect 290830 318815 290886 318824
rect 290844 317558 290872 318815
rect 290832 317552 290884 317558
rect 290832 317494 290884 317500
rect 290738 316840 290794 316849
rect 290738 316775 290794 316784
rect 290660 315982 290872 316010
rect 290568 315846 290780 315874
rect 290648 315784 290700 315790
rect 290476 315710 290596 315738
rect 290648 315726 290700 315732
rect 290384 311866 290504 311894
rect 290096 299056 290148 299062
rect 290096 298998 290148 299004
rect 289728 298104 289780 298110
rect 289728 298046 289780 298052
rect 289634 294536 289690 294545
rect 289634 294471 289690 294480
rect 289636 271176 289688 271182
rect 289636 271118 289688 271124
rect 289648 241466 289676 271118
rect 289728 253292 289780 253298
rect 289728 253234 289780 253240
rect 289636 241460 289688 241466
rect 289636 241402 289688 241408
rect 289740 237114 289768 253234
rect 289728 237108 289780 237114
rect 289728 237050 289780 237056
rect 289740 236026 289768 237050
rect 289728 236020 289780 236026
rect 289728 235962 289780 235968
rect 289728 231260 289780 231266
rect 289728 231202 289780 231208
rect 289740 230994 289768 231202
rect 289728 230988 289780 230994
rect 289728 230930 289780 230936
rect 290476 219366 290504 311866
rect 290568 220833 290596 315710
rect 290660 248033 290688 315726
rect 290752 257446 290780 315846
rect 290844 298858 290872 315982
rect 290936 299130 290964 319246
rect 291014 318880 291070 318889
rect 291014 318815 291070 318824
rect 291028 317490 291056 318815
rect 291120 318170 291148 319484
rect 291108 318164 291160 318170
rect 291108 318106 291160 318112
rect 291212 317694 291240 319756
rect 291292 319388 291344 319394
rect 291292 319330 291344 319336
rect 291304 318374 291332 319330
rect 291292 318368 291344 318374
rect 291292 318310 291344 318316
rect 291108 317688 291160 317694
rect 291108 317630 291160 317636
rect 291200 317688 291252 317694
rect 291200 317630 291252 317636
rect 291120 317490 291148 317630
rect 291200 317552 291252 317558
rect 291200 317494 291252 317500
rect 291016 317484 291068 317490
rect 291016 317426 291068 317432
rect 291108 317484 291160 317490
rect 291108 317426 291160 317432
rect 291212 315874 291240 317494
rect 291120 315846 291240 315874
rect 291120 315466 291148 315846
rect 291292 315784 291344 315790
rect 291198 315752 291254 315761
rect 291292 315726 291344 315732
rect 291198 315687 291254 315696
rect 291212 315586 291240 315687
rect 291200 315580 291252 315586
rect 291200 315522 291252 315528
rect 291120 315438 291240 315466
rect 291106 310448 291162 310457
rect 291106 310383 291162 310392
rect 291120 300830 291148 310383
rect 291108 300824 291160 300830
rect 291108 300766 291160 300772
rect 290924 299124 290976 299130
rect 290924 299066 290976 299072
rect 290832 298852 290884 298858
rect 290832 298794 290884 298800
rect 290740 257440 290792 257446
rect 290740 257382 290792 257388
rect 290646 248024 290702 248033
rect 290646 247959 290702 247968
rect 291120 235754 291148 300766
rect 291212 280838 291240 315438
rect 291304 298110 291332 315726
rect 291396 301889 291424 319756
rect 291488 318306 291516 319824
rect 291626 319784 291654 320076
rect 291810 319954 291838 320076
rect 291580 319756 291654 319784
rect 291764 319926 291838 319954
rect 291476 318300 291528 318306
rect 291476 318242 291528 318248
rect 291580 315790 291608 319756
rect 291660 318776 291712 318782
rect 291660 318718 291712 318724
rect 291568 315784 291620 315790
rect 291568 315726 291620 315732
rect 291476 315716 291528 315722
rect 291476 315658 291528 315664
rect 291488 305318 291516 315658
rect 291568 315648 291620 315654
rect 291568 315590 291620 315596
rect 291580 306270 291608 315590
rect 291568 306264 291620 306270
rect 291568 306206 291620 306212
rect 291580 305862 291608 306206
rect 291568 305856 291620 305862
rect 291568 305798 291620 305804
rect 291476 305312 291528 305318
rect 291476 305254 291528 305260
rect 291382 301880 291438 301889
rect 291382 301815 291438 301824
rect 291292 298104 291344 298110
rect 291292 298046 291344 298052
rect 291672 295118 291700 318718
rect 291764 318510 291792 319926
rect 291994 319852 292022 320076
rect 291948 319824 292022 319852
rect 291842 319288 291898 319297
rect 291842 319223 291898 319232
rect 291752 318504 291804 318510
rect 291752 318446 291804 318452
rect 291752 318368 291804 318374
rect 291752 318310 291804 318316
rect 291660 295112 291712 295118
rect 291660 295054 291712 295060
rect 291672 294409 291700 295054
rect 291658 294400 291714 294409
rect 291658 294335 291714 294344
rect 291200 280832 291252 280838
rect 291200 280774 291252 280780
rect 291764 279478 291792 318310
rect 291856 317801 291884 319223
rect 291948 318782 291976 319824
rect 292086 319784 292114 320076
rect 293452 320104 293508 320113
rect 292164 320039 292220 320048
rect 292270 319920 292298 320076
rect 292454 319920 292482 320076
rect 292040 319756 292114 319784
rect 292224 319892 292298 319920
rect 292408 319892 292482 319920
rect 292040 319394 292068 319756
rect 292118 319696 292174 319705
rect 292118 319631 292174 319640
rect 292028 319388 292080 319394
rect 292028 319330 292080 319336
rect 291936 318776 291988 318782
rect 291936 318718 291988 318724
rect 291936 318504 291988 318510
rect 291936 318446 291988 318452
rect 291842 317792 291898 317801
rect 291842 317727 291898 317736
rect 291948 317558 291976 318446
rect 292026 318200 292082 318209
rect 292026 318135 292082 318144
rect 291936 317552 291988 317558
rect 291936 317494 291988 317500
rect 292040 315382 292068 318135
rect 292132 318102 292160 319631
rect 292120 318096 292172 318102
rect 292120 318038 292172 318044
rect 292224 315654 292252 319892
rect 292408 319818 292436 319892
rect 292316 319790 292436 319818
rect 292316 318578 292344 319790
rect 292546 319784 292574 320076
rect 292730 319818 292758 320076
rect 292730 319790 292804 319818
rect 292546 319756 292620 319784
rect 292486 319696 292542 319705
rect 292486 319631 292488 319640
rect 292540 319631 292542 319640
rect 292488 319602 292540 319608
rect 292592 318794 292620 319756
rect 292672 319660 292724 319666
rect 292672 319602 292724 319608
rect 292684 319569 292712 319602
rect 292670 319560 292726 319569
rect 292670 319495 292726 319504
rect 292776 319326 292804 319790
rect 292914 319784 292942 320076
rect 292868 319756 292942 319784
rect 293006 319784 293034 320076
rect 293098 319852 293126 320076
rect 293282 319943 293310 320076
rect 293268 319934 293324 319943
rect 293268 319869 293324 319878
rect 293098 319824 293172 319852
rect 293006 319756 293080 319784
rect 292764 319320 292816 319326
rect 292764 319262 292816 319268
rect 292776 319054 292804 319262
rect 292764 319048 292816 319054
rect 292764 318990 292816 318996
rect 292408 318766 292620 318794
rect 292304 318572 292356 318578
rect 292304 318514 292356 318520
rect 292304 317688 292356 317694
rect 292304 317630 292356 317636
rect 292212 315648 292264 315654
rect 292212 315590 292264 315596
rect 292028 315376 292080 315382
rect 292028 315318 292080 315324
rect 292316 311894 292344 317630
rect 292408 315722 292436 318766
rect 292488 318300 292540 318306
rect 292488 318242 292540 318248
rect 292396 315716 292448 315722
rect 292396 315658 292448 315664
rect 292224 311866 292344 311894
rect 291844 310208 291896 310214
rect 291844 310150 291896 310156
rect 291856 309806 291884 310150
rect 291844 309800 291896 309806
rect 291844 309742 291896 309748
rect 292028 305312 292080 305318
rect 292028 305254 292080 305260
rect 291936 305040 291988 305046
rect 291936 304982 291988 304988
rect 291752 279472 291804 279478
rect 291752 279414 291804 279420
rect 291108 235748 291160 235754
rect 291108 235690 291160 235696
rect 291120 234666 291148 235690
rect 291108 234660 291160 234666
rect 291108 234602 291160 234608
rect 291844 234660 291896 234666
rect 291844 234602 291896 234608
rect 290648 231192 290700 231198
rect 290648 231134 290700 231140
rect 290554 220824 290610 220833
rect 290554 220759 290610 220768
rect 290464 219360 290516 219366
rect 290464 219302 290516 219308
rect 289544 219156 289596 219162
rect 289544 219098 289596 219104
rect 289360 155984 289412 155990
rect 289360 155926 289412 155932
rect 289372 146198 289400 155926
rect 289360 146192 289412 146198
rect 289360 146134 289412 146140
rect 290660 144158 290688 231134
rect 291752 227180 291804 227186
rect 291752 227122 291804 227128
rect 291764 227050 291792 227122
rect 291752 227044 291804 227050
rect 291752 226986 291804 226992
rect 290924 144288 290976 144294
rect 290924 144230 290976 144236
rect 290936 144158 290964 144230
rect 290648 144152 290700 144158
rect 290648 144094 290700 144100
rect 290924 144152 290976 144158
rect 290924 144094 290976 144100
rect 289176 142044 289228 142050
rect 289176 141986 289228 141992
rect 289188 141506 289216 141986
rect 289176 141500 289228 141506
rect 289176 141442 289228 141448
rect 289728 126880 289780 126886
rect 289728 126822 289780 126828
rect 289740 126274 289768 126822
rect 289728 126268 289780 126274
rect 289728 126210 289780 126216
rect 291384 3732 291436 3738
rect 291384 3674 291436 3680
rect 290188 3120 290240 3126
rect 290188 3062 290240 3068
rect 289084 3052 289136 3058
rect 289084 2994 289136 3000
rect 290200 480 290228 3062
rect 291396 480 291424 3674
rect 291856 2922 291884 234602
rect 291948 228342 291976 304982
rect 291936 228336 291988 228342
rect 291936 228278 291988 228284
rect 291936 227112 291988 227118
rect 291936 227054 291988 227060
rect 291948 133822 291976 227054
rect 292040 224738 292068 305254
rect 292118 301880 292174 301889
rect 292118 301815 292174 301824
rect 292028 224732 292080 224738
rect 292028 224674 292080 224680
rect 292132 220561 292160 301815
rect 292224 246430 292252 311866
rect 292394 300248 292450 300257
rect 292394 300183 292450 300192
rect 292304 298104 292356 298110
rect 292304 298046 292356 298052
rect 292316 297498 292344 298046
rect 292304 297492 292356 297498
rect 292304 297434 292356 297440
rect 292212 246424 292264 246430
rect 292212 246366 292264 246372
rect 292212 227180 292264 227186
rect 292212 227122 292264 227128
rect 292118 220552 292174 220561
rect 292118 220487 292174 220496
rect 292224 150414 292252 227122
rect 292316 220697 292344 297434
rect 292408 225554 292436 300183
rect 292500 253366 292528 318242
rect 292580 318096 292632 318102
rect 292580 318038 292632 318044
rect 292592 314022 292620 318038
rect 292868 316860 292896 319756
rect 293052 319705 293080 319756
rect 293038 319696 293094 319705
rect 293038 319631 293094 319640
rect 293144 319530 293172 319824
rect 293374 319784 293402 320076
rect 294280 320104 294336 320113
rect 293452 320039 293508 320048
rect 293558 319954 293586 320076
rect 293512 319926 293586 319954
rect 293512 319802 293540 319926
rect 293328 319756 293402 319784
rect 293500 319796 293552 319802
rect 293132 319524 293184 319530
rect 293132 319466 293184 319472
rect 292948 319048 293000 319054
rect 292948 318990 293000 318996
rect 292960 318850 292988 318990
rect 292948 318844 293000 318850
rect 292948 318786 293000 318792
rect 292684 316832 292896 316860
rect 292684 314537 292712 316832
rect 292764 316328 292816 316334
rect 292764 316270 292816 316276
rect 292776 316062 292804 316270
rect 292764 316056 292816 316062
rect 292764 315998 292816 316004
rect 293224 315648 293276 315654
rect 293224 315590 293276 315596
rect 293132 315376 293184 315382
rect 293132 315318 293184 315324
rect 292764 315308 292816 315314
rect 292764 315250 292816 315256
rect 292670 314528 292726 314537
rect 292670 314463 292726 314472
rect 292580 314016 292632 314022
rect 292580 313958 292632 313964
rect 292776 309126 292804 315250
rect 292764 309120 292816 309126
rect 292764 309062 292816 309068
rect 293144 301578 293172 315318
rect 293236 311166 293264 315590
rect 293328 315314 293356 319756
rect 293500 319738 293552 319744
rect 293650 319716 293678 320076
rect 293834 319852 293862 320076
rect 293788 319824 293862 319852
rect 293926 319852 293954 320076
rect 294110 319954 294138 320076
rect 294464 320104 294520 320113
rect 294280 320039 294336 320048
rect 294064 319926 294138 319954
rect 293926 319824 294000 319852
rect 293650 319688 293724 319716
rect 293590 319560 293646 319569
rect 293590 319495 293646 319504
rect 293604 318850 293632 319495
rect 293592 318844 293644 318850
rect 293592 318786 293644 318792
rect 293500 317688 293552 317694
rect 293500 317630 293552 317636
rect 293316 315308 293368 315314
rect 293316 315250 293368 315256
rect 293512 314226 293540 317630
rect 293500 314220 293552 314226
rect 293500 314162 293552 314168
rect 293224 311160 293276 311166
rect 293224 311102 293276 311108
rect 293132 301572 293184 301578
rect 293132 301514 293184 301520
rect 292488 253360 292540 253366
rect 292488 253302 292540 253308
rect 293236 231742 293264 311102
rect 293408 308780 293460 308786
rect 293408 308722 293460 308728
rect 293316 297084 293368 297090
rect 293316 297026 293368 297032
rect 293224 231736 293276 231742
rect 293224 231678 293276 231684
rect 292580 227248 292632 227254
rect 292580 227190 292632 227196
rect 292592 227050 292620 227190
rect 292580 227044 292632 227050
rect 292580 226986 292632 226992
rect 293224 227044 293276 227050
rect 293224 226986 293276 226992
rect 292396 225548 292448 225554
rect 292396 225490 292448 225496
rect 292302 220688 292358 220697
rect 292302 220623 292358 220632
rect 292212 150408 292264 150414
rect 292212 150350 292264 150356
rect 292224 149734 292252 150350
rect 292212 149728 292264 149734
rect 292212 149670 292264 149676
rect 291936 133816 291988 133822
rect 291936 133758 291988 133764
rect 291948 133210 291976 133758
rect 291936 133204 291988 133210
rect 291936 133146 291988 133152
rect 293236 132394 293264 226986
rect 293328 218657 293356 297026
rect 293420 232762 293448 308722
rect 293604 239766 293632 318786
rect 293696 317626 293724 319688
rect 293684 317620 293736 317626
rect 293684 317562 293736 317568
rect 293682 317520 293738 317529
rect 293682 317455 293738 317464
rect 293696 315518 293724 317455
rect 293788 315654 293816 319824
rect 293776 315648 293828 315654
rect 293776 315590 293828 315596
rect 293684 315512 293736 315518
rect 293684 315454 293736 315460
rect 293776 315512 293828 315518
rect 293776 315454 293828 315460
rect 293684 313540 293736 313546
rect 293684 313482 293736 313488
rect 293696 313342 293724 313482
rect 293684 313336 293736 313342
rect 293684 313278 293736 313284
rect 293788 298110 293816 315454
rect 293972 315382 294000 319824
rect 293960 315376 294012 315382
rect 293960 315318 294012 315324
rect 293866 313712 293922 313721
rect 293866 313647 293922 313656
rect 293880 313478 293908 313647
rect 293868 313472 293920 313478
rect 293868 313414 293920 313420
rect 293868 313336 293920 313342
rect 293868 313278 293920 313284
rect 293776 298104 293828 298110
rect 293776 298046 293828 298052
rect 293788 297090 293816 298046
rect 293776 297084 293828 297090
rect 293776 297026 293828 297032
rect 293592 239760 293644 239766
rect 293592 239702 293644 239708
rect 293880 239426 293908 313278
rect 294064 304910 294092 319926
rect 294386 319920 294414 320076
rect 294740 320104 294796 320113
rect 294464 320039 294520 320048
rect 294340 319892 294414 319920
rect 294512 319932 294564 319938
rect 294142 319832 294198 319841
rect 294142 319767 294198 319776
rect 294156 319297 294184 319767
rect 294142 319288 294198 319297
rect 294142 319223 294198 319232
rect 294156 315450 294184 319223
rect 294234 318472 294290 318481
rect 294234 318407 294290 318416
rect 294248 317694 294276 318407
rect 294236 317688 294288 317694
rect 294236 317630 294288 317636
rect 294340 316402 294368 319892
rect 294662 319920 294690 320076
rect 296120 320104 296176 320113
rect 294740 320039 294796 320048
rect 294662 319892 294736 319920
rect 294512 319874 294564 319880
rect 294418 319832 294474 319841
rect 294418 319767 294474 319776
rect 294432 319054 294460 319767
rect 294524 319161 294552 319874
rect 294604 319524 294656 319530
rect 294604 319466 294656 319472
rect 294510 319152 294566 319161
rect 294510 319087 294566 319096
rect 294420 319048 294472 319054
rect 294420 318990 294472 318996
rect 294524 318900 294552 319087
rect 294432 318872 294552 318900
rect 294432 316878 294460 318872
rect 294512 317960 294564 317966
rect 294512 317902 294564 317908
rect 294420 316872 294472 316878
rect 294420 316814 294472 316820
rect 294328 316396 294380 316402
rect 294328 316338 294380 316344
rect 294328 316056 294380 316062
rect 294328 315998 294380 316004
rect 294418 316024 294474 316033
rect 294236 315852 294288 315858
rect 294236 315794 294288 315800
rect 294144 315444 294196 315450
rect 294144 315386 294196 315392
rect 294248 306374 294276 315794
rect 294340 310146 294368 315998
rect 294418 315959 294474 315968
rect 294432 315790 294460 315959
rect 294420 315784 294472 315790
rect 294420 315726 294472 315732
rect 294328 310140 294380 310146
rect 294328 310082 294380 310088
rect 294248 306346 294460 306374
rect 294432 305998 294460 306346
rect 294420 305992 294472 305998
rect 294420 305934 294472 305940
rect 294052 304904 294104 304910
rect 294052 304846 294104 304852
rect 293960 301844 294012 301850
rect 293960 301786 294012 301792
rect 293972 298897 294000 301786
rect 293958 298888 294014 298897
rect 293958 298823 294014 298832
rect 293868 239420 293920 239426
rect 293868 239362 293920 239368
rect 293408 232756 293460 232762
rect 293408 232698 293460 232704
rect 294432 228818 294460 305934
rect 294524 301850 294552 317902
rect 294616 312798 294644 319466
rect 294708 316690 294736 319892
rect 294788 319864 294840 319870
rect 294788 319806 294840 319812
rect 294800 319054 294828 319806
rect 294938 319784 294966 320076
rect 295030 319938 295058 320076
rect 295018 319932 295070 319938
rect 295018 319874 295070 319880
rect 295122 319818 295150 320076
rect 295076 319790 295150 319818
rect 294938 319756 295012 319784
rect 294984 319530 295012 319756
rect 294972 319524 295024 319530
rect 294972 319466 295024 319472
rect 294788 319048 294840 319054
rect 294788 318990 294840 318996
rect 295076 317966 295104 319790
rect 295214 319682 295242 320076
rect 295168 319654 295242 319682
rect 295064 317960 295116 317966
rect 295064 317902 295116 317908
rect 295064 317620 295116 317626
rect 295064 317562 295116 317568
rect 294708 316662 294828 316690
rect 294694 315752 294750 315761
rect 294694 315687 294750 315696
rect 294708 315489 294736 315687
rect 294694 315480 294750 315489
rect 294694 315415 294750 315424
rect 294604 312792 294656 312798
rect 294604 312734 294656 312740
rect 294696 311636 294748 311642
rect 294696 311578 294748 311584
rect 294512 301844 294564 301850
rect 294512 301786 294564 301792
rect 294602 236600 294658 236609
rect 294602 236535 294658 236544
rect 294420 228812 294472 228818
rect 294420 228754 294472 228760
rect 293314 218648 293370 218657
rect 293314 218583 293370 218592
rect 294616 146266 294644 236535
rect 294708 224534 294736 311578
rect 294800 306134 294828 316662
rect 294880 316396 294932 316402
rect 294880 316338 294932 316344
rect 294788 306128 294840 306134
rect 294788 306070 294840 306076
rect 294800 305726 294828 306070
rect 294788 305720 294840 305726
rect 294788 305662 294840 305668
rect 294892 304502 294920 316338
rect 294972 310140 295024 310146
rect 294972 310082 295024 310088
rect 294880 304496 294932 304502
rect 294880 304438 294932 304444
rect 294788 304360 294840 304366
rect 294788 304302 294840 304308
rect 294800 230081 294828 304302
rect 294984 235006 295012 310082
rect 295076 306066 295104 317562
rect 295168 316062 295196 319654
rect 295306 319580 295334 320076
rect 295398 319784 295426 320076
rect 295490 319943 295518 320076
rect 295476 319934 295532 319943
rect 295476 319869 295532 319878
rect 295582 319784 295610 320076
rect 295398 319756 295472 319784
rect 295260 319552 295334 319580
rect 295156 316056 295208 316062
rect 295156 315998 295208 316004
rect 295260 315858 295288 319552
rect 295340 317416 295392 317422
rect 295340 317358 295392 317364
rect 295248 315852 295300 315858
rect 295248 315794 295300 315800
rect 295352 315738 295380 317358
rect 295260 315710 295380 315738
rect 295156 315444 295208 315450
rect 295156 315386 295208 315392
rect 295064 306060 295116 306066
rect 295064 306002 295116 306008
rect 295076 305930 295104 306002
rect 295064 305924 295116 305930
rect 295064 305866 295116 305872
rect 295168 299441 295196 315386
rect 295154 299432 295210 299441
rect 295154 299367 295210 299376
rect 295168 296714 295196 299367
rect 295076 296686 295196 296714
rect 294972 235000 295024 235006
rect 294972 234942 295024 234948
rect 294786 230072 294842 230081
rect 294786 230007 294842 230016
rect 295076 227225 295104 296686
rect 295260 238814 295288 315710
rect 295444 311894 295472 319756
rect 295536 319756 295610 319784
rect 295674 319784 295702 320076
rect 295766 319938 295794 320076
rect 295754 319932 295806 319938
rect 295754 319874 295806 319880
rect 295858 319784 295886 320076
rect 296042 319920 296070 320076
rect 296304 320104 296360 320113
rect 296120 320039 296176 320048
rect 296226 319954 296254 320076
rect 297224 320104 297280 320113
rect 296304 320039 296360 320048
rect 296226 319926 296300 319954
rect 295674 319756 295748 319784
rect 295536 317150 295564 319756
rect 295614 319696 295670 319705
rect 295614 319631 295670 319640
rect 295628 317218 295656 319631
rect 295616 317212 295668 317218
rect 295616 317154 295668 317160
rect 295524 317144 295576 317150
rect 295524 317086 295576 317092
rect 295536 316810 295564 317086
rect 295524 316804 295576 316810
rect 295524 316746 295576 316752
rect 295616 316396 295668 316402
rect 295616 316338 295668 316344
rect 295444 311866 295564 311894
rect 295536 304638 295564 311866
rect 295628 306202 295656 316338
rect 295720 316010 295748 319756
rect 295812 319756 295886 319784
rect 295950 319892 296070 319920
rect 295812 316402 295840 319756
rect 295950 319716 295978 319892
rect 296166 319832 296222 319841
rect 296272 319818 296300 319926
rect 296410 319852 296438 320076
rect 296410 319824 296484 319852
rect 296222 319790 296300 319818
rect 296166 319767 296222 319776
rect 295950 319688 296116 319716
rect 295892 319524 295944 319530
rect 295892 319466 295944 319472
rect 295904 318442 295932 319466
rect 295984 318912 296036 318918
rect 295984 318854 296036 318860
rect 295996 318782 296024 318854
rect 295984 318776 296036 318782
rect 295984 318718 296036 318724
rect 295892 318436 295944 318442
rect 295892 318378 295944 318384
rect 295984 316736 296036 316742
rect 295984 316678 296036 316684
rect 295800 316396 295852 316402
rect 295800 316338 295852 316344
rect 295720 315982 295932 316010
rect 295708 315852 295760 315858
rect 295708 315794 295760 315800
rect 295720 311234 295748 315794
rect 295708 311228 295760 311234
rect 295708 311170 295760 311176
rect 295616 306196 295668 306202
rect 295616 306138 295668 306144
rect 295628 305046 295656 306138
rect 295616 305040 295668 305046
rect 295616 304982 295668 304988
rect 295340 304632 295392 304638
rect 295340 304574 295392 304580
rect 295524 304632 295576 304638
rect 295524 304574 295576 304580
rect 295352 304473 295380 304574
rect 295338 304464 295394 304473
rect 295338 304399 295394 304408
rect 295904 301782 295932 315982
rect 295996 314090 296024 316678
rect 295984 314084 296036 314090
rect 295984 314026 296036 314032
rect 295984 311228 296036 311234
rect 295984 311170 296036 311176
rect 295340 301776 295392 301782
rect 295340 301718 295392 301724
rect 295892 301776 295944 301782
rect 295892 301718 295944 301724
rect 295352 301481 295380 301718
rect 295338 301472 295394 301481
rect 295338 301407 295394 301416
rect 295248 238808 295300 238814
rect 295248 238750 295300 238756
rect 295260 238474 295288 238750
rect 295248 238468 295300 238474
rect 295248 238410 295300 238416
rect 295340 236768 295392 236774
rect 295340 236710 295392 236716
rect 295352 235929 295380 236710
rect 295338 235920 295394 235929
rect 295338 235855 295394 235864
rect 295996 233102 296024 311170
rect 296088 310214 296116 319688
rect 296166 319696 296222 319705
rect 296456 319648 296484 319824
rect 296594 319784 296622 320076
rect 296166 319631 296222 319640
rect 296180 319530 296208 319631
rect 296364 319620 296484 319648
rect 296548 319756 296622 319784
rect 296168 319524 296220 319530
rect 296168 319466 296220 319472
rect 296364 319002 296392 319620
rect 296180 318974 296392 319002
rect 296076 310208 296128 310214
rect 296076 310150 296128 310156
rect 296076 309188 296128 309194
rect 296076 309130 296128 309136
rect 295984 233096 296036 233102
rect 295984 233038 296036 233044
rect 296088 231538 296116 309130
rect 296180 307834 296208 318974
rect 296444 318776 296496 318782
rect 296444 318718 296496 318724
rect 296456 318442 296484 318718
rect 296444 318436 296496 318442
rect 296444 318378 296496 318384
rect 296352 317212 296404 317218
rect 296352 317154 296404 317160
rect 296258 313984 296314 313993
rect 296258 313919 296314 313928
rect 296168 307828 296220 307834
rect 296168 307770 296220 307776
rect 296180 305794 296208 307770
rect 296168 305788 296220 305794
rect 296168 305730 296220 305736
rect 296168 302116 296220 302122
rect 296168 302058 296220 302064
rect 296076 231532 296128 231538
rect 296076 231474 296128 231480
rect 295062 227216 295118 227225
rect 295062 227151 295118 227160
rect 296180 224602 296208 302058
rect 296272 238542 296300 313919
rect 296364 311894 296392 317154
rect 296456 314226 296484 318378
rect 296548 315858 296576 319756
rect 296686 319716 296714 320076
rect 296778 319784 296806 320076
rect 296870 319938 296898 320076
rect 296858 319932 296910 319938
rect 296858 319874 296910 319880
rect 296962 319784 296990 320076
rect 297146 319954 297174 320076
rect 297592 320104 297648 320113
rect 297224 320039 297280 320048
rect 297146 319926 297220 319954
rect 297192 319920 297220 319926
rect 297192 319892 297266 319920
rect 297088 319864 297140 319870
rect 297238 319818 297266 319892
rect 297088 319806 297140 319812
rect 296778 319756 296852 319784
rect 296962 319756 297036 319784
rect 296640 319688 296714 319716
rect 296640 317626 296668 319688
rect 296628 317620 296680 317626
rect 296628 317562 296680 317568
rect 296720 317620 296772 317626
rect 296720 317562 296772 317568
rect 296732 317506 296760 317562
rect 296640 317478 296760 317506
rect 296536 315852 296588 315858
rect 296536 315794 296588 315800
rect 296444 314220 296496 314226
rect 296444 314162 296496 314168
rect 296364 311866 296484 311894
rect 296350 304600 296406 304609
rect 296350 304535 296406 304544
rect 296260 238536 296312 238542
rect 296260 238478 296312 238484
rect 296364 232966 296392 304535
rect 296456 304434 296484 311866
rect 296444 304428 296496 304434
rect 296444 304370 296496 304376
rect 296640 302122 296668 317478
rect 296824 315722 296852 319756
rect 296904 319660 296956 319666
rect 296904 319602 296956 319608
rect 296916 319530 296944 319602
rect 296904 319524 296956 319530
rect 296904 319466 296956 319472
rect 297008 317218 297036 319756
rect 297100 319297 297128 319806
rect 297192 319790 297266 319818
rect 297086 319288 297142 319297
rect 297086 319223 297142 319232
rect 297086 318608 297142 318617
rect 297086 318543 297142 318552
rect 297100 317529 297128 318543
rect 297192 318442 297220 319790
rect 297514 319784 297542 320076
rect 298052 320104 298108 320113
rect 297592 320039 297648 320048
rect 297698 319784 297726 320076
rect 297376 319756 297542 319784
rect 297652 319756 297726 319784
rect 297790 319784 297818 320076
rect 297974 319920 298002 320076
rect 299248 320104 299304 320113
rect 298052 320039 298108 320048
rect 298250 319920 298278 320076
rect 297928 319892 298002 319920
rect 298204 319892 298278 319920
rect 297790 319756 297864 319784
rect 297270 319696 297326 319705
rect 297270 319631 297326 319640
rect 297284 318782 297312 319631
rect 297272 318776 297324 318782
rect 297272 318718 297324 318724
rect 297180 318436 297232 318442
rect 297180 318378 297232 318384
rect 297178 318336 297234 318345
rect 297178 318271 297234 318280
rect 297192 317665 297220 318271
rect 297272 318164 297324 318170
rect 297272 318106 297324 318112
rect 297284 317694 297312 318106
rect 297272 317688 297324 317694
rect 297178 317656 297234 317665
rect 297272 317630 297324 317636
rect 297178 317591 297234 317600
rect 297086 317520 297142 317529
rect 297086 317455 297142 317464
rect 297272 317348 297324 317354
rect 297272 317290 297324 317296
rect 296996 317212 297048 317218
rect 296996 317154 297048 317160
rect 296902 316704 296958 316713
rect 297008 316674 297036 317154
rect 297284 316878 297312 317290
rect 297272 316872 297324 316878
rect 297272 316814 297324 316820
rect 296902 316639 296958 316648
rect 296996 316668 297048 316674
rect 296812 315716 296864 315722
rect 296812 315658 296864 315664
rect 296720 311024 296772 311030
rect 296720 310966 296772 310972
rect 296732 310350 296760 310966
rect 296720 310344 296772 310350
rect 296720 310286 296772 310292
rect 296916 305930 296944 316639
rect 296996 316610 297048 316616
rect 297376 316146 297404 319756
rect 297456 318776 297508 318782
rect 297456 318718 297508 318724
rect 297008 316118 297404 316146
rect 297008 308582 297036 316118
rect 297272 316056 297324 316062
rect 297272 315998 297324 316004
rect 297284 311710 297312 315998
rect 297364 315852 297416 315858
rect 297364 315794 297416 315800
rect 297272 311704 297324 311710
rect 297272 311646 297324 311652
rect 296996 308576 297048 308582
rect 296996 308518 297048 308524
rect 297284 308530 297312 311646
rect 297376 311438 297404 315794
rect 297364 311432 297416 311438
rect 297364 311374 297416 311380
rect 297376 310842 297404 311374
rect 297468 311030 297496 318718
rect 297652 316062 297680 319756
rect 297732 318504 297784 318510
rect 297732 318446 297784 318452
rect 297744 318306 297772 318446
rect 297732 318300 297784 318306
rect 297732 318242 297784 318248
rect 297730 317520 297786 317529
rect 297730 317455 297786 317464
rect 297640 316056 297692 316062
rect 297640 315998 297692 316004
rect 297456 311024 297508 311030
rect 297456 310966 297508 310972
rect 297376 310814 297680 310842
rect 297008 308310 297036 308518
rect 297284 308502 297588 308530
rect 296996 308304 297048 308310
rect 296996 308246 297048 308252
rect 297456 308304 297508 308310
rect 297456 308246 297508 308252
rect 296904 305924 296956 305930
rect 296904 305866 296956 305872
rect 297364 305040 297416 305046
rect 297364 304982 297416 304988
rect 296628 302116 296680 302122
rect 296628 302058 296680 302064
rect 296626 235920 296682 235929
rect 296626 235855 296682 235864
rect 296352 232960 296404 232966
rect 296352 232902 296404 232908
rect 296168 224596 296220 224602
rect 296168 224538 296220 224544
rect 294696 224528 294748 224534
rect 294696 224470 294748 224476
rect 296640 153338 296668 235855
rect 296720 225752 296772 225758
rect 296720 225694 296772 225700
rect 296628 153332 296680 153338
rect 296628 153274 296680 153280
rect 295984 151156 296036 151162
rect 295984 151098 296036 151104
rect 293960 146260 294012 146266
rect 293960 146202 294012 146208
rect 294604 146260 294656 146266
rect 294604 146202 294656 146208
rect 293972 145586 294000 146202
rect 293960 145580 294012 145586
rect 293960 145522 294012 145528
rect 293224 132388 293276 132394
rect 293224 132330 293276 132336
rect 293236 131782 293264 132330
rect 293224 131776 293276 131782
rect 293224 131718 293276 131724
rect 292580 3936 292632 3942
rect 292580 3878 292632 3884
rect 291844 2916 291896 2922
rect 291844 2858 291896 2864
rect 292592 480 292620 3878
rect 295996 3602 296024 151098
rect 296640 147626 296668 153274
rect 296628 147620 296680 147626
rect 296628 147562 296680 147568
rect 296732 16574 296760 225694
rect 297376 224670 297404 304982
rect 297468 228478 297496 308246
rect 297560 239018 297588 308502
rect 297652 239086 297680 310814
rect 297744 307086 297772 317455
rect 297732 307080 297784 307086
rect 297732 307022 297784 307028
rect 297836 306338 297864 319756
rect 297928 315858 297956 319892
rect 298006 319832 298062 319841
rect 298204 319784 298232 319892
rect 298342 319818 298370 320076
rect 298526 319954 298554 320076
rect 298006 319767 298062 319776
rect 297916 315852 297968 315858
rect 297916 315794 297968 315800
rect 297916 315716 297968 315722
rect 297916 315658 297968 315664
rect 297824 306332 297876 306338
rect 297824 306274 297876 306280
rect 297836 305046 297864 306274
rect 297824 305040 297876 305046
rect 297824 304982 297876 304988
rect 297822 304192 297878 304201
rect 297822 304127 297878 304136
rect 297732 295452 297784 295458
rect 297732 295394 297784 295400
rect 297640 239080 297692 239086
rect 297640 239022 297692 239028
rect 297548 239012 297600 239018
rect 297548 238954 297600 238960
rect 297456 228472 297508 228478
rect 297456 228414 297508 228420
rect 297744 225758 297772 295394
rect 297836 239630 297864 304127
rect 297928 301646 297956 315658
rect 298020 309806 298048 319767
rect 298112 319756 298232 319784
rect 298296 319790 298370 319818
rect 298480 319926 298554 319954
rect 298112 319530 298140 319756
rect 298190 319696 298246 319705
rect 298190 319631 298246 319640
rect 298100 319524 298152 319530
rect 298100 319466 298152 319472
rect 298100 318640 298152 318646
rect 298100 318582 298152 318588
rect 298112 317830 298140 318582
rect 298204 317937 298232 319631
rect 298190 317928 298246 317937
rect 298190 317863 298246 317872
rect 298100 317824 298152 317830
rect 298100 317766 298152 317772
rect 298296 317626 298324 319790
rect 298374 319288 298430 319297
rect 298374 319223 298430 319232
rect 298284 317620 298336 317626
rect 298284 317562 298336 317568
rect 298192 315852 298244 315858
rect 298192 315794 298244 315800
rect 298098 314256 298154 314265
rect 298098 314191 298154 314200
rect 298112 313410 298140 314191
rect 298100 313404 298152 313410
rect 298100 313346 298152 313352
rect 298100 312860 298152 312866
rect 298100 312802 298152 312808
rect 298008 309800 298060 309806
rect 298008 309742 298060 309748
rect 298112 308553 298140 312802
rect 298098 308544 298154 308553
rect 298098 308479 298154 308488
rect 298204 302938 298232 315794
rect 298284 315784 298336 315790
rect 298284 315726 298336 315732
rect 298296 303210 298324 315726
rect 298388 307766 298416 319223
rect 298480 318794 298508 319926
rect 298560 319864 298612 319870
rect 298710 319818 298738 320076
rect 298802 319938 298830 320076
rect 298894 319943 298922 320076
rect 298790 319932 298842 319938
rect 298790 319874 298842 319880
rect 298880 319934 298936 319943
rect 298880 319869 298936 319878
rect 298986 319852 299014 320076
rect 299170 319920 299198 320076
rect 299616 320104 299672 320113
rect 299248 320039 299304 320048
rect 299354 319920 299382 320076
rect 299124 319892 299198 319920
rect 299308 319892 299382 319920
rect 298986 319824 299060 319852
rect 298560 319806 298612 319812
rect 298572 319054 298600 319806
rect 298664 319790 298738 319818
rect 298560 319048 298612 319054
rect 298560 318990 298612 318996
rect 298480 318766 298600 318794
rect 298572 310486 298600 318766
rect 298664 312866 298692 319790
rect 298742 319696 298798 319705
rect 298742 319631 298798 319640
rect 298652 312860 298704 312866
rect 298652 312802 298704 312808
rect 298756 311894 298784 319631
rect 298664 311866 298784 311894
rect 298664 311386 298692 311866
rect 298928 311568 298980 311574
rect 298928 311510 298980 311516
rect 298940 311386 298968 311510
rect 298664 311358 298968 311386
rect 298560 310480 298612 310486
rect 298560 310422 298612 310428
rect 298836 310276 298888 310282
rect 298836 310218 298888 310224
rect 298848 310078 298876 310218
rect 298836 310072 298888 310078
rect 298836 310014 298888 310020
rect 298744 309664 298796 309670
rect 298744 309606 298796 309612
rect 298376 307760 298428 307766
rect 298376 307702 298428 307708
rect 298284 303204 298336 303210
rect 298284 303146 298336 303152
rect 298192 302932 298244 302938
rect 298192 302874 298244 302880
rect 297916 301640 297968 301646
rect 297916 301582 297968 301588
rect 297928 293185 297956 301582
rect 298296 296714 298324 303146
rect 298296 296686 298692 296714
rect 297914 293176 297970 293185
rect 297914 293111 297970 293120
rect 297824 239624 297876 239630
rect 297824 239566 297876 239572
rect 298190 236736 298246 236745
rect 298190 236671 298246 236680
rect 297732 225752 297784 225758
rect 297732 225694 297784 225700
rect 297364 224664 297416 224670
rect 297364 224606 297416 224612
rect 298100 168428 298152 168434
rect 298100 168370 298152 168376
rect 296732 16546 297312 16574
rect 294880 3596 294932 3602
rect 294880 3538 294932 3544
rect 295984 3596 296036 3602
rect 295984 3538 296036 3544
rect 293684 2916 293736 2922
rect 293684 2858 293736 2864
rect 293696 480 293724 2858
rect 294892 480 294920 3538
rect 296076 3052 296128 3058
rect 296076 2994 296128 3000
rect 296088 480 296116 2994
rect 297284 480 297312 16546
rect 287766 354 287878 480
rect 287348 326 287878 354
rect 287766 -960 287878 326
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298112 354 298140 168370
rect 298204 150385 298232 236671
rect 298664 230926 298692 296686
rect 298652 230920 298704 230926
rect 298652 230862 298704 230868
rect 298756 229090 298784 309606
rect 298834 308680 298890 308689
rect 298834 308615 298890 308624
rect 298848 230178 298876 308615
rect 298940 233646 298968 311358
rect 299032 302161 299060 319824
rect 299124 315858 299152 319892
rect 299308 319818 299336 319892
rect 299446 319852 299474 320076
rect 299216 319790 299336 319818
rect 299400 319824 299474 319852
rect 299216 316334 299244 319790
rect 299294 319696 299350 319705
rect 299294 319631 299350 319640
rect 299308 318170 299336 319631
rect 299296 318164 299348 318170
rect 299296 318106 299348 318112
rect 299294 318064 299350 318073
rect 299294 317999 299350 318008
rect 299204 316328 299256 316334
rect 299204 316270 299256 316276
rect 299112 315852 299164 315858
rect 299112 315794 299164 315800
rect 299216 314566 299244 316270
rect 299204 314560 299256 314566
rect 299204 314502 299256 314508
rect 299112 310480 299164 310486
rect 299112 310422 299164 310428
rect 299124 310214 299152 310422
rect 299112 310208 299164 310214
rect 299112 310150 299164 310156
rect 299018 302152 299074 302161
rect 299018 302087 299074 302096
rect 299124 239834 299152 310150
rect 299204 307760 299256 307766
rect 299204 307702 299256 307708
rect 299216 307494 299244 307702
rect 299204 307488 299256 307494
rect 299204 307430 299256 307436
rect 299216 240786 299244 307430
rect 299308 293457 299336 317999
rect 299400 315790 299428 319824
rect 299538 319784 299566 320076
rect 300720 320104 300776 320113
rect 299616 320039 299672 320048
rect 299722 319784 299750 320076
rect 299492 319756 299566 319784
rect 299676 319756 299750 319784
rect 299814 319784 299842 320076
rect 299998 319852 300026 320076
rect 299952 319824 300026 319852
rect 299814 319756 299888 319784
rect 299388 315784 299440 315790
rect 299388 315726 299440 315732
rect 299388 303408 299440 303414
rect 299388 303350 299440 303356
rect 299400 302938 299428 303350
rect 299388 302932 299440 302938
rect 299388 302874 299440 302880
rect 299492 301578 299520 319756
rect 299570 319696 299626 319705
rect 299570 319631 299626 319640
rect 299584 307766 299612 319631
rect 299572 307760 299624 307766
rect 299572 307702 299624 307708
rect 299676 303074 299704 319756
rect 299756 319660 299808 319666
rect 299756 319602 299808 319608
rect 299664 303068 299716 303074
rect 299664 303010 299716 303016
rect 299676 302258 299704 303010
rect 299768 302870 299796 319602
rect 299860 316062 299888 319756
rect 299848 316056 299900 316062
rect 299848 315998 299900 316004
rect 299952 316010 299980 319824
rect 300090 319784 300118 320076
rect 300182 319938 300210 320076
rect 300170 319932 300222 319938
rect 300170 319874 300222 319880
rect 300274 319818 300302 320076
rect 300228 319790 300302 319818
rect 300228 319784 300256 319790
rect 300044 319756 300118 319784
rect 300182 319756 300256 319784
rect 300044 317529 300072 319756
rect 300182 319682 300210 319756
rect 300366 319716 300394 320076
rect 300320 319688 300394 319716
rect 300182 319654 300256 319682
rect 300030 317520 300086 317529
rect 300030 317455 300086 317464
rect 299952 315982 300164 316010
rect 300032 315852 300084 315858
rect 300032 315794 300084 315800
rect 299940 315784 299992 315790
rect 299940 315726 299992 315732
rect 299846 314528 299902 314537
rect 299846 314463 299902 314472
rect 299860 313342 299888 314463
rect 299848 313336 299900 313342
rect 299848 313278 299900 313284
rect 299846 312624 299902 312633
rect 299846 312559 299902 312568
rect 299860 303142 299888 312559
rect 299952 305046 299980 315726
rect 300044 307154 300072 315794
rect 300136 312526 300164 315982
rect 300228 315790 300256 319654
rect 300320 317937 300348 319688
rect 300458 319648 300486 320076
rect 300550 319870 300578 320076
rect 300538 319864 300590 319870
rect 300538 319806 300590 319812
rect 300642 319784 300670 320076
rect 300904 320104 300960 320113
rect 300720 320039 300776 320048
rect 300826 319954 300854 320076
rect 301732 320104 301788 320113
rect 300904 320039 300960 320048
rect 300826 319926 300900 319954
rect 300768 319864 300820 319870
rect 300768 319806 300820 319812
rect 300642 319756 300716 319784
rect 300412 319620 300486 319648
rect 300306 317928 300362 317937
rect 300306 317863 300362 317872
rect 300412 315858 300440 319620
rect 300492 318164 300544 318170
rect 300492 318106 300544 318112
rect 300400 315852 300452 315858
rect 300400 315794 300452 315800
rect 300216 315784 300268 315790
rect 300216 315726 300268 315732
rect 300124 312520 300176 312526
rect 300124 312462 300176 312468
rect 300136 311894 300164 312462
rect 300136 311866 300256 311894
rect 300228 311642 300256 311866
rect 300216 311636 300268 311642
rect 300216 311578 300268 311584
rect 300504 309670 300532 318106
rect 300584 316056 300636 316062
rect 300584 315998 300636 316004
rect 300492 309664 300544 309670
rect 300492 309606 300544 309612
rect 300400 308712 300452 308718
rect 300400 308654 300452 308660
rect 300308 307284 300360 307290
rect 300308 307226 300360 307232
rect 300032 307148 300084 307154
rect 300032 307090 300084 307096
rect 299940 305040 299992 305046
rect 299940 304982 299992 304988
rect 299848 303136 299900 303142
rect 299848 303078 299900 303084
rect 299756 302864 299808 302870
rect 299756 302806 299808 302812
rect 299664 302252 299716 302258
rect 299664 302194 299716 302200
rect 299480 301572 299532 301578
rect 299480 301514 299532 301520
rect 299768 296714 299796 302806
rect 300216 302252 300268 302258
rect 300216 302194 300268 302200
rect 299768 296686 300164 296714
rect 299294 293448 299350 293457
rect 299294 293383 299350 293392
rect 299204 240780 299256 240786
rect 299204 240722 299256 240728
rect 299112 239828 299164 239834
rect 299112 239770 299164 239776
rect 299020 237448 299072 237454
rect 299020 237390 299072 237396
rect 299032 236745 299060 237390
rect 299018 236736 299074 236745
rect 299018 236671 299074 236680
rect 298928 233640 298980 233646
rect 298928 233582 298980 233588
rect 298836 230172 298888 230178
rect 298836 230114 298888 230120
rect 298744 229084 298796 229090
rect 298744 229026 298796 229032
rect 299572 225820 299624 225826
rect 299572 225762 299624 225768
rect 298190 150376 298246 150385
rect 298190 150311 298246 150320
rect 299386 150376 299442 150385
rect 299386 150311 299442 150320
rect 299400 149705 299428 150311
rect 299386 149696 299442 149705
rect 299386 149631 299442 149640
rect 299584 3602 299612 225762
rect 300136 224913 300164 296686
rect 300228 226234 300256 302194
rect 300320 230353 300348 307226
rect 300412 234462 300440 308654
rect 300492 307760 300544 307766
rect 300492 307702 300544 307708
rect 300504 307222 300532 307702
rect 300492 307216 300544 307222
rect 300492 307158 300544 307164
rect 300504 235074 300532 307158
rect 300596 302297 300624 315998
rect 300582 302288 300638 302297
rect 300582 302223 300638 302232
rect 300596 301986 300624 302223
rect 300688 302054 300716 319756
rect 300780 303278 300808 319806
rect 300872 319666 300900 319926
rect 301010 319852 301038 320076
rect 300964 319824 301038 319852
rect 300860 319660 300912 319666
rect 300860 319602 300912 319608
rect 300964 319598 300992 319824
rect 301102 319784 301130 320076
rect 301056 319756 301130 319784
rect 301194 319784 301222 320076
rect 301286 319943 301314 320076
rect 301272 319934 301328 319943
rect 301272 319869 301328 319878
rect 301378 319818 301406 320076
rect 301332 319802 301406 319818
rect 301320 319796 301406 319802
rect 301194 319756 301268 319784
rect 300952 319592 301004 319598
rect 300952 319534 301004 319540
rect 300860 318708 300912 318714
rect 300860 318650 300912 318656
rect 300872 316266 300900 318650
rect 300860 316260 300912 316266
rect 300860 316202 300912 316208
rect 300872 315042 300900 316202
rect 301056 316146 301084 319756
rect 301136 319660 301188 319666
rect 301136 319602 301188 319608
rect 301148 319054 301176 319602
rect 301136 319048 301188 319054
rect 301136 318990 301188 318996
rect 300964 316118 301084 316146
rect 300860 315036 300912 315042
rect 300860 314978 300912 314984
rect 300964 314022 300992 316118
rect 301044 316056 301096 316062
rect 301044 315998 301096 316004
rect 300952 314016 301004 314022
rect 300952 313958 301004 313964
rect 300952 313880 301004 313886
rect 300952 313822 301004 313828
rect 300858 313576 300914 313585
rect 300858 313511 300860 313520
rect 300912 313511 300914 313520
rect 300860 313482 300912 313488
rect 300860 305652 300912 305658
rect 300860 305594 300912 305600
rect 300872 305046 300900 305594
rect 300860 305040 300912 305046
rect 300860 304982 300912 304988
rect 300768 303272 300820 303278
rect 300768 303214 300820 303220
rect 300676 302048 300728 302054
rect 300676 301990 300728 301996
rect 300584 301980 300636 301986
rect 300584 301922 300636 301928
rect 300688 301753 300716 301990
rect 300674 301744 300730 301753
rect 300674 301679 300730 301688
rect 300584 301572 300636 301578
rect 300584 301514 300636 301520
rect 300596 293321 300624 301514
rect 300582 293312 300638 293321
rect 300582 293247 300638 293256
rect 300584 289604 300636 289610
rect 300584 289546 300636 289552
rect 300492 235068 300544 235074
rect 300492 235010 300544 235016
rect 300400 234456 300452 234462
rect 300400 234398 300452 234404
rect 300306 230344 300362 230353
rect 300306 230279 300362 230288
rect 300216 226228 300268 226234
rect 300216 226170 300268 226176
rect 300596 225826 300624 289546
rect 300584 225820 300636 225826
rect 300584 225762 300636 225768
rect 300122 224904 300178 224913
rect 300122 224839 300178 224848
rect 300872 224058 300900 304982
rect 300964 303346 300992 313822
rect 301056 307766 301084 315998
rect 301136 315852 301188 315858
rect 301136 315794 301188 315800
rect 301044 307760 301096 307766
rect 301044 307702 301096 307708
rect 301148 307290 301176 315794
rect 301240 314401 301268 319756
rect 301372 319790 301406 319796
rect 301320 319738 301372 319744
rect 301470 319716 301498 320076
rect 301562 319938 301590 320076
rect 301550 319932 301602 319938
rect 301550 319874 301602 319880
rect 301654 319818 301682 320076
rect 302192 320104 302248 320113
rect 301732 320039 301788 320048
rect 301654 319790 301728 319818
rect 301318 319696 301374 319705
rect 301318 319631 301374 319640
rect 301424 319688 301498 319716
rect 301226 314392 301282 314401
rect 301226 314327 301282 314336
rect 301332 314106 301360 319631
rect 301424 315874 301452 319688
rect 301504 319592 301556 319598
rect 301700 319580 301728 319790
rect 301838 319784 301866 320076
rect 301504 319534 301556 319540
rect 301608 319552 301728 319580
rect 301792 319756 301866 319784
rect 301930 319784 301958 320076
rect 302114 319954 302142 320076
rect 302836 320104 302892 320113
rect 302192 320039 302248 320048
rect 302068 319926 302142 319954
rect 301930 319756 302004 319784
rect 301516 318510 301544 319534
rect 301504 318504 301556 318510
rect 301504 318446 301556 318452
rect 301502 315888 301558 315897
rect 301424 315846 301502 315874
rect 301502 315823 301558 315832
rect 301410 315616 301466 315625
rect 301410 315551 301466 315560
rect 301240 314078 301360 314106
rect 301240 313449 301268 314078
rect 301320 314016 301372 314022
rect 301320 313958 301372 313964
rect 301226 313440 301282 313449
rect 301226 313375 301282 313384
rect 301332 310078 301360 313958
rect 301320 310072 301372 310078
rect 301320 310014 301372 310020
rect 301424 308446 301452 315551
rect 301516 315217 301544 315823
rect 301502 315208 301558 315217
rect 301502 315143 301558 315152
rect 301608 313886 301636 319552
rect 301688 319048 301740 319054
rect 301688 318990 301740 318996
rect 301700 316266 301728 318990
rect 301688 316260 301740 316266
rect 301688 316202 301740 316208
rect 301792 315858 301820 319756
rect 301870 319696 301926 319705
rect 301870 319631 301926 319640
rect 301780 315852 301832 315858
rect 301780 315794 301832 315800
rect 301778 315752 301834 315761
rect 301778 315687 301834 315696
rect 301686 314256 301742 314265
rect 301686 314191 301742 314200
rect 301596 313880 301648 313886
rect 301596 313822 301648 313828
rect 301412 308440 301464 308446
rect 301412 308382 301464 308388
rect 301596 307760 301648 307766
rect 301596 307702 301648 307708
rect 301504 307556 301556 307562
rect 301504 307498 301556 307504
rect 301136 307284 301188 307290
rect 301136 307226 301188 307232
rect 301148 307086 301176 307226
rect 301136 307080 301188 307086
rect 301136 307022 301188 307028
rect 301134 303512 301190 303521
rect 301134 303447 301190 303456
rect 300952 303340 301004 303346
rect 300952 303282 301004 303288
rect 300964 302938 300992 303282
rect 301148 303006 301176 303447
rect 301136 303000 301188 303006
rect 301134 302968 301136 302977
rect 301188 302968 301190 302977
rect 300952 302932 301004 302938
rect 301134 302903 301190 302912
rect 300952 302874 301004 302880
rect 301516 225962 301544 307498
rect 301608 307290 301636 307702
rect 301596 307284 301648 307290
rect 301596 307226 301648 307232
rect 301608 230382 301636 307226
rect 301700 237454 301728 314191
rect 301792 307698 301820 315687
rect 301884 311894 301912 319631
rect 301976 317529 302004 319756
rect 301962 317520 302018 317529
rect 301962 317455 302018 317464
rect 302068 316062 302096 319926
rect 302148 319864 302200 319870
rect 302298 319818 302326 320076
rect 302390 319938 302418 320076
rect 302378 319932 302430 319938
rect 302378 319874 302430 319880
rect 302482 319870 302510 320076
rect 302574 319943 302602 320076
rect 302560 319934 302616 319943
rect 302148 319806 302200 319812
rect 302160 319161 302188 319806
rect 302252 319802 302326 319818
rect 302470 319864 302522 319870
rect 302560 319869 302616 319878
rect 302470 319806 302522 319812
rect 302240 319796 302326 319802
rect 302292 319790 302326 319796
rect 302666 319784 302694 320076
rect 302758 319920 302786 320076
rect 303940 320104 303996 320113
rect 302836 320039 302892 320048
rect 302758 319892 302832 319920
rect 302240 319738 302292 319744
rect 302620 319756 302694 319784
rect 302620 319716 302648 319756
rect 302436 319688 302648 319716
rect 302804 319716 302832 319892
rect 302942 319784 302970 320076
rect 303034 319938 303062 320076
rect 303022 319932 303074 319938
rect 303022 319874 303074 319880
rect 302942 319756 303016 319784
rect 302698 319696 302754 319705
rect 302240 319660 302292 319666
rect 302240 319602 302292 319608
rect 302146 319152 302202 319161
rect 302146 319087 302202 319096
rect 302252 316878 302280 319602
rect 302332 319592 302384 319598
rect 302332 319534 302384 319540
rect 302344 318209 302372 319534
rect 302436 318714 302464 319688
rect 302804 319688 302924 319716
rect 302698 319631 302754 319640
rect 302608 319592 302660 319598
rect 302608 319534 302660 319540
rect 302516 319048 302568 319054
rect 302516 318990 302568 318996
rect 302424 318708 302476 318714
rect 302424 318650 302476 318656
rect 302330 318200 302386 318209
rect 302330 318135 302386 318144
rect 302240 316872 302292 316878
rect 302240 316814 302292 316820
rect 302148 316260 302200 316266
rect 302148 316202 302200 316208
rect 302424 316260 302476 316266
rect 302424 316202 302476 316208
rect 302056 316056 302108 316062
rect 302056 315998 302108 316004
rect 301884 311866 302004 311894
rect 301780 307692 301832 307698
rect 301780 307634 301832 307640
rect 301780 304700 301832 304706
rect 301780 304642 301832 304648
rect 301688 237448 301740 237454
rect 301688 237390 301740 237396
rect 301792 231674 301820 304642
rect 301976 303482 302004 311866
rect 302160 310010 302188 316202
rect 302240 316056 302292 316062
rect 302240 315998 302292 316004
rect 302148 310004 302200 310010
rect 302148 309946 302200 309952
rect 302252 307426 302280 315998
rect 302436 307562 302464 316202
rect 302528 309126 302556 318990
rect 302620 317966 302648 319534
rect 302712 318753 302740 319631
rect 302792 319592 302844 319598
rect 302792 319534 302844 319540
rect 302698 318744 302754 318753
rect 302698 318679 302754 318688
rect 302700 318504 302752 318510
rect 302700 318446 302752 318452
rect 302608 317960 302660 317966
rect 302608 317902 302660 317908
rect 302608 317824 302660 317830
rect 302608 317766 302660 317772
rect 302516 309120 302568 309126
rect 302516 309062 302568 309068
rect 302620 308514 302648 317766
rect 302608 308508 302660 308514
rect 302608 308450 302660 308456
rect 302424 307556 302476 307562
rect 302424 307498 302476 307504
rect 302240 307420 302292 307426
rect 302240 307362 302292 307368
rect 302252 306950 302280 307362
rect 302240 306944 302292 306950
rect 302240 306886 302292 306892
rect 301964 303476 302016 303482
rect 301964 303418 302016 303424
rect 302240 300416 302292 300422
rect 302240 300358 302292 300364
rect 302252 300257 302280 300358
rect 302238 300248 302294 300257
rect 302238 300183 302294 300192
rect 302620 296714 302648 308450
rect 302712 307193 302740 318446
rect 302698 307184 302754 307193
rect 302698 307119 302754 307128
rect 302804 303482 302832 319534
rect 302896 311506 302924 319688
rect 302988 316062 303016 319756
rect 303126 319682 303154 320076
rect 303218 319938 303246 320076
rect 303206 319932 303258 319938
rect 303206 319874 303258 319880
rect 303310 319784 303338 320076
rect 303494 319954 303522 320076
rect 303080 319654 303154 319682
rect 303264 319756 303338 319784
rect 303448 319926 303522 319954
rect 303080 317937 303108 319654
rect 303160 319592 303212 319598
rect 303160 319534 303212 319540
rect 303172 319054 303200 319534
rect 303160 319048 303212 319054
rect 303160 318990 303212 318996
rect 303160 318028 303212 318034
rect 303160 317970 303212 317976
rect 303066 317928 303122 317937
rect 303066 317863 303122 317872
rect 303066 316704 303122 316713
rect 303066 316639 303122 316648
rect 302976 316056 303028 316062
rect 302976 315998 303028 316004
rect 303080 311894 303108 316639
rect 303172 316198 303200 317970
rect 303264 317529 303292 319756
rect 303342 319696 303398 319705
rect 303342 319631 303344 319640
rect 303396 319631 303398 319640
rect 303344 319602 303396 319608
rect 303448 317830 303476 319926
rect 303586 319818 303614 320076
rect 303678 319870 303706 320076
rect 303540 319790 303614 319818
rect 303666 319864 303718 319870
rect 303666 319806 303718 319812
rect 303436 317824 303488 317830
rect 303436 317766 303488 317772
rect 303436 317620 303488 317626
rect 303436 317562 303488 317568
rect 303250 317520 303306 317529
rect 303250 317455 303306 317464
rect 303252 317348 303304 317354
rect 303252 317290 303304 317296
rect 303264 316441 303292 317290
rect 303344 316872 303396 316878
rect 303344 316814 303396 316820
rect 303356 316538 303384 316814
rect 303344 316532 303396 316538
rect 303344 316474 303396 316480
rect 303250 316432 303306 316441
rect 303250 316367 303306 316376
rect 303160 316192 303212 316198
rect 303160 316134 303212 316140
rect 303344 316192 303396 316198
rect 303344 316134 303396 316140
rect 303356 315654 303384 316134
rect 303344 315648 303396 315654
rect 303344 315590 303396 315596
rect 302988 311866 303108 311894
rect 303448 311894 303476 317562
rect 303540 316266 303568 319790
rect 303620 319728 303672 319734
rect 303770 319716 303798 320076
rect 303862 319784 303890 320076
rect 304216 320104 304272 320113
rect 303940 320039 303996 320048
rect 304046 319938 304074 320076
rect 304034 319932 304086 319938
rect 304034 319874 304086 319880
rect 304138 319852 304166 320076
rect 304584 320104 304640 320113
rect 304216 320039 304272 320048
rect 304322 319938 304350 320076
rect 304414 319938 304442 320076
rect 304310 319932 304362 319938
rect 304310 319874 304362 319880
rect 304402 319932 304454 319938
rect 304402 319874 304454 319880
rect 304506 319870 304534 320076
rect 305872 320104 305928 320113
rect 304584 320039 304640 320048
rect 304494 319864 304546 319870
rect 304138 319824 304212 319852
rect 303862 319756 303936 319784
rect 303770 319688 303844 319716
rect 303620 319670 303672 319676
rect 303528 316260 303580 316266
rect 303528 316202 303580 316208
rect 303632 312730 303660 319670
rect 303712 319048 303764 319054
rect 303712 318990 303764 318996
rect 303724 318850 303752 318990
rect 303712 318844 303764 318850
rect 303712 318786 303764 318792
rect 303712 317824 303764 317830
rect 303712 317766 303764 317772
rect 303724 316130 303752 317766
rect 303816 317082 303844 319688
rect 303804 317076 303856 317082
rect 303804 317018 303856 317024
rect 303712 316124 303764 316130
rect 303712 316066 303764 316072
rect 303804 316124 303856 316130
rect 303804 316066 303856 316072
rect 303724 313002 303752 316066
rect 303712 312996 303764 313002
rect 303712 312938 303764 312944
rect 303620 312724 303672 312730
rect 303620 312666 303672 312672
rect 303448 311866 303568 311894
rect 302884 311500 302936 311506
rect 302884 311442 302936 311448
rect 302792 303476 302844 303482
rect 302792 303418 302844 303424
rect 302804 302258 302832 303418
rect 302792 302252 302844 302258
rect 302792 302194 302844 302200
rect 302620 296686 302924 296714
rect 301780 231668 301832 231674
rect 301780 231610 301832 231616
rect 301596 230376 301648 230382
rect 301596 230318 301648 230324
rect 302896 229498 302924 296686
rect 302988 238406 303016 311866
rect 303068 309120 303120 309126
rect 303068 309062 303120 309068
rect 303540 309074 303568 311866
rect 303632 310418 303660 312666
rect 303620 310412 303672 310418
rect 303620 310354 303672 310360
rect 303080 308650 303108 309062
rect 303540 309046 303660 309074
rect 303068 308644 303120 308650
rect 303068 308586 303120 308592
rect 302976 238400 303028 238406
rect 302976 238342 303028 238348
rect 303080 234530 303108 308586
rect 303632 308446 303660 309046
rect 303620 308440 303672 308446
rect 303620 308382 303672 308388
rect 303528 307624 303580 307630
rect 303528 307566 303580 307572
rect 303540 306406 303568 307566
rect 303528 306400 303580 306406
rect 303528 306342 303580 306348
rect 303160 304836 303212 304842
rect 303160 304778 303212 304784
rect 303172 239193 303200 304778
rect 303436 303612 303488 303618
rect 303436 303554 303488 303560
rect 303448 303521 303476 303554
rect 303434 303512 303490 303521
rect 303434 303447 303490 303456
rect 303540 303249 303568 306342
rect 303526 303240 303582 303249
rect 303526 303175 303582 303184
rect 303252 302252 303304 302258
rect 303252 302194 303304 302200
rect 303264 247858 303292 302194
rect 303526 297664 303582 297673
rect 303526 297599 303528 297608
rect 303580 297599 303582 297608
rect 303528 297570 303580 297576
rect 303252 247852 303304 247858
rect 303252 247794 303304 247800
rect 303158 239184 303214 239193
rect 303158 239119 303214 239128
rect 303068 234524 303120 234530
rect 303068 234466 303120 234472
rect 303632 230314 303660 308382
rect 303816 302802 303844 316066
rect 303908 307358 303936 319756
rect 303988 319728 304040 319734
rect 303988 319670 304040 319676
rect 304000 318646 304028 319670
rect 304078 319560 304134 319569
rect 304078 319495 304134 319504
rect 303988 318640 304040 318646
rect 303988 318582 304040 318588
rect 303988 318504 304040 318510
rect 303988 318446 304040 318452
rect 304000 309058 304028 318446
rect 304092 314158 304120 319495
rect 304184 316010 304212 319824
rect 304690 319852 304718 320076
rect 304494 319806 304546 319812
rect 304644 319824 304718 319852
rect 304262 319696 304318 319705
rect 304262 319631 304318 319640
rect 304538 319696 304594 319705
rect 304538 319631 304594 319640
rect 304276 317937 304304 319631
rect 304356 319592 304408 319598
rect 304356 319534 304408 319540
rect 304262 317928 304318 317937
rect 304262 317863 304318 317872
rect 304368 316130 304396 319534
rect 304448 319524 304500 319530
rect 304448 319466 304500 319472
rect 304460 317529 304488 319466
rect 304552 318073 304580 319631
rect 304644 318510 304672 319824
rect 304782 319784 304810 320076
rect 304874 319870 304902 320076
rect 304862 319864 304914 319870
rect 304862 319806 304914 319812
rect 304736 319756 304810 319784
rect 304632 318504 304684 318510
rect 304632 318446 304684 318452
rect 304632 318164 304684 318170
rect 304632 318106 304684 318112
rect 304538 318064 304594 318073
rect 304538 317999 304594 318008
rect 304446 317520 304502 317529
rect 304446 317455 304502 317464
rect 304356 316124 304408 316130
rect 304356 316066 304408 316072
rect 304184 315982 304580 316010
rect 304172 315920 304224 315926
rect 304172 315862 304224 315868
rect 304080 314152 304132 314158
rect 304080 314094 304132 314100
rect 303988 309052 304040 309058
rect 303988 308994 304040 309000
rect 303896 307352 303948 307358
rect 303896 307294 303948 307300
rect 303804 302796 303856 302802
rect 303804 302738 303856 302744
rect 303712 300620 303764 300626
rect 303712 300562 303764 300568
rect 303724 300150 303752 300562
rect 303712 300144 303764 300150
rect 303712 300086 303764 300092
rect 304184 297945 304212 315862
rect 304448 307828 304500 307834
rect 304448 307770 304500 307776
rect 304264 307760 304316 307766
rect 304264 307702 304316 307708
rect 304276 300286 304304 307702
rect 304356 305856 304408 305862
rect 304356 305798 304408 305804
rect 304264 300280 304316 300286
rect 304264 300222 304316 300228
rect 304170 297936 304226 297945
rect 304170 297871 304226 297880
rect 304184 290873 304212 297871
rect 304170 290864 304226 290873
rect 304170 290799 304226 290808
rect 303620 230308 303672 230314
rect 303620 230250 303672 230256
rect 302884 229492 302936 229498
rect 302884 229434 302936 229440
rect 301504 225956 301556 225962
rect 301504 225898 301556 225904
rect 300860 224052 300912 224058
rect 300860 223994 300912 224000
rect 304276 217462 304304 300222
rect 304368 227390 304396 305798
rect 304460 230246 304488 307770
rect 304552 307630 304580 315982
rect 304540 307624 304592 307630
rect 304540 307566 304592 307572
rect 304540 302796 304592 302802
rect 304540 302738 304592 302744
rect 304552 244934 304580 302738
rect 304644 300626 304672 318106
rect 304736 315926 304764 319756
rect 304816 319660 304868 319666
rect 304966 319648 304994 320076
rect 305058 319784 305086 320076
rect 305150 319943 305178 320076
rect 305136 319934 305192 319943
rect 305136 319869 305192 319878
rect 305242 319784 305270 320076
rect 305334 319938 305362 320076
rect 305322 319932 305374 319938
rect 305322 319874 305374 319880
rect 305426 319818 305454 320076
rect 305058 319756 305132 319784
rect 304816 319602 304868 319608
rect 304920 319620 304994 319648
rect 304828 317626 304856 319602
rect 304920 318170 304948 319620
rect 304998 319560 305054 319569
rect 304998 319495 305054 319504
rect 304908 318164 304960 318170
rect 304908 318106 304960 318112
rect 305012 318034 305040 319495
rect 305000 318028 305052 318034
rect 305000 317970 305052 317976
rect 304816 317620 304868 317626
rect 304816 317562 304868 317568
rect 304908 317620 304960 317626
rect 304908 317562 304960 317568
rect 304920 316305 304948 317562
rect 304906 316296 304962 316305
rect 304906 316231 304962 316240
rect 304724 315920 304776 315926
rect 304724 315862 304776 315868
rect 304920 314634 304948 316231
rect 304908 314628 304960 314634
rect 304908 314570 304960 314576
rect 304998 309904 305054 309913
rect 304998 309839 305054 309848
rect 305012 309738 305040 309839
rect 305000 309732 305052 309738
rect 305000 309674 305052 309680
rect 304632 300620 304684 300626
rect 304632 300562 304684 300568
rect 305104 298042 305132 319756
rect 305196 319756 305270 319784
rect 305380 319790 305454 319818
rect 305518 319818 305546 320076
rect 305702 319852 305730 320076
rect 305656 319824 305730 319852
rect 305518 319790 305592 319818
rect 305196 319297 305224 319756
rect 305182 319288 305238 319297
rect 305182 319223 305238 319232
rect 305380 317830 305408 319790
rect 305460 319728 305512 319734
rect 305460 319670 305512 319676
rect 305368 317824 305420 317830
rect 305368 317766 305420 317772
rect 305276 316260 305328 316266
rect 305276 316202 305328 316208
rect 305184 315852 305236 315858
rect 305184 315794 305236 315800
rect 305196 300150 305224 315794
rect 305288 300354 305316 316202
rect 305472 316146 305500 319670
rect 305564 316266 305592 319790
rect 305552 316260 305604 316266
rect 305552 316202 305604 316208
rect 305656 316146 305684 319824
rect 305794 319784 305822 320076
rect 306332 320104 306388 320113
rect 305872 320039 305928 320048
rect 305978 319852 306006 320076
rect 305380 316118 305500 316146
rect 305564 316118 305684 316146
rect 305748 319756 305822 319784
rect 305932 319824 306006 319852
rect 305380 307154 305408 316118
rect 305460 316056 305512 316062
rect 305460 315998 305512 316004
rect 305472 308854 305500 315998
rect 305460 308848 305512 308854
rect 305460 308790 305512 308796
rect 305564 308718 305592 316118
rect 305748 315858 305776 319756
rect 305828 319660 305880 319666
rect 305828 319602 305880 319608
rect 305736 315852 305788 315858
rect 305736 315794 305788 315800
rect 305840 315738 305868 319602
rect 305932 316062 305960 319824
rect 306070 319784 306098 320076
rect 306024 319756 306098 319784
rect 305920 316056 305972 316062
rect 305920 315998 305972 316004
rect 305656 315710 305868 315738
rect 305656 309738 305684 315710
rect 306024 311894 306052 319756
rect 306162 319648 306190 320076
rect 306254 319870 306282 320076
rect 306976 320104 307032 320113
rect 306332 320039 306388 320048
rect 306438 319954 306466 320076
rect 306392 319926 306466 319954
rect 306242 319864 306294 319870
rect 306242 319806 306294 319812
rect 306162 319620 306328 319648
rect 305840 311866 306052 311894
rect 305644 309732 305696 309738
rect 305644 309674 305696 309680
rect 305552 308712 305604 308718
rect 305552 308654 305604 308660
rect 305840 307766 305868 311866
rect 306104 308848 306156 308854
rect 306104 308790 306156 308796
rect 305828 307760 305880 307766
rect 305828 307702 305880 307708
rect 305368 307148 305420 307154
rect 305368 307090 305420 307096
rect 305380 306374 305408 307090
rect 305380 306346 305776 306374
rect 305644 300688 305696 300694
rect 305644 300630 305696 300636
rect 305276 300348 305328 300354
rect 305276 300290 305328 300296
rect 305552 300348 305604 300354
rect 305552 300290 305604 300296
rect 305184 300144 305236 300150
rect 305184 300086 305236 300092
rect 305092 298036 305144 298042
rect 305092 297978 305144 297984
rect 305460 298036 305512 298042
rect 305460 297978 305512 297984
rect 305472 289785 305500 297978
rect 305564 295458 305592 300290
rect 305552 295452 305604 295458
rect 305552 295394 305604 295400
rect 305458 289776 305514 289785
rect 305458 289711 305514 289720
rect 304540 244928 304592 244934
rect 304540 244870 304592 244876
rect 304448 230240 304500 230246
rect 304448 230182 304500 230188
rect 304356 227384 304408 227390
rect 304356 227326 304408 227332
rect 305656 226098 305684 300630
rect 305748 233034 305776 306346
rect 306010 305688 306066 305697
rect 306010 305623 306066 305632
rect 305826 301472 305882 301481
rect 305826 301407 305882 301416
rect 305736 233028 305788 233034
rect 305736 232970 305788 232976
rect 305644 226092 305696 226098
rect 305644 226034 305696 226040
rect 303620 217456 303672 217462
rect 303620 217398 303672 217404
rect 304264 217456 304316 217462
rect 304264 217398 304316 217404
rect 303632 217326 303660 217398
rect 303620 217320 303672 217326
rect 303620 217262 303672 217268
rect 302884 140208 302936 140214
rect 302884 140150 302936 140156
rect 301504 131912 301556 131918
rect 301504 131854 301556 131860
rect 301516 3874 301544 131854
rect 301962 6080 302018 6089
rect 301962 6015 302018 6024
rect 301504 3868 301556 3874
rect 301504 3810 301556 3816
rect 299480 3596 299532 3602
rect 299480 3538 299532 3544
rect 299572 3596 299624 3602
rect 299572 3538 299624 3544
rect 300768 3596 300820 3602
rect 300768 3538 300820 3544
rect 299492 1850 299520 3538
rect 299492 1822 299704 1850
rect 299676 480 299704 1822
rect 300780 480 300808 3538
rect 301976 480 302004 6015
rect 302896 4146 302924 140150
rect 303632 16574 303660 217262
rect 305000 171148 305052 171154
rect 305000 171090 305052 171096
rect 305012 16574 305040 171090
rect 303632 16546 303936 16574
rect 305012 16546 305592 16574
rect 302884 4140 302936 4146
rect 302884 4082 302936 4088
rect 303160 4072 303212 4078
rect 303160 4014 303212 4020
rect 303172 480 303200 4014
rect 298438 354 298550 480
rect 298112 326 298550 354
rect 298438 -960 298550 326
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 303908 354 303936 16546
rect 305564 480 305592 16546
rect 305656 3738 305684 226034
rect 305840 221785 305868 301407
rect 305920 296744 305972 296750
rect 305920 296686 305972 296692
rect 305932 225690 305960 296686
rect 306024 234326 306052 305623
rect 306116 240922 306144 308790
rect 306196 300144 306248 300150
rect 306196 300086 306248 300092
rect 306208 289610 306236 300086
rect 306300 297702 306328 319620
rect 306392 315518 306420 319926
rect 306530 319818 306558 320076
rect 306484 319790 306558 319818
rect 306622 319818 306650 320076
rect 306806 319938 306834 320076
rect 306794 319932 306846 319938
rect 306794 319874 306846 319880
rect 306746 319832 306802 319841
rect 306622 319790 306696 319818
rect 306484 317626 306512 319790
rect 306564 319728 306616 319734
rect 306564 319670 306616 319676
rect 306472 317620 306524 317626
rect 306472 317562 306524 317568
rect 306472 315784 306524 315790
rect 306472 315726 306524 315732
rect 306380 315512 306432 315518
rect 306380 315454 306432 315460
rect 306288 297696 306340 297702
rect 306288 297638 306340 297644
rect 306196 289604 306248 289610
rect 306196 289546 306248 289552
rect 306104 240916 306156 240922
rect 306104 240858 306156 240864
rect 306012 234320 306064 234326
rect 306012 234262 306064 234268
rect 305920 225684 305972 225690
rect 305920 225626 305972 225632
rect 305826 221776 305882 221785
rect 305826 221711 305882 221720
rect 305932 219434 305960 225626
rect 306484 223038 306512 315726
rect 306576 300762 306604 319670
rect 306668 315926 306696 319790
rect 306746 319767 306802 319776
rect 306898 319784 306926 320076
rect 307528 320104 307584 320113
rect 306976 320039 307032 320048
rect 307082 319954 307110 320076
rect 307036 319926 307110 319954
rect 306760 317529 306788 319767
rect 306898 319756 306972 319784
rect 306840 317824 306892 317830
rect 306840 317766 306892 317772
rect 306746 317520 306802 317529
rect 306852 317490 306880 317766
rect 306746 317455 306802 317464
rect 306840 317484 306892 317490
rect 306840 317426 306892 317432
rect 306748 316056 306800 316062
rect 306748 315998 306800 316004
rect 306656 315920 306708 315926
rect 306656 315862 306708 315868
rect 306760 307834 306788 315998
rect 306840 315988 306892 315994
rect 306840 315930 306892 315936
rect 306852 309058 306880 315930
rect 306840 309052 306892 309058
rect 306840 308994 306892 309000
rect 306748 307828 306800 307834
rect 306748 307770 306800 307776
rect 306564 300756 306616 300762
rect 306564 300698 306616 300704
rect 306944 299946 306972 319756
rect 307036 315994 307064 319926
rect 307174 319852 307202 320076
rect 307128 319824 307202 319852
rect 307024 315988 307076 315994
rect 307024 315930 307076 315936
rect 307024 315852 307076 315858
rect 307024 315794 307076 315800
rect 307036 309194 307064 315794
rect 307024 309188 307076 309194
rect 307024 309130 307076 309136
rect 307024 300756 307076 300762
rect 307024 300698 307076 300704
rect 307036 300014 307064 300698
rect 307128 300558 307156 319824
rect 307266 319784 307294 320076
rect 307220 319756 307294 319784
rect 307358 319784 307386 320076
rect 307450 319938 307478 320076
rect 308632 320104 308688 320113
rect 307528 320039 307584 320048
rect 307542 319938 307570 320039
rect 307438 319932 307490 319938
rect 307438 319874 307490 319880
rect 307530 319932 307582 319938
rect 307530 319874 307582 319880
rect 307634 319784 307662 320076
rect 307358 319756 307432 319784
rect 307220 317937 307248 319756
rect 307404 318050 307432 319756
rect 307588 319756 307662 319784
rect 307484 319728 307536 319734
rect 307484 319670 307536 319676
rect 307496 318345 307524 319670
rect 307482 318336 307538 318345
rect 307482 318271 307538 318280
rect 307312 318022 307432 318050
rect 307206 317928 307262 317937
rect 307206 317863 307262 317872
rect 307312 316062 307340 318022
rect 307392 317960 307444 317966
rect 307392 317902 307444 317908
rect 307404 317626 307432 317902
rect 307392 317620 307444 317626
rect 307392 317562 307444 317568
rect 307300 316056 307352 316062
rect 307300 315998 307352 316004
rect 307588 315858 307616 319756
rect 307726 319716 307754 320076
rect 307818 319784 307846 320076
rect 308094 319784 308122 320076
rect 307818 319756 307984 319784
rect 307680 319688 307754 319716
rect 307680 316010 307708 319688
rect 307852 316192 307904 316198
rect 307852 316134 307904 316140
rect 307680 315982 307800 316010
rect 307668 315920 307720 315926
rect 307668 315862 307720 315868
rect 307576 315852 307628 315858
rect 307576 315794 307628 315800
rect 307574 314664 307630 314673
rect 307574 314599 307630 314608
rect 307484 309188 307536 309194
rect 307484 309130 307536 309136
rect 307208 309052 307260 309058
rect 307208 308994 307260 309000
rect 307220 308922 307248 308994
rect 307496 308990 307524 309130
rect 307484 308984 307536 308990
rect 307484 308926 307536 308932
rect 307208 308916 307260 308922
rect 307208 308858 307260 308864
rect 307116 300552 307168 300558
rect 307116 300494 307168 300500
rect 307024 300008 307076 300014
rect 307024 299950 307076 299956
rect 306932 299940 306984 299946
rect 306932 299882 306984 299888
rect 306944 296750 306972 299882
rect 306932 296744 306984 296750
rect 306932 296686 306984 296692
rect 307036 226030 307064 299950
rect 307116 292120 307168 292126
rect 307116 292062 307168 292068
rect 307128 228449 307156 292062
rect 307220 261526 307248 308858
rect 307484 308304 307536 308310
rect 307484 308246 307536 308252
rect 307496 307834 307524 308246
rect 307484 307828 307536 307834
rect 307484 307770 307536 307776
rect 307588 297770 307616 314599
rect 307680 303346 307708 315862
rect 307772 315790 307800 315982
rect 307760 315784 307812 315790
rect 307760 315726 307812 315732
rect 307864 315602 307892 316134
rect 307772 315574 307892 315602
rect 307772 313206 307800 315574
rect 307760 313200 307812 313206
rect 307758 313168 307760 313177
rect 307812 313168 307814 313177
rect 307758 313103 307814 313112
rect 307668 303340 307720 303346
rect 307668 303282 307720 303288
rect 307680 300694 307708 303282
rect 307758 302016 307814 302025
rect 307758 301951 307814 301960
rect 307668 300688 307720 300694
rect 307668 300630 307720 300636
rect 307668 300552 307720 300558
rect 307668 300494 307720 300500
rect 307576 297764 307628 297770
rect 307576 297706 307628 297712
rect 307588 290465 307616 297706
rect 307574 290456 307630 290465
rect 307574 290391 307630 290400
rect 307208 261520 307260 261526
rect 307208 261462 307260 261468
rect 307680 247858 307708 300494
rect 307772 300218 307800 301951
rect 307760 300212 307812 300218
rect 307760 300154 307812 300160
rect 307668 247852 307720 247858
rect 307668 247794 307720 247800
rect 307114 228440 307170 228449
rect 307114 228375 307170 228384
rect 307024 226024 307076 226030
rect 307024 225966 307076 225972
rect 306472 223032 306524 223038
rect 306472 222974 306524 222980
rect 305748 219406 305960 219434
rect 305644 3732 305696 3738
rect 305644 3674 305696 3680
rect 305748 3602 305776 219406
rect 307036 4146 307064 225966
rect 307116 223032 307168 223038
rect 307116 222974 307168 222980
rect 307128 158030 307156 222974
rect 307116 158024 307168 158030
rect 307116 157966 307168 157972
rect 307116 152652 307168 152658
rect 307116 152594 307168 152600
rect 306748 4140 306800 4146
rect 306748 4082 306800 4088
rect 307024 4140 307076 4146
rect 307024 4082 307076 4088
rect 305736 3596 305788 3602
rect 305736 3538 305788 3544
rect 306760 480 306788 4082
rect 307128 3126 307156 152594
rect 307668 3596 307720 3602
rect 307668 3538 307720 3544
rect 307680 3398 307708 3538
rect 307772 3482 307800 300154
rect 307956 297362 307984 319756
rect 308048 319756 308122 319784
rect 308186 319784 308214 320076
rect 308278 319920 308306 320076
rect 308462 319954 308490 320076
rect 308416 319926 308490 319954
rect 308278 319892 308352 319920
rect 308186 319756 308260 319784
rect 308048 316198 308076 319756
rect 308232 317354 308260 319756
rect 308220 317348 308272 317354
rect 308220 317290 308272 317296
rect 308232 317014 308260 317290
rect 308220 317008 308272 317014
rect 308220 316950 308272 316956
rect 308036 316192 308088 316198
rect 308036 316134 308088 316140
rect 308036 316056 308088 316062
rect 308036 315998 308088 316004
rect 308048 300082 308076 315998
rect 308220 315988 308272 315994
rect 308220 315930 308272 315936
rect 308128 315920 308180 315926
rect 308128 315862 308180 315868
rect 308140 310010 308168 315862
rect 308232 311098 308260 315930
rect 308324 313274 308352 319892
rect 308416 317286 308444 319926
rect 308554 319784 308582 320076
rect 309736 320104 309792 320113
rect 308632 320039 308688 320048
rect 308738 319784 308766 320076
rect 308922 319852 308950 320076
rect 308508 319756 308582 319784
rect 308692 319756 308766 319784
rect 308876 319824 308950 319852
rect 308404 317280 308456 317286
rect 308404 317222 308456 317228
rect 308416 316606 308444 317222
rect 308404 316600 308456 316606
rect 308404 316542 308456 316548
rect 308508 316062 308536 319756
rect 308496 316056 308548 316062
rect 308496 315998 308548 316004
rect 308588 316056 308640 316062
rect 308588 315998 308640 316004
rect 308312 313268 308364 313274
rect 308312 313210 308364 313216
rect 308220 311092 308272 311098
rect 308220 311034 308272 311040
rect 308128 310004 308180 310010
rect 308128 309946 308180 309952
rect 308140 306374 308168 309946
rect 308600 307902 308628 315998
rect 308692 315926 308720 319756
rect 308680 315920 308732 315926
rect 308680 315862 308732 315868
rect 308876 311894 308904 319824
rect 309014 319784 309042 320076
rect 308968 319756 309042 319784
rect 308968 316062 308996 319756
rect 309106 319716 309134 320076
rect 309060 319688 309134 319716
rect 309198 319716 309226 320076
rect 309290 319784 309318 320076
rect 309382 319852 309410 320076
rect 309474 319954 309502 320076
rect 309658 319954 309686 320076
rect 309920 320104 309976 320113
rect 309736 320039 309792 320048
rect 309474 319926 309548 319954
rect 309658 319926 309732 319954
rect 309382 319824 309456 319852
rect 309290 319756 309364 319784
rect 309198 319688 309272 319716
rect 308956 316056 309008 316062
rect 308956 315998 309008 316004
rect 309060 315994 309088 319688
rect 309048 315988 309100 315994
rect 309048 315930 309100 315936
rect 309048 313268 309100 313274
rect 309048 313210 309100 313216
rect 309060 313138 309088 313210
rect 309048 313132 309100 313138
rect 309048 313074 309100 313080
rect 308692 311866 308904 311894
rect 308588 307896 308640 307902
rect 308588 307838 308640 307844
rect 308140 306346 308444 306374
rect 308036 300076 308088 300082
rect 308036 300018 308088 300024
rect 307944 297356 307996 297362
rect 307944 297298 307996 297304
rect 307956 296714 307984 297298
rect 307864 296686 307984 296714
rect 307864 291825 307892 296686
rect 307850 291816 307906 291825
rect 307850 291751 307906 291760
rect 308416 240990 308444 306346
rect 308692 297838 308720 311866
rect 308956 307896 309008 307902
rect 308956 307838 309008 307844
rect 308968 307329 308996 307838
rect 308954 307320 309010 307329
rect 308954 307255 309010 307264
rect 308680 297832 308732 297838
rect 308680 297774 308732 297780
rect 308692 296714 308720 297774
rect 308508 296686 308720 296714
rect 308508 254590 308536 296686
rect 308496 254584 308548 254590
rect 308496 254526 308548 254532
rect 309060 250510 309088 313074
rect 309138 312216 309194 312225
rect 309138 312151 309194 312160
rect 309152 312050 309180 312151
rect 309140 312044 309192 312050
rect 309140 311986 309192 311992
rect 309244 311894 309272 319688
rect 309336 317490 309364 319756
rect 309324 317484 309376 317490
rect 309324 317426 309376 317432
rect 309244 311866 309364 311894
rect 309336 297974 309364 311866
rect 309428 299878 309456 319824
rect 309520 318617 309548 319926
rect 309598 319832 309654 319841
rect 309598 319767 309654 319776
rect 309506 318608 309562 318617
rect 309506 318543 309562 318552
rect 309508 318504 309560 318510
rect 309508 318446 309560 318452
rect 309520 304434 309548 318446
rect 309612 315450 309640 319767
rect 309704 315858 309732 319926
rect 309842 319920 309870 320076
rect 310932 320104 310988 320113
rect 309920 320039 309976 320048
rect 309796 319892 309870 319920
rect 309796 319462 309824 319892
rect 309874 319832 309930 319841
rect 309874 319767 309930 319776
rect 310026 319784 310054 320076
rect 310210 319954 310238 320076
rect 310486 319954 310514 320076
rect 310210 319938 310284 319954
rect 310210 319932 310296 319938
rect 310210 319926 310244 319932
rect 310244 319874 310296 319880
rect 310440 319926 310514 319954
rect 310152 319864 310204 319870
rect 310150 319832 310152 319841
rect 310204 319832 310206 319841
rect 309784 319456 309836 319462
rect 309784 319398 309836 319404
rect 309888 318170 309916 319767
rect 310026 319756 310100 319784
rect 310150 319767 310206 319776
rect 309968 319456 310020 319462
rect 309968 319398 310020 319404
rect 309876 318164 309928 318170
rect 309876 318106 309928 318112
rect 309876 317960 309928 317966
rect 309876 317902 309928 317908
rect 309888 316742 309916 317902
rect 309876 316736 309928 316742
rect 309876 316678 309928 316684
rect 309784 315988 309836 315994
rect 309784 315930 309836 315936
rect 309692 315852 309744 315858
rect 309692 315794 309744 315800
rect 309600 315444 309652 315450
rect 309600 315386 309652 315392
rect 309796 309058 309824 315930
rect 309876 313268 309928 313274
rect 309876 313210 309928 313216
rect 309888 312662 309916 313210
rect 309876 312656 309928 312662
rect 309876 312598 309928 312604
rect 309784 309052 309836 309058
rect 309784 308994 309836 309000
rect 309796 308417 309824 308994
rect 309782 308408 309838 308417
rect 309782 308343 309838 308352
rect 309508 304428 309560 304434
rect 309508 304370 309560 304376
rect 309520 303822 309548 304370
rect 309508 303816 309560 303822
rect 309508 303758 309560 303764
rect 309416 299872 309468 299878
rect 309416 299814 309468 299820
rect 309324 297968 309376 297974
rect 309324 297910 309376 297916
rect 309428 296714 309456 299814
rect 309428 296686 309824 296714
rect 309048 250504 309100 250510
rect 309048 250446 309100 250452
rect 308404 240984 308456 240990
rect 308404 240926 308456 240932
rect 309796 220114 309824 296686
rect 309784 220108 309836 220114
rect 309784 220050 309836 220056
rect 307852 126404 307904 126410
rect 307852 126346 307904 126352
rect 307864 3602 307892 126346
rect 309796 3942 309824 220050
rect 309888 219298 309916 312598
rect 309980 311370 310008 319398
rect 310072 313274 310100 319756
rect 310336 319592 310388 319598
rect 310150 319560 310206 319569
rect 310336 319534 310388 319540
rect 310150 319495 310206 319504
rect 310164 318322 310192 319495
rect 310242 319288 310298 319297
rect 310242 319223 310298 319232
rect 310256 318510 310284 319223
rect 310244 318504 310296 318510
rect 310244 318446 310296 318452
rect 310164 318294 310284 318322
rect 310152 318164 310204 318170
rect 310152 318106 310204 318112
rect 310060 313268 310112 313274
rect 310060 313210 310112 313216
rect 309968 311364 310020 311370
rect 309968 311306 310020 311312
rect 309968 303816 310020 303822
rect 309968 303758 310020 303764
rect 309980 233170 310008 303758
rect 310060 297968 310112 297974
rect 310060 297910 310112 297916
rect 310072 289241 310100 297910
rect 310164 291825 310192 318106
rect 310256 315994 310284 318294
rect 310244 315988 310296 315994
rect 310244 315930 310296 315936
rect 310244 315852 310296 315858
rect 310244 315794 310296 315800
rect 310150 291816 310206 291825
rect 310150 291751 310206 291760
rect 310058 289232 310114 289241
rect 310058 289167 310114 289176
rect 310060 285728 310112 285734
rect 310060 285670 310112 285676
rect 309968 233164 310020 233170
rect 309968 233106 310020 233112
rect 310072 224874 310100 285670
rect 310164 234297 310192 291751
rect 310256 286346 310284 315794
rect 310348 312934 310376 319534
rect 310440 317966 310468 319926
rect 310578 319784 310606 320076
rect 310762 319852 310790 320076
rect 310854 319920 310882 320076
rect 311668 320104 311724 320113
rect 310932 320039 310988 320048
rect 310854 319892 310928 319920
rect 310762 319824 310836 319852
rect 310532 319756 310606 319784
rect 310532 319666 310560 319756
rect 310520 319660 310572 319666
rect 310520 319602 310572 319608
rect 310612 319660 310664 319666
rect 310612 319602 310664 319608
rect 310428 317960 310480 317966
rect 310428 317902 310480 317908
rect 310520 317484 310572 317490
rect 310520 317426 310572 317432
rect 310336 312928 310388 312934
rect 310336 312870 310388 312876
rect 310348 311894 310376 312870
rect 310348 311866 310468 311894
rect 310440 296714 310468 311866
rect 310532 308786 310560 317426
rect 310520 308780 310572 308786
rect 310520 308722 310572 308728
rect 310624 304706 310652 319602
rect 310702 319560 310758 319569
rect 310702 319495 310758 319504
rect 310716 316946 310744 319495
rect 310704 316940 310756 316946
rect 310704 316882 310756 316888
rect 310704 315988 310756 315994
rect 310704 315930 310756 315936
rect 310612 304700 310664 304706
rect 310612 304642 310664 304648
rect 310716 304473 310744 315930
rect 310808 310962 310836 319824
rect 310900 317472 310928 319892
rect 311038 319784 311066 320076
rect 310992 319756 311066 319784
rect 310992 318782 311020 319756
rect 311130 319716 311158 320076
rect 311222 319938 311250 320076
rect 311210 319932 311262 319938
rect 311210 319874 311262 319880
rect 311314 319784 311342 320076
rect 311498 319784 311526 320076
rect 311084 319688 311158 319716
rect 311268 319756 311342 319784
rect 311452 319756 311526 319784
rect 311590 319784 311618 320076
rect 311944 320104 312000 320113
rect 311668 320039 311724 320048
rect 311774 319852 311802 320076
rect 311728 319824 311802 319852
rect 311590 319756 311664 319784
rect 310980 318776 311032 318782
rect 310980 318718 311032 318724
rect 310900 317444 311020 317472
rect 310888 316056 310940 316062
rect 310888 315998 310940 316004
rect 310796 310956 310848 310962
rect 310796 310898 310848 310904
rect 310702 304464 310758 304473
rect 310702 304399 310758 304408
rect 310716 303793 310744 304399
rect 310900 304337 310928 315998
rect 310992 315586 311020 317444
rect 310980 315580 311032 315586
rect 310980 315522 311032 315528
rect 311084 315466 311112 319688
rect 310992 315438 311112 315466
rect 310992 313886 311020 315438
rect 310980 313880 311032 313886
rect 310980 313822 311032 313828
rect 310992 312594 311020 313822
rect 310980 312588 311032 312594
rect 310980 312530 311032 312536
rect 311268 311894 311296 319756
rect 311452 315994 311480 319756
rect 311440 315988 311492 315994
rect 311440 315930 311492 315936
rect 311532 315988 311584 315994
rect 311532 315930 311584 315936
rect 310992 311866 311296 311894
rect 310992 311778 311020 311866
rect 310980 311772 311032 311778
rect 310980 311714 311032 311720
rect 311164 310956 311216 310962
rect 311164 310898 311216 310904
rect 310886 304328 310942 304337
rect 310886 304263 310942 304272
rect 310702 303784 310758 303793
rect 310702 303719 310758 303728
rect 310900 303657 310928 304263
rect 310886 303648 310942 303657
rect 310886 303583 310942 303592
rect 310348 296686 310468 296714
rect 310244 286340 310296 286346
rect 310244 286282 310296 286288
rect 310256 285734 310284 286282
rect 310244 285728 310296 285734
rect 310244 285670 310296 285676
rect 310348 258126 310376 296686
rect 310336 258120 310388 258126
rect 310256 258068 310336 258074
rect 310256 258062 310388 258068
rect 310256 258046 310376 258062
rect 310256 238338 310284 258046
rect 310244 238332 310296 238338
rect 310244 238274 310296 238280
rect 310150 234288 310206 234297
rect 310150 234223 310206 234232
rect 310060 224868 310112 224874
rect 310060 224810 310112 224816
rect 309876 219292 309928 219298
rect 309876 219234 309928 219240
rect 311176 213246 311204 310898
rect 311544 306374 311572 315930
rect 311636 313138 311664 319756
rect 311728 316062 311756 319824
rect 311866 319784 311894 320076
rect 312772 320104 312828 320113
rect 311944 320039 312000 320048
rect 311992 319864 312044 319870
rect 312142 319852 312170 320076
rect 311992 319806 312044 319812
rect 312096 319824 312170 319852
rect 311820 319756 311894 319784
rect 311716 316056 311768 316062
rect 311716 315998 311768 316004
rect 311820 315994 311848 319756
rect 311898 319696 311954 319705
rect 311898 319631 311900 319640
rect 311952 319631 311954 319640
rect 311900 319602 311952 319608
rect 311808 315988 311860 315994
rect 311808 315930 311860 315936
rect 311900 314084 311952 314090
rect 311900 314026 311952 314032
rect 311912 313342 311940 314026
rect 311900 313336 311952 313342
rect 311900 313278 311952 313284
rect 311624 313132 311676 313138
rect 311624 313074 311676 313080
rect 311636 311894 311664 313074
rect 311912 312905 311940 313278
rect 311898 312896 311954 312905
rect 311898 312831 311954 312840
rect 311636 311866 311756 311894
rect 311544 306346 311664 306374
rect 311254 303784 311310 303793
rect 311254 303719 311310 303728
rect 311268 239562 311296 303719
rect 311438 303648 311494 303657
rect 311438 303583 311494 303592
rect 311348 300552 311400 300558
rect 311348 300494 311400 300500
rect 311360 300014 311388 300494
rect 311348 300008 311400 300014
rect 311348 299950 311400 299956
rect 311348 262200 311400 262206
rect 311348 262142 311400 262148
rect 311360 260982 311388 262142
rect 311348 260976 311400 260982
rect 311348 260918 311400 260924
rect 311256 239556 311308 239562
rect 311256 239498 311308 239504
rect 311360 226166 311388 260918
rect 311452 253230 311480 303583
rect 311530 299296 311586 299305
rect 311530 299231 311586 299240
rect 311544 298926 311572 299231
rect 311532 298920 311584 298926
rect 311532 298862 311584 298868
rect 311636 292534 311664 306346
rect 311624 292528 311676 292534
rect 311624 292470 311676 292476
rect 311636 292126 311664 292470
rect 311624 292120 311676 292126
rect 311624 292062 311676 292068
rect 311728 262206 311756 311866
rect 311808 311772 311860 311778
rect 311808 311714 311860 311720
rect 311716 262200 311768 262206
rect 311716 262142 311768 262148
rect 311820 258074 311848 311714
rect 312004 304774 312032 319806
rect 312096 316266 312124 319824
rect 312234 319784 312262 320076
rect 312188 319756 312262 319784
rect 312084 316260 312136 316266
rect 312084 316202 312136 316208
rect 312188 316146 312216 319756
rect 312326 319682 312354 320076
rect 312418 319784 312446 320076
rect 312510 319852 312538 320076
rect 312602 319954 312630 320076
rect 313416 320104 313472 320113
rect 312772 320039 312828 320048
rect 312878 319954 312906 320076
rect 312602 319926 312676 319954
rect 312510 319824 312584 319852
rect 312418 319756 312492 319784
rect 312326 319654 312400 319682
rect 312268 319592 312320 319598
rect 312268 319534 312320 319540
rect 312096 316118 312216 316146
rect 312096 314090 312124 316118
rect 312176 315988 312228 315994
rect 312176 315930 312228 315936
rect 312084 314084 312136 314090
rect 312084 314026 312136 314032
rect 312084 313812 312136 313818
rect 312084 313754 312136 313760
rect 311992 304768 312044 304774
rect 311992 304710 312044 304716
rect 312004 304366 312032 304710
rect 312096 304609 312124 313754
rect 312188 307426 312216 315930
rect 312280 310418 312308 319534
rect 312372 315489 312400 319654
rect 312358 315480 312414 315489
rect 312358 315415 312414 315424
rect 312464 315382 312492 319756
rect 312556 317529 312584 319824
rect 312542 317520 312598 317529
rect 312542 317455 312598 317464
rect 312648 315994 312676 319926
rect 312740 319926 312906 319954
rect 312636 315988 312688 315994
rect 312636 315930 312688 315936
rect 312452 315376 312504 315382
rect 312452 315318 312504 315324
rect 312452 315172 312504 315178
rect 312452 315114 312504 315120
rect 312464 311846 312492 315114
rect 312740 313818 312768 319926
rect 312818 319832 312874 319841
rect 312818 319767 312874 319776
rect 312970 319784 312998 320076
rect 313154 319938 313182 320076
rect 313142 319932 313194 319938
rect 313142 319874 313194 319880
rect 313094 319832 313150 319841
rect 312832 319530 312860 319767
rect 312970 319756 313044 319784
rect 313246 319784 313274 320076
rect 313094 319767 313150 319776
rect 312820 319524 312872 319530
rect 312820 319466 312872 319472
rect 312820 316260 312872 316266
rect 312820 316202 312872 316208
rect 312728 313812 312780 313818
rect 312728 313754 312780 313760
rect 312452 311840 312504 311846
rect 312452 311782 312504 311788
rect 312268 310412 312320 310418
rect 312268 310354 312320 310360
rect 312176 307420 312228 307426
rect 312176 307362 312228 307368
rect 312188 306374 312216 307362
rect 312188 306346 312584 306374
rect 312082 304600 312138 304609
rect 312082 304535 312138 304544
rect 311992 304360 312044 304366
rect 311992 304302 312044 304308
rect 311544 258046 311848 258074
rect 311544 255406 311572 258046
rect 311532 255400 311584 255406
rect 311532 255342 311584 255348
rect 311440 253224 311492 253230
rect 311440 253166 311492 253172
rect 311348 226160 311400 226166
rect 311348 226102 311400 226108
rect 311544 224806 311572 255342
rect 312556 240854 312584 306346
rect 312832 301918 312860 316202
rect 313016 315178 313044 319756
rect 313108 315790 313136 319767
rect 313200 319756 313274 319784
rect 313338 319784 313366 320076
rect 314428 320104 314484 320113
rect 313416 320039 313472 320048
rect 313522 319784 313550 320076
rect 313706 319841 313734 320076
rect 313798 319938 313826 320076
rect 313786 319932 313838 319938
rect 313786 319874 313838 319880
rect 313692 319832 313748 319841
rect 313338 319756 313412 319784
rect 313522 319756 313596 319784
rect 313890 319784 313918 320076
rect 313982 319818 314010 320076
rect 314074 319938 314102 320076
rect 314258 319954 314286 320076
rect 314062 319932 314114 319938
rect 314062 319874 314114 319880
rect 314212 319926 314286 319954
rect 313982 319790 314056 319818
rect 313692 319767 313748 319776
rect 313200 319598 313228 319756
rect 313278 319696 313334 319705
rect 313278 319631 313334 319640
rect 313188 319592 313240 319598
rect 313188 319534 313240 319540
rect 313292 317801 313320 319631
rect 313384 317937 313412 319756
rect 313568 319716 313596 319756
rect 313844 319756 313918 319784
rect 313568 319688 313780 319716
rect 313556 319592 313608 319598
rect 313556 319534 313608 319540
rect 313646 319560 313702 319569
rect 313464 318912 313516 318918
rect 313464 318854 313516 318860
rect 313370 317928 313426 317937
rect 313370 317863 313426 317872
rect 313278 317792 313334 317801
rect 313278 317727 313334 317736
rect 313096 315784 313148 315790
rect 313096 315726 313148 315732
rect 313004 315172 313056 315178
rect 313004 315114 313056 315120
rect 313016 314974 313044 315114
rect 313004 314968 313056 314974
rect 313004 314910 313056 314916
rect 312912 310412 312964 310418
rect 312912 310354 312964 310360
rect 312820 301912 312872 301918
rect 312820 301854 312872 301860
rect 312924 259486 312952 310354
rect 313004 301912 313056 301918
rect 313004 301854 313056 301860
rect 312912 259480 312964 259486
rect 312912 259422 312964 259428
rect 312924 258074 312952 259422
rect 312648 258046 312952 258074
rect 312544 240848 312596 240854
rect 312544 240790 312596 240796
rect 311532 224800 311584 224806
rect 311532 224742 311584 224748
rect 312648 221814 312676 258046
rect 312912 256760 312964 256766
rect 312912 256702 312964 256708
rect 312728 253972 312780 253978
rect 312728 253914 312780 253920
rect 312636 221808 312688 221814
rect 312636 221750 312688 221756
rect 312740 221746 312768 253914
rect 312820 253224 312872 253230
rect 312820 253166 312872 253172
rect 312832 222086 312860 253166
rect 312924 230858 312952 256702
rect 313016 251326 313044 301854
rect 313108 256766 313136 315726
rect 313186 312624 313242 312633
rect 313186 312559 313242 312568
rect 313200 312254 313228 312559
rect 313188 312248 313240 312254
rect 313188 312190 313240 312196
rect 313188 311840 313240 311846
rect 313188 311782 313240 311788
rect 313096 256760 313148 256766
rect 313096 256702 313148 256708
rect 313200 253978 313228 311782
rect 313280 311636 313332 311642
rect 313280 311578 313332 311584
rect 313292 311302 313320 311578
rect 313280 311296 313332 311302
rect 313280 311238 313332 311244
rect 313476 310486 313504 318854
rect 313568 311846 313596 319534
rect 313646 319495 313702 319504
rect 313660 319025 313688 319495
rect 313646 319016 313702 319025
rect 313646 318951 313702 318960
rect 313648 317620 313700 317626
rect 313648 317562 313700 317568
rect 313660 317490 313688 317562
rect 313648 317484 313700 317490
rect 313648 317426 313700 317432
rect 313752 315314 313780 319688
rect 313844 317937 313872 319756
rect 314028 318794 314056 319790
rect 314106 319696 314162 319705
rect 314106 319631 314162 319640
rect 313936 318766 314056 318794
rect 313830 317928 313886 317937
rect 313830 317863 313886 317872
rect 313936 316010 313964 318766
rect 314014 317928 314070 317937
rect 314014 317863 314070 317872
rect 313844 315982 313964 316010
rect 313740 315308 313792 315314
rect 313740 315250 313792 315256
rect 313844 311894 313872 315982
rect 313924 315716 313976 315722
rect 313924 315658 313976 315664
rect 313936 315178 313964 315658
rect 313924 315172 313976 315178
rect 313924 315114 313976 315120
rect 313660 311866 313872 311894
rect 313556 311840 313608 311846
rect 313556 311782 313608 311788
rect 313660 311642 313688 311866
rect 313648 311636 313700 311642
rect 313648 311578 313700 311584
rect 313464 310480 313516 310486
rect 313464 310422 313516 310428
rect 313280 303680 313332 303686
rect 313280 303622 313332 303628
rect 313292 303385 313320 303622
rect 313278 303376 313334 303385
rect 313278 303311 313334 303320
rect 313188 253972 313240 253978
rect 313188 253914 313240 253920
rect 313004 251320 313056 251326
rect 313004 251262 313056 251268
rect 312912 230852 312964 230858
rect 312912 230794 312964 230800
rect 313016 227594 313044 251262
rect 313004 227588 313056 227594
rect 313004 227530 313056 227536
rect 312820 222080 312872 222086
rect 312820 222022 312872 222028
rect 312728 221740 312780 221746
rect 312728 221682 312780 221688
rect 313936 214606 313964 315114
rect 314028 219230 314056 317863
rect 314120 316033 314148 319631
rect 314212 319297 314240 319926
rect 314350 319784 314378 320076
rect 314888 320104 314944 320113
rect 314428 320039 314484 320048
rect 314534 319784 314562 320076
rect 314626 319938 314654 320076
rect 314718 319938 314746 320076
rect 314614 319932 314666 319938
rect 314614 319874 314666 319880
rect 314706 319932 314758 319938
rect 314706 319874 314758 319880
rect 314304 319756 314378 319784
rect 314488 319756 314562 319784
rect 314658 319832 314714 319841
rect 314810 319818 314838 320076
rect 315256 320104 315312 320113
rect 314888 320039 314944 320048
rect 314994 319954 315022 320076
rect 314658 319767 314714 319776
rect 314764 319790 314838 319818
rect 314948 319926 315022 319954
rect 314198 319288 314254 319297
rect 314198 319223 314254 319232
rect 314106 316024 314162 316033
rect 314162 315982 314240 316010
rect 314106 315959 314162 315968
rect 314106 314528 314162 314537
rect 314106 314463 314162 314472
rect 314120 225894 314148 314463
rect 314212 313954 314240 315982
rect 314200 313948 314252 313954
rect 314200 313890 314252 313896
rect 314200 310480 314252 310486
rect 314200 310422 314252 310428
rect 314108 225888 314160 225894
rect 314108 225830 314160 225836
rect 314212 223106 314240 310422
rect 314304 307766 314332 319756
rect 314384 319592 314436 319598
rect 314384 319534 314436 319540
rect 314396 315722 314424 319534
rect 314384 315716 314436 315722
rect 314384 315658 314436 315664
rect 314488 311894 314516 319756
rect 314568 319660 314620 319666
rect 314568 319602 314620 319608
rect 314580 318918 314608 319602
rect 314568 318912 314620 318918
rect 314568 318854 314620 318860
rect 314568 318776 314620 318782
rect 314568 318718 314620 318724
rect 314580 316878 314608 318718
rect 314568 316872 314620 316878
rect 314568 316814 314620 316820
rect 314672 315518 314700 319767
rect 314764 318646 314792 319790
rect 314844 319592 314896 319598
rect 314844 319534 314896 319540
rect 314752 318640 314804 318646
rect 314752 318582 314804 318588
rect 314752 316668 314804 316674
rect 314752 316610 314804 316616
rect 314660 315512 314712 315518
rect 314660 315454 314712 315460
rect 314396 311866 314516 311894
rect 314292 307760 314344 307766
rect 314292 307702 314344 307708
rect 314304 223174 314332 307702
rect 314396 304201 314424 311866
rect 314568 311840 314620 311846
rect 314568 311782 314620 311788
rect 314382 304192 314438 304201
rect 314382 304127 314438 304136
rect 314580 248606 314608 311782
rect 314660 304836 314712 304842
rect 314660 304778 314712 304784
rect 314672 304230 314700 304778
rect 314660 304224 314712 304230
rect 314660 304166 314712 304172
rect 314764 300626 314792 316610
rect 314856 303657 314884 319534
rect 314948 315994 314976 319926
rect 315086 319852 315114 320076
rect 315040 319824 315114 319852
rect 315040 318238 315068 319824
rect 315178 319784 315206 320076
rect 316176 320104 316232 320113
rect 315256 320039 315312 320048
rect 315362 319938 315390 320076
rect 315350 319932 315402 319938
rect 315350 319874 315402 319880
rect 315454 319818 315482 320076
rect 315546 319938 315574 320076
rect 315534 319932 315586 319938
rect 315534 319874 315586 319880
rect 315454 319790 315528 319818
rect 315178 319756 315252 319784
rect 315120 319660 315172 319666
rect 315120 319602 315172 319608
rect 315028 318232 315080 318238
rect 315028 318174 315080 318180
rect 315028 316056 315080 316062
rect 315028 315998 315080 316004
rect 314936 315988 314988 315994
rect 314936 315930 314988 315936
rect 314936 315852 314988 315858
rect 314936 315794 314988 315800
rect 314948 304366 314976 315794
rect 315040 304842 315068 315998
rect 315132 308242 315160 319602
rect 315224 315926 315252 319756
rect 315500 319682 315528 319790
rect 315638 319784 315666 320076
rect 315730 319852 315758 320076
rect 315914 319954 315942 320076
rect 315868 319926 315942 319954
rect 315730 319824 315804 319852
rect 315638 319756 315712 319784
rect 315408 319654 315528 319682
rect 315578 319696 315634 319705
rect 315408 316674 315436 319654
rect 315578 319631 315580 319640
rect 315632 319631 315634 319640
rect 315580 319602 315632 319608
rect 315488 319592 315540 319598
rect 315488 319534 315540 319540
rect 315396 316668 315448 316674
rect 315396 316610 315448 316616
rect 315396 316396 315448 316402
rect 315396 316338 315448 316344
rect 315212 315920 315264 315926
rect 315212 315862 315264 315868
rect 315120 308236 315172 308242
rect 315120 308178 315172 308184
rect 315028 304836 315080 304842
rect 315028 304778 315080 304784
rect 314936 304360 314988 304366
rect 314936 304302 314988 304308
rect 315304 304360 315356 304366
rect 315304 304302 315356 304308
rect 314842 303648 314898 303657
rect 314842 303583 314898 303592
rect 314752 300620 314804 300626
rect 314752 300562 314804 300568
rect 314568 248600 314620 248606
rect 314568 248542 314620 248548
rect 314580 238754 314608 248542
rect 315316 246362 315344 304302
rect 315408 258777 315436 316338
rect 315500 316062 315528 319534
rect 315592 317937 315620 319602
rect 315684 319598 315712 319756
rect 315672 319592 315724 319598
rect 315672 319534 315724 319540
rect 315578 317928 315634 317937
rect 315578 317863 315634 317872
rect 315776 317529 315804 319824
rect 315762 317520 315818 317529
rect 315762 317455 315818 317464
rect 315488 316056 315540 316062
rect 315488 315998 315540 316004
rect 315672 315988 315724 315994
rect 315672 315930 315724 315936
rect 315488 308236 315540 308242
rect 315488 308178 315540 308184
rect 315500 285054 315528 308178
rect 315684 297430 315712 315930
rect 315868 315858 315896 319926
rect 316006 319818 316034 320076
rect 316098 319954 316126 320076
rect 316912 320104 316968 320113
rect 316176 320039 316232 320048
rect 316098 319926 316172 319954
rect 315960 319790 316034 319818
rect 315960 317286 315988 319790
rect 316038 319696 316094 319705
rect 316038 319631 316094 319640
rect 315948 317280 316000 317286
rect 315948 317222 316000 317228
rect 315960 316402 315988 317222
rect 315948 316396 316000 316402
rect 315948 316338 316000 316344
rect 315948 315920 316000 315926
rect 315948 315862 316000 315868
rect 315856 315852 315908 315858
rect 315856 315794 315908 315800
rect 315856 300620 315908 300626
rect 315856 300562 315908 300568
rect 315672 297424 315724 297430
rect 315672 297366 315724 297372
rect 315488 285048 315540 285054
rect 315488 284990 315540 284996
rect 315488 272536 315540 272542
rect 315488 272478 315540 272484
rect 315394 258768 315450 258777
rect 315394 258703 315450 258712
rect 315396 247104 315448 247110
rect 315396 247046 315448 247052
rect 315304 246356 315356 246362
rect 315304 246298 315356 246304
rect 315304 243092 315356 243098
rect 315304 243034 315356 243040
rect 314396 238726 314608 238754
rect 314292 223168 314344 223174
rect 314292 223110 314344 223116
rect 314200 223100 314252 223106
rect 314200 223042 314252 223048
rect 314396 221882 314424 238726
rect 315316 222018 315344 243034
rect 315408 238202 315436 247046
rect 315396 238196 315448 238202
rect 315396 238138 315448 238144
rect 315500 222193 315528 272478
rect 315868 247110 315896 300562
rect 315856 247104 315908 247110
rect 315856 247046 315908 247052
rect 315960 243098 315988 315862
rect 316052 299334 316080 319631
rect 316144 317665 316172 319926
rect 316282 319784 316310 320076
rect 316374 319852 316402 320076
rect 316558 319954 316586 320076
rect 316558 319926 316632 319954
rect 316374 319824 316540 319852
rect 316282 319756 316448 319784
rect 316130 317656 316186 317665
rect 316130 317591 316186 317600
rect 316132 316056 316184 316062
rect 316132 315998 316184 316004
rect 316144 299470 316172 315998
rect 316224 315988 316276 315994
rect 316224 315930 316276 315936
rect 316236 305862 316264 315930
rect 316420 315450 316448 319756
rect 316512 316062 316540 319824
rect 316500 316056 316552 316062
rect 316500 315998 316552 316004
rect 316408 315444 316460 315450
rect 316408 315386 316460 315392
rect 316604 311817 316632 319926
rect 316742 319784 316770 320076
rect 316834 319852 316862 320076
rect 318292 320104 318348 320113
rect 316912 320039 316968 320048
rect 316834 319824 316908 319852
rect 316742 319756 316816 319784
rect 316684 317348 316736 317354
rect 316684 317290 316736 317296
rect 316696 317014 316724 317290
rect 316684 317008 316736 317014
rect 316684 316950 316736 316956
rect 316788 315586 316816 319756
rect 316880 318617 316908 319824
rect 317018 319784 317046 320076
rect 317202 319920 317230 320076
rect 317294 319938 317322 320076
rect 317156 319892 317230 319920
rect 317282 319932 317334 319938
rect 317156 319802 317184 319892
rect 317282 319874 317334 319880
rect 317386 319818 317414 320076
rect 316972 319756 317046 319784
rect 317144 319796 317196 319802
rect 316866 318608 316922 318617
rect 316866 318543 316922 318552
rect 316866 318472 316922 318481
rect 316866 318407 316922 318416
rect 316776 315580 316828 315586
rect 316776 315522 316828 315528
rect 316880 314362 316908 318407
rect 316972 315994 317000 319756
rect 317144 319738 317196 319744
rect 317236 319796 317288 319802
rect 317236 319738 317288 319744
rect 317340 319790 317414 319818
rect 317050 319696 317106 319705
rect 317050 319631 317106 319640
rect 317144 319660 317196 319666
rect 317064 317121 317092 319631
rect 317144 319602 317196 319608
rect 317156 318753 317184 319602
rect 317142 318744 317198 318753
rect 317142 318679 317198 318688
rect 317142 318608 317198 318617
rect 317142 318543 317198 318552
rect 317050 317112 317106 317121
rect 317050 317047 317106 317056
rect 317064 317014 317092 317047
rect 317052 317008 317104 317014
rect 317052 316950 317104 316956
rect 316960 315988 317012 315994
rect 316960 315930 317012 315936
rect 316868 314356 316920 314362
rect 316868 314298 316920 314304
rect 316880 311894 316908 314298
rect 317156 313070 317184 318543
rect 317248 317529 317276 319738
rect 317234 317520 317290 317529
rect 317234 317455 317290 317464
rect 317340 313750 317368 319790
rect 317478 319784 317506 320076
rect 317570 319852 317598 320076
rect 317846 319938 317874 320076
rect 317834 319932 317886 319938
rect 317834 319874 317886 319880
rect 317938 319870 317966 320076
rect 317926 319864 317978 319870
rect 317570 319824 317644 319852
rect 317478 319756 317552 319784
rect 317524 319648 317552 319756
rect 317616 319716 317644 319824
rect 317926 319806 317978 319812
rect 318122 319818 318150 320076
rect 318568 320104 318624 320113
rect 318292 320039 318348 320048
rect 318398 319954 318426 320076
rect 318352 319926 318426 319954
rect 317788 319796 317840 319802
rect 318122 319790 318196 319818
rect 317788 319738 317840 319744
rect 317616 319688 317736 319716
rect 317524 319620 317598 319648
rect 317570 319580 317598 319620
rect 317570 319552 317644 319580
rect 317510 319152 317566 319161
rect 317510 319087 317566 319096
rect 317418 319016 317474 319025
rect 317418 318951 317474 318960
rect 317328 313744 317380 313750
rect 317328 313686 317380 313692
rect 317144 313064 317196 313070
rect 317144 313006 317196 313012
rect 316880 311866 317092 311894
rect 316590 311808 316646 311817
rect 316590 311743 316646 311752
rect 316224 305856 316276 305862
rect 316224 305798 316276 305804
rect 316960 305856 317012 305862
rect 316960 305798 317012 305804
rect 316972 305454 317000 305798
rect 316960 305448 317012 305454
rect 316960 305390 317012 305396
rect 316132 299464 316184 299470
rect 316132 299406 316184 299412
rect 316776 299464 316828 299470
rect 316776 299406 316828 299412
rect 316040 299328 316092 299334
rect 316040 299270 316092 299276
rect 316682 299296 316738 299305
rect 316682 299231 316738 299240
rect 316696 251841 316724 299231
rect 316788 264217 316816 299406
rect 316868 299328 316920 299334
rect 316868 299270 316920 299276
rect 316880 267073 316908 299270
rect 316866 267064 316922 267073
rect 316866 266999 316922 267008
rect 316774 264208 316830 264217
rect 316774 264143 316830 264152
rect 317064 258074 317092 311866
rect 316972 258046 317092 258074
rect 316972 255338 317000 258046
rect 316960 255332 317012 255338
rect 316960 255274 317012 255280
rect 316776 251864 316828 251870
rect 316682 251832 316738 251841
rect 316776 251806 316828 251812
rect 316682 251767 316738 251776
rect 316040 248532 316092 248538
rect 316040 248474 316092 248480
rect 316052 247790 316080 248474
rect 316040 247784 316092 247790
rect 316040 247726 316092 247732
rect 316684 245676 316736 245682
rect 316684 245618 316736 245624
rect 315948 243092 316000 243098
rect 315948 243034 316000 243040
rect 316696 223310 316724 245618
rect 316684 223304 316736 223310
rect 316684 223246 316736 223252
rect 315486 222184 315542 222193
rect 315486 222119 315542 222128
rect 315304 222012 315356 222018
rect 315304 221954 315356 221960
rect 316788 221950 316816 251806
rect 316868 244316 316920 244322
rect 316868 244258 316920 244264
rect 316880 223242 316908 244258
rect 316972 238270 317000 255274
rect 317156 248538 317184 313006
rect 317234 311808 317290 311817
rect 317234 311743 317290 311752
rect 317144 248532 317196 248538
rect 317144 248474 317196 248480
rect 317248 245682 317276 311743
rect 317236 245676 317288 245682
rect 317236 245618 317288 245624
rect 317340 244526 317368 313686
rect 317432 299305 317460 318951
rect 317524 318102 317552 319087
rect 317512 318096 317564 318102
rect 317512 318038 317564 318044
rect 317616 316282 317644 319552
rect 317708 318510 317736 319688
rect 317800 318782 317828 319738
rect 317880 319728 317932 319734
rect 317878 319696 317880 319705
rect 317932 319696 317934 319705
rect 318168 319648 318196 319790
rect 318248 319796 318300 319802
rect 318248 319738 318300 319744
rect 317878 319631 317934 319640
rect 317984 319620 318196 319648
rect 317878 319560 317934 319569
rect 317878 319495 317934 319504
rect 317788 318776 317840 318782
rect 317788 318718 317840 318724
rect 317696 318504 317748 318510
rect 317696 318446 317748 318452
rect 317892 316810 317920 319495
rect 317984 318918 318012 319620
rect 318154 319560 318210 319569
rect 318064 319524 318116 319530
rect 318260 319530 318288 319738
rect 318352 319648 318380 319926
rect 318490 319920 318518 320076
rect 319120 320104 319176 320113
rect 318568 320039 318624 320048
rect 318490 319892 318564 319920
rect 318352 319620 318472 319648
rect 318154 319495 318210 319504
rect 318248 319524 318300 319530
rect 318064 319466 318116 319472
rect 317972 318912 318024 318918
rect 317972 318854 318024 318860
rect 318076 317830 318104 319466
rect 318064 317824 318116 317830
rect 318064 317766 318116 317772
rect 317880 316804 317932 316810
rect 317880 316746 317932 316752
rect 317616 316254 318104 316282
rect 317696 316124 317748 316130
rect 317696 316066 317748 316072
rect 317512 316056 317564 316062
rect 317512 315998 317564 316004
rect 317524 310282 317552 315998
rect 317604 315784 317656 315790
rect 317604 315726 317656 315732
rect 317512 310276 317564 310282
rect 317512 310218 317564 310224
rect 317616 304978 317644 315726
rect 317708 306377 317736 316066
rect 317880 315988 317932 315994
rect 317880 315930 317932 315936
rect 317892 311273 317920 315930
rect 318076 314378 318104 316254
rect 318168 314498 318196 319495
rect 318248 319466 318300 319472
rect 318340 319524 318392 319530
rect 318340 319466 318392 319472
rect 318246 319424 318302 319433
rect 318246 319359 318302 319368
rect 318260 316062 318288 319359
rect 318352 319161 318380 319466
rect 318338 319152 318394 319161
rect 318338 319087 318394 319096
rect 318340 318912 318392 318918
rect 318340 318854 318392 318860
rect 318352 316130 318380 318854
rect 318444 317529 318472 319620
rect 318430 317520 318486 317529
rect 318430 317455 318486 317464
rect 318340 316124 318392 316130
rect 318340 316066 318392 316072
rect 318248 316056 318300 316062
rect 318248 315998 318300 316004
rect 318536 315994 318564 319892
rect 318674 319852 318702 320076
rect 318628 319824 318702 319852
rect 318524 315988 318576 315994
rect 318524 315930 318576 315936
rect 318628 315790 318656 319824
rect 318766 319784 318794 320076
rect 318858 319954 318886 320076
rect 319042 319954 319070 320076
rect 319672 320104 319728 320113
rect 319120 320039 319176 320048
rect 318858 319926 318932 319954
rect 319042 319926 319116 319954
rect 318720 319756 318794 319784
rect 318616 315784 318668 315790
rect 318616 315726 318668 315732
rect 318156 314492 318208 314498
rect 318156 314434 318208 314440
rect 318616 314492 318668 314498
rect 318616 314434 318668 314440
rect 318076 314350 318288 314378
rect 318156 313812 318208 313818
rect 318156 313754 318208 313760
rect 317878 311264 317934 311273
rect 317878 311199 317934 311208
rect 317694 306368 317750 306377
rect 317694 306303 317750 306312
rect 317708 305017 317736 306303
rect 317694 305008 317750 305017
rect 317604 304972 317656 304978
rect 317694 304943 317750 304952
rect 317604 304914 317656 304920
rect 317616 304298 317644 304914
rect 317604 304292 317656 304298
rect 317604 304234 317656 304240
rect 317418 299296 317474 299305
rect 317418 299231 317474 299240
rect 318062 299296 318118 299305
rect 318062 299231 318118 299240
rect 317420 247852 317472 247858
rect 317420 247794 317472 247800
rect 317328 244520 317380 244526
rect 317328 244462 317380 244468
rect 317340 244322 317368 244462
rect 317328 244316 317380 244322
rect 317328 244258 317380 244264
rect 316960 238264 317012 238270
rect 316960 238206 317012 238212
rect 316868 223236 316920 223242
rect 316868 223178 316920 223184
rect 316776 221944 316828 221950
rect 316776 221886 316828 221892
rect 314384 221876 314436 221882
rect 314384 221818 314436 221824
rect 314016 219224 314068 219230
rect 314016 219166 314068 219172
rect 317432 215966 317460 247794
rect 318076 244905 318104 299231
rect 318168 262857 318196 313754
rect 318260 300801 318288 314350
rect 318628 311894 318656 314434
rect 318720 314294 318748 319756
rect 318904 318753 318932 319926
rect 318982 319424 319038 319433
rect 318982 319359 319038 319368
rect 318890 318744 318946 318753
rect 318890 318679 318946 318688
rect 318904 318073 318932 318679
rect 318890 318064 318946 318073
rect 318890 317999 318946 318008
rect 318708 314288 318760 314294
rect 318708 314230 318760 314236
rect 318720 313818 318748 314230
rect 318708 313812 318760 313818
rect 318708 313754 318760 313760
rect 318628 311866 318748 311894
rect 318522 311264 318578 311273
rect 318522 311199 318578 311208
rect 318338 305008 318394 305017
rect 318338 304943 318394 304952
rect 318246 300792 318302 300801
rect 318246 300727 318302 300736
rect 318154 262848 318210 262857
rect 318154 262783 318210 262792
rect 318156 256760 318208 256766
rect 318156 256702 318208 256708
rect 318062 244896 318118 244905
rect 318062 244831 318118 244840
rect 318168 223378 318196 256702
rect 318260 250481 318288 300727
rect 318352 271182 318380 304943
rect 318340 271176 318392 271182
rect 318340 271118 318392 271124
rect 318536 260914 318564 311199
rect 318616 310276 318668 310282
rect 318616 310218 318668 310224
rect 318524 260908 318576 260914
rect 318524 260850 318576 260856
rect 318536 258074 318564 260850
rect 318352 258046 318564 258074
rect 318246 250472 318302 250481
rect 318246 250407 318302 250416
rect 318248 247716 318300 247722
rect 318248 247658 318300 247664
rect 318260 223446 318288 247658
rect 318352 238134 318380 258046
rect 318628 257378 318656 310218
rect 318616 257372 318668 257378
rect 318616 257314 318668 257320
rect 318720 256766 318748 311866
rect 318996 309097 319024 319359
rect 319088 314430 319116 319926
rect 319318 319920 319346 320076
rect 319180 319892 319346 319920
rect 319076 314424 319128 314430
rect 319076 314366 319128 314372
rect 319180 314090 319208 319892
rect 319258 319832 319314 319841
rect 319258 319767 319314 319776
rect 319272 319161 319300 319767
rect 319410 319682 319438 320076
rect 319364 319654 319438 319682
rect 319258 319152 319314 319161
rect 319258 319087 319314 319096
rect 319260 315852 319312 315858
rect 319260 315794 319312 315800
rect 319272 314974 319300 315794
rect 319260 314968 319312 314974
rect 319260 314910 319312 314916
rect 319168 314084 319220 314090
rect 319168 314026 319220 314032
rect 318982 309088 319038 309097
rect 318982 309023 319038 309032
rect 319364 297974 319392 319654
rect 319502 319580 319530 320076
rect 319594 319870 319622 320076
rect 320684 320104 320740 320113
rect 319672 320039 319728 320048
rect 319582 319864 319634 319870
rect 319582 319806 319634 319812
rect 319778 319716 319806 320076
rect 319870 319870 319898 320076
rect 319858 319864 319910 319870
rect 319858 319806 319910 319812
rect 319962 319784 319990 320076
rect 320054 319920 320082 320076
rect 320054 319892 320128 319920
rect 320100 319852 320128 319892
rect 320238 319852 320266 320076
rect 320422 319954 320450 320076
rect 320376 319926 320450 319954
rect 320100 319824 320174 319852
rect 320238 319824 320312 319852
rect 320146 319784 320174 319824
rect 319962 319756 320036 319784
rect 319778 319688 319852 319716
rect 319628 319660 319680 319666
rect 319628 319602 319680 319608
rect 319502 319552 319576 319580
rect 319548 318918 319576 319552
rect 319536 318912 319588 318918
rect 319536 318854 319588 318860
rect 319640 318794 319668 319602
rect 319720 318912 319772 318918
rect 319824 318889 319852 319688
rect 319904 319660 319956 319666
rect 319904 319602 319956 319608
rect 319720 318854 319772 318860
rect 319810 318880 319866 318889
rect 319548 318766 319668 318794
rect 319442 315208 319498 315217
rect 319442 315143 319498 315152
rect 319352 297968 319404 297974
rect 319352 297910 319404 297916
rect 318708 256760 318760 256766
rect 318708 256702 318760 256708
rect 318340 238128 318392 238134
rect 318340 238070 318392 238076
rect 319456 228410 319484 315143
rect 319548 313857 319576 318766
rect 319534 313848 319590 313857
rect 319534 313783 319590 313792
rect 319548 250753 319576 313783
rect 319628 313336 319680 313342
rect 319628 313278 319680 313284
rect 319640 305862 319668 313278
rect 319732 305969 319760 318854
rect 319810 318815 319866 318824
rect 319824 315110 319852 318815
rect 319916 318617 319944 319602
rect 319902 318608 319958 318617
rect 319902 318543 319958 318552
rect 320008 315217 320036 319756
rect 320100 319756 320174 319784
rect 320100 318918 320128 319756
rect 320178 319696 320234 319705
rect 320178 319631 320234 319640
rect 320088 318912 320140 318918
rect 320088 318854 320140 318860
rect 320100 315246 320128 318854
rect 320192 318850 320220 319631
rect 320180 318844 320232 318850
rect 320180 318786 320232 318792
rect 320284 317529 320312 319824
rect 320270 317520 320326 317529
rect 320270 317455 320326 317464
rect 320376 317422 320404 319926
rect 320514 319784 320542 320076
rect 320606 319954 320634 320076
rect 321328 320104 321384 320113
rect 320684 320039 320740 320048
rect 320606 319926 320680 319954
rect 320882 319938 320910 320076
rect 320974 319938 321002 320076
rect 320514 319756 320588 319784
rect 320454 319424 320510 319433
rect 320454 319359 320510 319368
rect 320364 317416 320416 317422
rect 320364 317358 320416 317364
rect 320178 316160 320234 316169
rect 320178 316095 320234 316104
rect 320192 315994 320220 316095
rect 320468 316062 320496 319359
rect 320456 316056 320508 316062
rect 320456 315998 320508 316004
rect 320180 315988 320232 315994
rect 320180 315930 320232 315936
rect 320456 315920 320508 315926
rect 320456 315862 320508 315868
rect 320468 315722 320496 315862
rect 320560 315722 320588 319756
rect 320652 317626 320680 319926
rect 320870 319932 320922 319938
rect 320870 319874 320922 319880
rect 320962 319932 321014 319938
rect 320962 319874 321014 319880
rect 320732 319796 320784 319802
rect 320732 319738 320784 319744
rect 320640 317620 320692 317626
rect 320640 317562 320692 317568
rect 320744 315994 320772 319738
rect 320916 319728 320968 319734
rect 321066 319682 321094 320076
rect 321158 319784 321186 320076
rect 321250 319943 321278 320076
rect 322524 320104 322580 320113
rect 321328 320039 321384 320048
rect 321236 319934 321292 319943
rect 321434 319938 321462 320076
rect 321236 319869 321292 319878
rect 321422 319932 321474 319938
rect 321526 319920 321554 320076
rect 321526 319892 321600 319920
rect 321422 319874 321474 319880
rect 321572 319818 321600 319892
rect 321710 319870 321738 320076
rect 321526 319790 321600 319818
rect 321698 319864 321750 319870
rect 321698 319806 321750 319812
rect 321158 319756 321232 319784
rect 320916 319670 320968 319676
rect 320822 319424 320878 319433
rect 320822 319359 320878 319368
rect 320732 315988 320784 315994
rect 320732 315930 320784 315936
rect 320836 315761 320864 319359
rect 320928 317937 320956 319670
rect 321020 319654 321094 319682
rect 321020 319025 321048 319654
rect 321006 319016 321062 319025
rect 321006 318951 321062 318960
rect 320914 317928 320970 317937
rect 320914 317863 320970 317872
rect 321020 317801 321048 318951
rect 321006 317792 321062 317801
rect 321006 317727 321062 317736
rect 320916 316192 320968 316198
rect 320916 316134 320968 316140
rect 320822 315752 320878 315761
rect 320456 315716 320508 315722
rect 320456 315658 320508 315664
rect 320548 315716 320600 315722
rect 320822 315687 320878 315696
rect 320548 315658 320600 315664
rect 320088 315240 320140 315246
rect 319994 315208 320050 315217
rect 320088 315182 320140 315188
rect 319994 315143 320050 315152
rect 319812 315104 319864 315110
rect 319812 315046 319864 315052
rect 320088 314424 320140 314430
rect 320088 314366 320140 314372
rect 319996 314084 320048 314090
rect 319996 314026 320048 314032
rect 319812 312452 319864 312458
rect 319812 312394 319864 312400
rect 319824 311982 319852 312394
rect 319812 311976 319864 311982
rect 319812 311918 319864 311924
rect 319718 305960 319774 305969
rect 319718 305895 319774 305904
rect 319628 305856 319680 305862
rect 319628 305798 319680 305804
rect 319628 297968 319680 297974
rect 319628 297910 319680 297916
rect 319534 250744 319590 250753
rect 319534 250679 319590 250688
rect 319640 242185 319668 297910
rect 319732 287706 319760 305895
rect 319824 304842 319852 311918
rect 319902 309088 319958 309097
rect 319902 309023 319958 309032
rect 319916 308553 319944 309023
rect 319902 308544 319958 308553
rect 319902 308479 319958 308488
rect 319812 304836 319864 304842
rect 319812 304778 319864 304784
rect 319720 287700 319772 287706
rect 319720 287642 319772 287648
rect 319720 253088 319772 253094
rect 319720 253030 319772 253036
rect 319732 252686 319760 253030
rect 319720 252680 319772 252686
rect 319720 252622 319772 252628
rect 319626 242176 319682 242185
rect 319626 242111 319682 242120
rect 319444 228404 319496 228410
rect 319444 228346 319496 228352
rect 319732 223514 319760 252622
rect 319812 251184 319864 251190
rect 319812 251126 319864 251132
rect 319824 249830 319852 251126
rect 319812 249824 319864 249830
rect 319812 249766 319864 249772
rect 319824 223582 319852 249766
rect 319916 248414 319944 308479
rect 320008 253094 320036 314026
rect 319996 253088 320048 253094
rect 319996 253030 320048 253036
rect 320100 251190 320128 314366
rect 320928 313120 320956 316134
rect 321006 315752 321062 315761
rect 321006 315687 321062 315696
rect 321100 315716 321152 315722
rect 320744 313092 320956 313120
rect 320640 312588 320692 312594
rect 320640 312530 320692 312536
rect 320652 311914 320680 312530
rect 320744 312458 320772 313092
rect 320914 313032 320970 313041
rect 320914 312967 320970 312976
rect 320732 312452 320784 312458
rect 320732 312394 320784 312400
rect 320824 312384 320876 312390
rect 320824 312326 320876 312332
rect 320640 311908 320692 311914
rect 320640 311850 320692 311856
rect 320652 307562 320680 311850
rect 320640 307556 320692 307562
rect 320640 307498 320692 307504
rect 320730 304464 320786 304473
rect 320730 304399 320786 304408
rect 320744 304298 320772 304399
rect 320732 304292 320784 304298
rect 320732 304234 320784 304240
rect 320088 251184 320140 251190
rect 320088 251126 320140 251132
rect 320088 248464 320140 248470
rect 319916 248412 320088 248414
rect 319916 248406 320140 248412
rect 319916 248386 320128 248406
rect 319916 247926 319944 248386
rect 319904 247920 319956 247926
rect 319904 247862 319956 247868
rect 320836 239494 320864 312326
rect 320928 242350 320956 312967
rect 321020 247625 321048 315687
rect 321100 315658 321152 315664
rect 321112 307737 321140 315658
rect 321204 312594 321232 319756
rect 321526 319716 321554 319790
rect 321802 319784 321830 320076
rect 321894 319852 321922 320076
rect 321986 319920 322014 320076
rect 322170 319938 322198 320076
rect 322354 319954 322382 320076
rect 322158 319932 322210 319938
rect 321986 319892 322060 319920
rect 321894 319824 321968 319852
rect 321802 319756 321876 319784
rect 321374 319696 321430 319705
rect 321284 319660 321336 319666
rect 321374 319631 321430 319640
rect 321480 319688 321554 319716
rect 321742 319696 321798 319705
rect 321284 319602 321336 319608
rect 321296 316198 321324 319602
rect 321284 316192 321336 316198
rect 321284 316134 321336 316140
rect 321284 316056 321336 316062
rect 321284 315998 321336 316004
rect 321192 312588 321244 312594
rect 321192 312530 321244 312536
rect 321296 309602 321324 315998
rect 321388 312390 321416 319631
rect 321480 313041 321508 319688
rect 321742 319631 321744 319640
rect 321796 319631 321798 319640
rect 321744 319602 321796 319608
rect 321560 319592 321612 319598
rect 321560 319534 321612 319540
rect 321652 319592 321704 319598
rect 321652 319534 321704 319540
rect 321742 319560 321798 319569
rect 321572 318345 321600 319534
rect 321558 318336 321614 318345
rect 321558 318271 321614 318280
rect 321560 316056 321612 316062
rect 321560 315998 321612 316004
rect 321466 313032 321522 313041
rect 321466 312967 321522 312976
rect 321376 312384 321428 312390
rect 321376 312326 321428 312332
rect 321284 309596 321336 309602
rect 321284 309538 321336 309544
rect 321098 307728 321154 307737
rect 321098 307663 321154 307672
rect 321112 257281 321140 307663
rect 321296 306374 321324 309538
rect 321296 306346 321508 306374
rect 321282 304328 321338 304337
rect 321282 304263 321284 304272
rect 321336 304263 321338 304272
rect 321284 304234 321336 304240
rect 321098 257272 321154 257281
rect 321098 257207 321154 257216
rect 321480 252618 321508 306346
rect 321572 301510 321600 315998
rect 321664 302734 321692 319534
rect 321742 319495 321798 319504
rect 321756 316010 321784 319495
rect 321848 319433 321876 319756
rect 321834 319424 321890 319433
rect 321834 319359 321890 319368
rect 321756 315982 321876 316010
rect 321744 315716 321796 315722
rect 321744 315658 321796 315664
rect 321756 306241 321784 315658
rect 321848 309097 321876 315982
rect 321940 310185 321968 319824
rect 322032 319802 322060 319892
rect 322158 319874 322210 319880
rect 322308 319926 322382 319954
rect 322446 319954 322474 320076
rect 324916 320104 324972 320113
rect 322524 320039 322580 320048
rect 322446 319926 322520 319954
rect 322110 319832 322166 319841
rect 322020 319796 322072 319802
rect 322110 319767 322166 319776
rect 322308 319784 322336 319926
rect 322020 319738 322072 319744
rect 322020 319660 322072 319666
rect 322020 319602 322072 319608
rect 322032 311137 322060 319602
rect 322124 319161 322152 319767
rect 322308 319756 322428 319784
rect 322294 319696 322350 319705
rect 322204 319660 322256 319666
rect 322294 319631 322350 319640
rect 322204 319602 322256 319608
rect 322110 319152 322166 319161
rect 322110 319087 322166 319096
rect 322110 319016 322166 319025
rect 322110 318951 322166 318960
rect 322124 312322 322152 318951
rect 322216 317529 322244 319602
rect 322308 318170 322336 319631
rect 322296 318164 322348 318170
rect 322296 318106 322348 318112
rect 322202 317520 322258 317529
rect 322202 317455 322258 317464
rect 322400 316849 322428 319756
rect 322492 319666 322520 319926
rect 322630 319784 322658 320076
rect 322722 319870 322750 320076
rect 322814 319938 322842 320076
rect 322802 319932 322854 319938
rect 322802 319874 322854 319880
rect 322710 319864 322762 319870
rect 322710 319806 322762 319812
rect 322906 319784 322934 320076
rect 322584 319756 322658 319784
rect 322860 319756 322934 319784
rect 322480 319660 322532 319666
rect 322480 319602 322532 319608
rect 322478 319560 322534 319569
rect 322478 319495 322534 319504
rect 322492 318782 322520 319495
rect 322480 318776 322532 318782
rect 322480 318718 322532 318724
rect 322386 316840 322442 316849
rect 322386 316775 322442 316784
rect 322584 315722 322612 319756
rect 322756 319728 322808 319734
rect 322662 319696 322718 319705
rect 322756 319670 322808 319676
rect 322662 319631 322718 319640
rect 322676 316674 322704 319631
rect 322664 316668 322716 316674
rect 322664 316610 322716 316616
rect 322572 315716 322624 315722
rect 322572 315658 322624 315664
rect 322388 313948 322440 313954
rect 322388 313890 322440 313896
rect 322112 312316 322164 312322
rect 322112 312258 322164 312264
rect 322018 311128 322074 311137
rect 322018 311063 322074 311072
rect 322124 311001 322152 312258
rect 322202 311128 322258 311137
rect 322202 311063 322258 311072
rect 322110 310992 322166 311001
rect 322110 310927 322166 310936
rect 321926 310176 321982 310185
rect 321926 310111 321982 310120
rect 321834 309088 321890 309097
rect 321834 309023 321890 309032
rect 321742 306232 321798 306241
rect 321742 306167 321798 306176
rect 321756 305017 321784 306167
rect 321742 305008 321798 305017
rect 321742 304943 321798 304952
rect 321652 302728 321704 302734
rect 321652 302670 321704 302676
rect 321652 302184 321704 302190
rect 321652 302126 321704 302132
rect 321560 301504 321612 301510
rect 321664 301481 321692 302126
rect 321560 301446 321612 301452
rect 321650 301472 321706 301481
rect 321650 301407 321706 301416
rect 321468 252612 321520 252618
rect 321468 252554 321520 252560
rect 321480 248414 321508 252554
rect 321112 248386 321508 248414
rect 321006 247616 321062 247625
rect 321006 247551 321062 247560
rect 320916 242344 320968 242350
rect 320916 242286 320968 242292
rect 320824 239488 320876 239494
rect 320824 239430 320876 239436
rect 321112 227526 321140 248386
rect 322216 243545 322244 311063
rect 322294 309088 322350 309097
rect 322294 309023 322350 309032
rect 322202 243536 322258 243545
rect 322202 243471 322258 243480
rect 322308 242894 322336 309023
rect 322400 253298 322428 313890
rect 322676 311894 322704 316610
rect 322768 313954 322796 319670
rect 322860 316062 322888 319756
rect 322998 319682 323026 320076
rect 323090 319784 323118 320076
rect 323182 319852 323210 320076
rect 323458 319954 323486 320076
rect 323642 319954 323670 320076
rect 323458 319926 323532 319954
rect 323504 319870 323532 319926
rect 323596 319926 323670 319954
rect 323492 319864 323544 319870
rect 323182 319824 323348 319852
rect 323090 319756 323164 319784
rect 322998 319654 323072 319682
rect 322938 319152 322994 319161
rect 322938 319087 322994 319096
rect 322952 318850 322980 319087
rect 322940 318844 322992 318850
rect 322940 318786 322992 318792
rect 323044 316266 323072 319654
rect 323136 318102 323164 319756
rect 323214 319696 323270 319705
rect 323214 319631 323270 319640
rect 323124 318096 323176 318102
rect 323124 318038 323176 318044
rect 323228 317937 323256 319631
rect 323214 317928 323270 317937
rect 323214 317863 323270 317872
rect 323320 316282 323348 319824
rect 323492 319806 323544 319812
rect 323400 319728 323452 319734
rect 323400 319670 323452 319676
rect 323032 316260 323084 316266
rect 323032 316202 323084 316208
rect 323228 316254 323348 316282
rect 322940 316192 322992 316198
rect 322940 316134 322992 316140
rect 322848 316056 322900 316062
rect 322848 315998 322900 316004
rect 322756 313948 322808 313954
rect 322756 313890 322808 313896
rect 322768 313750 322796 313890
rect 322756 313744 322808 313750
rect 322756 313686 322808 313692
rect 322952 311894 322980 316134
rect 323032 316056 323084 316062
rect 323032 315998 323084 316004
rect 322676 311866 322796 311894
rect 322570 310176 322626 310185
rect 322570 310111 322626 310120
rect 322480 302728 322532 302734
rect 322480 302670 322532 302676
rect 322388 253292 322440 253298
rect 322388 253234 322440 253240
rect 322492 246401 322520 302670
rect 322584 253201 322612 310111
rect 322664 301504 322716 301510
rect 322664 301446 322716 301452
rect 322676 265674 322704 301446
rect 322768 290601 322796 311866
rect 322860 311866 322980 311894
rect 322860 311114 322888 311866
rect 322860 311086 322980 311114
rect 322952 310049 322980 311086
rect 322938 310040 322994 310049
rect 322938 309975 322994 309984
rect 322952 309777 322980 309975
rect 322938 309768 322994 309777
rect 322938 309703 322994 309712
rect 323044 309097 323072 315998
rect 323228 312905 323256 316254
rect 323308 316124 323360 316130
rect 323308 316066 323360 316072
rect 323214 312896 323270 312905
rect 323214 312831 323270 312840
rect 323124 312248 323176 312254
rect 323124 312190 323176 312196
rect 323136 311302 323164 312190
rect 323124 311296 323176 311302
rect 323124 311238 323176 311244
rect 323320 310321 323348 316066
rect 323412 314673 323440 319670
rect 323492 319660 323544 319666
rect 323492 319602 323544 319608
rect 323504 319462 323532 319602
rect 323492 319456 323544 319462
rect 323492 319398 323544 319404
rect 323490 319016 323546 319025
rect 323490 318951 323546 318960
rect 323504 318209 323532 318951
rect 323490 318200 323546 318209
rect 323490 318135 323546 318144
rect 323492 316260 323544 316266
rect 323492 316202 323544 316208
rect 323398 314664 323454 314673
rect 323398 314599 323454 314608
rect 323306 310312 323362 310321
rect 323306 310247 323362 310256
rect 323030 309088 323086 309097
rect 323030 309023 323086 309032
rect 322846 305008 322902 305017
rect 322846 304943 322902 304952
rect 322754 290592 322810 290601
rect 322754 290527 322810 290536
rect 322664 265668 322716 265674
rect 322664 265610 322716 265616
rect 322570 253192 322626 253201
rect 322570 253127 322626 253136
rect 322478 246392 322534 246401
rect 322478 246327 322534 246336
rect 322860 244458 322888 304943
rect 323504 300665 323532 316202
rect 323596 314401 323624 319926
rect 323734 319784 323762 320076
rect 323918 319818 323946 320076
rect 324010 319938 324038 320076
rect 323998 319932 324050 319938
rect 323998 319874 324050 319880
rect 323918 319790 323992 319818
rect 323688 319756 323762 319784
rect 323688 316062 323716 319756
rect 323860 319728 323912 319734
rect 323860 319670 323912 319676
rect 323676 316056 323728 316062
rect 323676 315998 323728 316004
rect 323582 314392 323638 314401
rect 323582 314327 323638 314336
rect 323872 313177 323900 319670
rect 323858 313168 323914 313177
rect 323858 313103 323914 313112
rect 323490 300656 323546 300665
rect 323490 300591 323546 300600
rect 323504 296714 323532 300591
rect 323872 296714 323900 313103
rect 323964 312594 323992 319790
rect 324194 319784 324222 320076
rect 324148 319756 324222 319784
rect 324042 319696 324098 319705
rect 324042 319631 324098 319640
rect 324056 318481 324084 319631
rect 324042 318472 324098 318481
rect 324042 318407 324098 318416
rect 324044 318164 324096 318170
rect 324044 318106 324096 318112
rect 324056 318073 324084 318106
rect 324042 318064 324098 318073
rect 324042 317999 324098 318008
rect 324044 316940 324096 316946
rect 324044 316882 324096 316888
rect 324056 315722 324084 316882
rect 324148 316198 324176 319756
rect 324470 319682 324498 320076
rect 324562 319784 324590 320076
rect 324746 319954 324774 320076
rect 324700 319926 324774 319954
rect 324562 319756 324636 319784
rect 324470 319654 324544 319682
rect 324226 319016 324282 319025
rect 324226 318951 324282 318960
rect 324136 316192 324188 316198
rect 324136 316134 324188 316140
rect 324240 316130 324268 318951
rect 324516 318753 324544 319654
rect 324502 318744 324558 318753
rect 324502 318679 324558 318688
rect 324608 316470 324636 319756
rect 324596 316464 324648 316470
rect 324596 316406 324648 316412
rect 324228 316124 324280 316130
rect 324228 316066 324280 316072
rect 324412 316056 324464 316062
rect 324412 315998 324464 316004
rect 324044 315716 324096 315722
rect 324044 315658 324096 315664
rect 324134 312896 324190 312905
rect 324134 312831 324190 312840
rect 323952 312588 324004 312594
rect 323952 312530 324004 312536
rect 324042 309088 324098 309097
rect 324042 309023 324098 309032
rect 323504 296686 323624 296714
rect 322940 273964 322992 273970
rect 322940 273906 322992 273912
rect 322952 273873 322980 273906
rect 322938 273864 322994 273873
rect 322938 273799 322994 273808
rect 323596 247761 323624 296686
rect 323780 296686 323900 296714
rect 323780 287745 323808 296686
rect 323766 287736 323822 287745
rect 323766 287671 323822 287680
rect 324056 273970 324084 309023
rect 324044 273964 324096 273970
rect 324044 273906 324096 273912
rect 324148 268258 324176 312831
rect 324424 311273 324452 315998
rect 324608 314974 324636 316406
rect 324596 314968 324648 314974
rect 324596 314910 324648 314916
rect 324700 313721 324728 319926
rect 324838 319920 324866 320076
rect 326848 320104 326904 320113
rect 324916 320039 324972 320048
rect 324838 319892 324912 319920
rect 324780 318708 324832 318714
rect 324780 318650 324832 318656
rect 324792 318510 324820 318650
rect 324780 318504 324832 318510
rect 324780 318446 324832 318452
rect 324780 317620 324832 317626
rect 324780 317562 324832 317568
rect 324792 313954 324820 317562
rect 324884 317393 324912 319892
rect 325022 319818 325050 320076
rect 325114 319938 325142 320076
rect 325102 319932 325154 319938
rect 325102 319874 325154 319880
rect 325298 319870 325326 320076
rect 325286 319864 325338 319870
rect 325022 319790 325188 319818
rect 325286 319806 325338 319812
rect 325056 319728 325108 319734
rect 324962 319696 325018 319705
rect 325056 319670 325108 319676
rect 324962 319631 325018 319640
rect 324870 317384 324926 317393
rect 324870 317319 324926 317328
rect 324884 315110 324912 317319
rect 324872 315104 324924 315110
rect 324872 315046 324924 315052
rect 324780 313948 324832 313954
rect 324780 313890 324832 313896
rect 324686 313712 324742 313721
rect 324686 313647 324742 313656
rect 324976 311894 325004 319631
rect 325068 319462 325096 319670
rect 325056 319456 325108 319462
rect 325056 319398 325108 319404
rect 325054 319016 325110 319025
rect 325054 318951 325110 318960
rect 325068 316130 325096 318951
rect 325056 316124 325108 316130
rect 325056 316066 325108 316072
rect 325160 314537 325188 319790
rect 325390 319784 325418 320076
rect 325574 319920 325602 320076
rect 325528 319892 325602 319920
rect 325390 319756 325464 319784
rect 325332 319456 325384 319462
rect 325332 319398 325384 319404
rect 325238 319016 325294 319025
rect 325238 318951 325294 318960
rect 325252 317257 325280 318951
rect 325344 317626 325372 319398
rect 325436 319025 325464 319756
rect 325422 319016 325478 319025
rect 325422 318951 325478 318960
rect 325424 318844 325476 318850
rect 325424 318786 325476 318792
rect 325332 317620 325384 317626
rect 325332 317562 325384 317568
rect 325436 317490 325464 318786
rect 325424 317484 325476 317490
rect 325424 317426 325476 317432
rect 325238 317248 325294 317257
rect 325238 317183 325294 317192
rect 325146 314528 325202 314537
rect 325146 314463 325202 314472
rect 324976 311866 325096 311894
rect 324410 311264 324466 311273
rect 324410 311199 324466 311208
rect 324962 311264 325018 311273
rect 324962 311199 325018 311208
rect 324226 310312 324282 310321
rect 324226 310247 324282 310256
rect 323676 268252 323728 268258
rect 323676 268194 323728 268200
rect 324136 268252 324188 268258
rect 324136 268194 324188 268200
rect 323688 267782 323716 268194
rect 323676 267776 323728 267782
rect 323676 267718 323728 267724
rect 323582 247752 323638 247761
rect 323582 247687 323638 247696
rect 322388 244452 322440 244458
rect 322388 244394 322440 244400
rect 322848 244452 322900 244458
rect 322848 244394 322900 244400
rect 321468 242888 321520 242894
rect 321468 242830 321520 242836
rect 322296 242888 322348 242894
rect 322296 242830 322348 242836
rect 321480 241534 321508 242830
rect 321468 241528 321520 241534
rect 321468 241470 321520 241476
rect 321100 227520 321152 227526
rect 321100 227462 321152 227468
rect 319812 223576 319864 223582
rect 319812 223518 319864 223524
rect 319720 223508 319772 223514
rect 319720 223450 319772 223456
rect 318248 223440 318300 223446
rect 318248 223382 318300 223388
rect 318156 223372 318208 223378
rect 318156 223314 318208 223320
rect 317420 215960 317472 215966
rect 317420 215902 317472 215908
rect 313924 214600 313976 214606
rect 313924 214542 313976 214548
rect 311164 213240 311216 213246
rect 311164 213182 311216 213188
rect 309876 142928 309928 142934
rect 309876 142870 309928 142876
rect 309784 3936 309836 3942
rect 309784 3878 309836 3884
rect 307852 3596 307904 3602
rect 307852 3538 307904 3544
rect 309048 3596 309100 3602
rect 309048 3538 309100 3544
rect 307772 3454 307984 3482
rect 307668 3392 307720 3398
rect 307668 3334 307720 3340
rect 307116 3120 307168 3126
rect 307116 3062 307168 3068
rect 307956 480 307984 3454
rect 309060 480 309088 3538
rect 309888 3262 309916 142870
rect 311176 4010 311204 213182
rect 311898 106992 311954 107001
rect 311898 106927 311954 106936
rect 311912 16574 311940 106927
rect 311912 16546 312216 16574
rect 311164 4004 311216 4010
rect 311164 3946 311216 3952
rect 311440 3732 311492 3738
rect 311440 3674 311492 3680
rect 309876 3256 309928 3262
rect 309876 3198 309928 3204
rect 310244 3120 310296 3126
rect 310244 3062 310296 3068
rect 310256 480 310284 3062
rect 311452 480 311480 3674
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312188 354 312216 16546
rect 313936 3806 313964 214542
rect 316684 147076 316736 147082
rect 316684 147018 316736 147024
rect 314016 138848 314068 138854
rect 314016 138790 314068 138796
rect 313924 3800 313976 3806
rect 313924 3742 313976 3748
rect 314028 3738 314056 138790
rect 315302 100192 315358 100201
rect 315302 100127 315358 100136
rect 315316 4078 315344 100127
rect 315304 4072 315356 4078
rect 315304 4014 315356 4020
rect 316224 4072 316276 4078
rect 316224 4014 316276 4020
rect 314016 3732 314068 3738
rect 314016 3674 314068 3680
rect 315028 3392 315080 3398
rect 315028 3334 315080 3340
rect 313832 3256 313884 3262
rect 313832 3198 313884 3204
rect 313844 480 313872 3198
rect 315040 480 315068 3334
rect 316236 480 316264 4014
rect 316696 3602 316724 147018
rect 317432 6914 317460 215902
rect 319444 144356 319496 144362
rect 319444 144298 319496 144304
rect 318062 69592 318118 69601
rect 318062 69527 318118 69536
rect 318076 16574 318104 69527
rect 318076 16546 318196 16574
rect 317432 6886 318104 6914
rect 317328 3732 317380 3738
rect 317328 3674 317380 3680
rect 316684 3596 316736 3602
rect 316684 3538 316736 3544
rect 317340 480 317368 3674
rect 312606 354 312718 480
rect 312188 326 312718 354
rect 312606 -960 312718 326
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 6886
rect 318168 2922 318196 16546
rect 319456 4078 319484 144298
rect 320180 133340 320232 133346
rect 320180 133282 320232 133288
rect 320192 16574 320220 133282
rect 320192 16546 320496 16574
rect 319444 4072 319496 4078
rect 319444 4014 319496 4020
rect 318156 2916 318208 2922
rect 318156 2858 318208 2864
rect 319720 2916 319772 2922
rect 319720 2858 319772 2864
rect 319732 480 319760 2858
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320468 354 320496 16546
rect 321100 4072 321152 4078
rect 321100 4014 321152 4020
rect 320824 4004 320876 4010
rect 320824 3946 320876 3952
rect 320836 3738 320864 3946
rect 320824 3732 320876 3738
rect 320824 3674 320876 3680
rect 321112 3602 321140 4014
rect 321480 3602 321508 241470
rect 322400 229809 322428 244394
rect 322386 229800 322442 229809
rect 322386 229735 322442 229744
rect 323688 228954 323716 267718
rect 324240 251258 324268 310247
rect 323768 251252 323820 251258
rect 323768 251194 323820 251200
rect 324228 251252 324280 251258
rect 324228 251194 324280 251200
rect 323676 228948 323728 228954
rect 323676 228890 323728 228896
rect 323780 228750 323808 251194
rect 324976 242214 325004 311199
rect 325068 245041 325096 311866
rect 325146 302016 325202 302025
rect 325146 301951 325202 301960
rect 325160 264353 325188 301951
rect 325252 283626 325280 317183
rect 325424 316124 325476 316130
rect 325424 316066 325476 316072
rect 325330 314528 325386 314537
rect 325330 314463 325386 314472
rect 325344 313993 325372 314463
rect 325330 313984 325386 313993
rect 325330 313919 325386 313928
rect 325436 302025 325464 316066
rect 325528 315246 325556 319892
rect 325666 319818 325694 320076
rect 325850 319852 325878 320076
rect 325620 319790 325694 319818
rect 325804 319824 325878 319852
rect 325620 316062 325648 319790
rect 325700 319728 325752 319734
rect 325804 319716 325832 319824
rect 325942 319784 325970 320076
rect 326034 319920 326062 320076
rect 326034 319892 326154 319920
rect 326126 319784 326154 319892
rect 326218 319852 326246 320076
rect 326310 319954 326338 320076
rect 326310 319926 326384 319954
rect 326218 319824 326292 319852
rect 325942 319756 326016 319784
rect 326126 319756 326200 319784
rect 325804 319688 325924 319716
rect 325700 319670 325752 319676
rect 325712 318794 325740 319670
rect 325712 318766 325832 318794
rect 325896 318782 325924 319688
rect 325988 318794 326016 319756
rect 325700 317960 325752 317966
rect 325700 317902 325752 317908
rect 325608 316056 325660 316062
rect 325608 315998 325660 316004
rect 325516 315240 325568 315246
rect 325516 315182 325568 315188
rect 325608 315104 325660 315110
rect 325608 315046 325660 315052
rect 325516 314968 325568 314974
rect 325516 314910 325568 314916
rect 325422 302016 325478 302025
rect 325422 301951 325478 301960
rect 325240 283620 325292 283626
rect 325240 283562 325292 283568
rect 325146 264344 325202 264353
rect 325146 264279 325202 264288
rect 325054 245032 325110 245041
rect 325054 244967 325110 244976
rect 325528 244390 325556 314910
rect 325148 244384 325200 244390
rect 325148 244326 325200 244332
rect 325516 244384 325568 244390
rect 325516 244326 325568 244332
rect 325056 243024 325108 243030
rect 325056 242966 325108 242972
rect 324964 242208 325016 242214
rect 324964 242150 325016 242156
rect 325068 228886 325096 242966
rect 325160 229022 325188 244326
rect 325620 243030 325648 315046
rect 325712 291174 325740 317902
rect 325804 302841 325832 318766
rect 325884 318776 325936 318782
rect 325988 318766 326108 318794
rect 325884 318718 325936 318724
rect 325884 316124 325936 316130
rect 325884 316066 325936 316072
rect 325896 306105 325924 316066
rect 325976 316056 326028 316062
rect 325976 315998 326028 316004
rect 325988 307601 326016 315998
rect 326080 312769 326108 318766
rect 326172 315625 326200 319756
rect 326264 316130 326292 319824
rect 326356 319648 326384 319926
rect 326494 319920 326522 320076
rect 326448 319892 326522 319920
rect 326448 319802 326476 319892
rect 326586 319818 326614 320076
rect 326678 319938 326706 320076
rect 326666 319932 326718 319938
rect 326666 319874 326718 319880
rect 326770 319870 326798 320076
rect 327216 320104 327272 320113
rect 326848 320039 326904 320048
rect 326954 319920 326982 320076
rect 327138 319938 327166 320076
rect 327216 320039 327272 320048
rect 327126 319932 327178 319938
rect 326954 319892 327028 319920
rect 326436 319796 326488 319802
rect 326436 319738 326488 319744
rect 326540 319790 326614 319818
rect 326758 319864 326810 319870
rect 326758 319806 326810 319812
rect 326356 319620 326476 319648
rect 326342 319560 326398 319569
rect 326342 319495 326344 319504
rect 326396 319495 326398 319504
rect 326344 319466 326396 319472
rect 326252 316124 326304 316130
rect 326252 316066 326304 316072
rect 326448 316062 326476 319620
rect 326436 316056 326488 316062
rect 326436 315998 326488 316004
rect 326158 315616 326214 315625
rect 326158 315551 326214 315560
rect 326066 312760 326122 312769
rect 326066 312695 326122 312704
rect 326172 311894 326200 315551
rect 326540 314265 326568 319790
rect 326620 319728 326672 319734
rect 326620 319670 326672 319676
rect 326804 319728 326856 319734
rect 327000 319716 327028 319892
rect 327126 319874 327178 319880
rect 327080 319796 327132 319802
rect 327080 319738 327132 319744
rect 327172 319796 327224 319802
rect 327322 319784 327350 320076
rect 327552 319920 327580 330375
rect 327630 321600 327686 321609
rect 327630 321535 327686 321544
rect 327644 320793 327672 321535
rect 327630 320784 327686 320793
rect 327630 320719 327686 320728
rect 327632 320544 327684 320550
rect 327630 320512 327632 320521
rect 327684 320512 327686 320521
rect 327630 320447 327686 320456
rect 327630 320376 327686 320385
rect 327630 320311 327686 320320
rect 327644 320074 327672 320311
rect 327632 320068 327684 320074
rect 327632 320010 327684 320016
rect 327632 319932 327684 319938
rect 327552 319892 327632 319920
rect 327632 319874 327684 319880
rect 327172 319738 327224 319744
rect 327276 319756 327350 319784
rect 326856 319688 327028 319716
rect 326804 319670 326856 319676
rect 326632 317665 326660 319670
rect 326802 319560 326858 319569
rect 326802 319495 326858 319504
rect 326710 319016 326766 319025
rect 326710 318951 326766 318960
rect 326618 317656 326674 317665
rect 326618 317591 326674 317600
rect 326618 316296 326674 316305
rect 326618 316231 326674 316240
rect 326526 314256 326582 314265
rect 326526 314191 326582 314200
rect 326172 311866 326384 311894
rect 325974 307592 326030 307601
rect 325974 307527 326030 307536
rect 325882 306096 325938 306105
rect 325882 306031 325938 306040
rect 325790 302832 325846 302841
rect 325790 302767 325846 302776
rect 325700 291168 325752 291174
rect 325700 291110 325752 291116
rect 326356 249121 326384 311866
rect 326434 307592 326490 307601
rect 326434 307527 326490 307536
rect 326342 249112 326398 249121
rect 326342 249047 326398 249056
rect 326448 246265 326476 307527
rect 326540 260137 326568 314191
rect 326632 271153 326660 316231
rect 326724 309777 326752 318951
rect 326816 317121 326844 319495
rect 326802 317112 326858 317121
rect 326802 317047 326858 317056
rect 326816 316305 326844 317047
rect 326908 316713 326936 319688
rect 327092 319648 327120 319738
rect 327000 319620 327120 319648
rect 327000 317966 327028 319620
rect 327078 319560 327134 319569
rect 327184 319530 327212 319738
rect 327078 319495 327134 319504
rect 327172 319524 327224 319530
rect 326988 317960 327040 317966
rect 326988 317902 327040 317908
rect 326988 317620 327040 317626
rect 326988 317562 327040 317568
rect 327000 317529 327028 317562
rect 326986 317520 327042 317529
rect 326986 317455 327042 317464
rect 326894 316704 326950 316713
rect 326894 316639 326950 316648
rect 326802 316296 326858 316305
rect 326802 316231 326858 316240
rect 327092 313274 327120 319495
rect 327172 319466 327224 319472
rect 327172 317824 327224 317830
rect 327276 317801 327304 319756
rect 327356 319524 327408 319530
rect 327356 319466 327408 319472
rect 327368 318850 327396 319466
rect 327446 319016 327502 319025
rect 327446 318951 327502 318960
rect 327356 318844 327408 318850
rect 327356 318786 327408 318792
rect 327172 317766 327224 317772
rect 327262 317792 327318 317801
rect 327080 313268 327132 313274
rect 327080 313210 327132 313216
rect 326986 312760 327042 312769
rect 326986 312695 327042 312704
rect 326710 309768 326766 309777
rect 326710 309703 326766 309712
rect 326724 284986 326752 309703
rect 326802 306096 326858 306105
rect 326802 306031 326858 306040
rect 326816 296714 326844 306031
rect 326894 303512 326950 303521
rect 326894 303447 326950 303456
rect 326908 302841 326936 303447
rect 326894 302832 326950 302841
rect 326894 302767 326950 302776
rect 326816 296686 326936 296714
rect 326712 284980 326764 284986
rect 326712 284922 326764 284928
rect 326618 271144 326674 271153
rect 326618 271079 326674 271088
rect 326526 260128 326582 260137
rect 326526 260063 326582 260072
rect 326434 246256 326490 246265
rect 326434 246191 326490 246200
rect 326344 244316 326396 244322
rect 326344 244258 326396 244264
rect 325608 243024 325660 243030
rect 325608 242966 325660 242972
rect 326252 242956 326304 242962
rect 326252 242898 326304 242904
rect 326264 242282 326292 242898
rect 326252 242276 326304 242282
rect 326252 242218 326304 242224
rect 325148 229016 325200 229022
rect 325148 228958 325200 228964
rect 325056 228880 325108 228886
rect 326356 228857 326384 244258
rect 326908 242962 326936 296686
rect 327000 244322 327028 312695
rect 327184 253337 327212 317766
rect 327262 317727 327318 317736
rect 327264 316872 327316 316878
rect 327264 316814 327316 316820
rect 327170 253328 327226 253337
rect 327170 253263 327226 253272
rect 326988 244316 327040 244322
rect 326988 244258 327040 244264
rect 326896 242956 326948 242962
rect 326896 242898 326948 242904
rect 325056 228822 325108 228828
rect 326342 228848 326398 228857
rect 326342 228783 326398 228792
rect 323768 228744 323820 228750
rect 323768 228686 323820 228692
rect 327276 204882 327304 316814
rect 327368 315466 327396 318786
rect 327460 317830 327488 318951
rect 327448 317824 327500 317830
rect 327448 317766 327500 317772
rect 327540 317484 327592 317490
rect 327540 317426 327592 317432
rect 327368 315438 327488 315466
rect 327354 315344 327410 315353
rect 327354 315279 327410 315288
rect 327368 313721 327396 315279
rect 327354 313712 327410 313721
rect 327354 313647 327410 313656
rect 327460 313562 327488 315438
rect 327368 313534 327488 313562
rect 327368 226302 327396 313534
rect 327448 313472 327500 313478
rect 327448 313414 327500 313420
rect 327356 226296 327408 226302
rect 327356 226238 327408 226244
rect 327460 225622 327488 313414
rect 327552 308378 327580 317426
rect 327540 308372 327592 308378
rect 327540 308314 327592 308320
rect 327540 291168 327592 291174
rect 327540 291110 327592 291116
rect 327552 290494 327580 291110
rect 327540 290488 327592 290494
rect 327540 290430 327592 290436
rect 327552 229945 327580 290430
rect 327644 247897 327672 319874
rect 327736 305590 327764 398754
rect 327828 370938 327856 455738
rect 327908 453280 327960 453286
rect 327908 453222 327960 453228
rect 327816 370932 327868 370938
rect 327816 370874 327868 370880
rect 327920 368626 327948 453222
rect 329196 398608 329248 398614
rect 329196 398550 329248 398556
rect 329104 396976 329156 396982
rect 329104 396918 329156 396924
rect 328000 389020 328052 389026
rect 328000 388962 328052 388968
rect 327908 368620 327960 368626
rect 327908 368562 327960 368568
rect 327814 358048 327870 358057
rect 327814 357983 327870 357992
rect 327828 321162 327856 357983
rect 328012 345014 328040 388962
rect 328368 372088 328420 372094
rect 328368 372030 328420 372036
rect 328380 366489 328408 372030
rect 328366 366480 328422 366489
rect 328366 366415 328422 366424
rect 328012 344986 328316 345014
rect 327906 341592 327962 341601
rect 327906 341527 327962 341536
rect 327920 321434 327948 341527
rect 327998 327720 328054 327729
rect 327998 327655 328054 327664
rect 327908 321428 327960 321434
rect 327908 321370 327960 321376
rect 327906 321192 327962 321201
rect 327816 321156 327868 321162
rect 327906 321127 327962 321136
rect 327816 321098 327868 321104
rect 327814 321056 327870 321065
rect 327814 320991 327870 321000
rect 327828 320521 327856 320991
rect 327814 320512 327870 320521
rect 327814 320447 327870 320456
rect 327920 320385 327948 321127
rect 327906 320376 327962 320385
rect 327906 320311 327962 320320
rect 328012 317801 328040 327655
rect 328184 321428 328236 321434
rect 328184 321370 328236 321376
rect 328092 321156 328144 321162
rect 328092 321098 328144 321104
rect 328104 318306 328132 321098
rect 328092 318300 328144 318306
rect 328092 318242 328144 318248
rect 328196 318238 328224 321370
rect 328288 320142 328316 344986
rect 329012 338768 329064 338774
rect 329012 338710 329064 338716
rect 329024 325694 329052 338710
rect 328932 325666 329052 325694
rect 328366 321464 328422 321473
rect 328366 321399 328422 321408
rect 328380 321201 328408 321399
rect 328366 321192 328422 321201
rect 328366 321127 328422 321136
rect 328276 320136 328328 320142
rect 328276 320078 328328 320084
rect 328184 318232 328236 318238
rect 328184 318174 328236 318180
rect 327998 317792 328054 317801
rect 327998 317727 328054 317736
rect 328196 317490 328224 318174
rect 328380 317642 328408 321127
rect 328460 320680 328512 320686
rect 328460 320622 328512 320628
rect 328472 320278 328500 320622
rect 328460 320272 328512 320278
rect 328460 320214 328512 320220
rect 328932 320113 328960 325666
rect 329116 321554 329144 396918
rect 329024 321526 329144 321554
rect 328918 320104 328974 320113
rect 328918 320039 328974 320048
rect 328736 318300 328788 318306
rect 328736 318242 328788 318248
rect 328644 318164 328696 318170
rect 328644 318106 328696 318112
rect 328460 318028 328512 318034
rect 328460 317970 328512 317976
rect 328288 317614 328408 317642
rect 328184 317484 328236 317490
rect 328184 317426 328236 317432
rect 328288 313478 328316 317614
rect 328368 317484 328420 317490
rect 328368 317426 328420 317432
rect 328380 316962 328408 317426
rect 328472 317082 328500 317970
rect 328552 317960 328604 317966
rect 328552 317902 328604 317908
rect 328460 317076 328512 317082
rect 328460 317018 328512 317024
rect 328564 317014 328592 317902
rect 328552 317008 328604 317014
rect 328380 316934 328500 316962
rect 328552 316950 328604 316956
rect 328472 316826 328500 316934
rect 328472 316798 328592 316826
rect 328458 316704 328514 316713
rect 328458 316639 328514 316648
rect 328276 313472 328328 313478
rect 328276 313414 328328 313420
rect 327816 313268 327868 313274
rect 327816 313210 327868 313216
rect 327724 305584 327776 305590
rect 327724 305526 327776 305532
rect 327630 247888 327686 247897
rect 327630 247823 327686 247832
rect 327828 238754 327856 313210
rect 328472 309641 328500 316639
rect 328458 309632 328514 309641
rect 328458 309567 328514 309576
rect 328460 309528 328512 309534
rect 328460 309470 328512 309476
rect 327736 238726 327856 238754
rect 327736 236434 327764 238726
rect 327724 236428 327776 236434
rect 327724 236370 327776 236376
rect 327538 229936 327594 229945
rect 327538 229871 327594 229880
rect 327448 225616 327500 225622
rect 327448 225558 327500 225564
rect 327264 204876 327316 204882
rect 327264 204818 327316 204824
rect 325700 175296 325752 175302
rect 325700 175238 325752 175244
rect 324412 158024 324464 158030
rect 324412 157966 324464 157972
rect 323584 141568 323636 141574
rect 323584 141510 323636 141516
rect 322938 13016 322994 13025
rect 322938 12951 322994 12960
rect 322112 4140 322164 4146
rect 322112 4082 322164 4088
rect 321100 3596 321152 3602
rect 321100 3538 321152 3544
rect 321468 3596 321520 3602
rect 321468 3538 321520 3544
rect 322124 480 322152 4082
rect 320886 354 320998 480
rect 320468 326 320998 354
rect 320886 -960 320998 326
rect 322082 -960 322194 480
rect 322952 354 322980 12951
rect 323596 4146 323624 141510
rect 323584 4140 323636 4146
rect 323584 4082 323636 4088
rect 324320 3868 324372 3874
rect 324320 3810 324372 3816
rect 324332 1986 324360 3810
rect 324424 3398 324452 157966
rect 325712 16574 325740 175238
rect 327080 149796 327132 149802
rect 327080 149738 327132 149744
rect 327092 16574 327120 149738
rect 325712 16546 326384 16574
rect 327092 16546 327672 16574
rect 324412 3392 324464 3398
rect 324412 3334 324464 3340
rect 325608 3392 325660 3398
rect 325608 3334 325660 3340
rect 324332 1958 324452 1986
rect 324424 480 324452 1958
rect 325620 480 325648 3334
rect 323278 354 323390 480
rect 322952 326 323390 354
rect 323278 -960 323390 326
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326356 354 326384 16546
rect 327540 4140 327592 4146
rect 327540 4082 327592 4088
rect 327552 3398 327580 4082
rect 327644 3482 327672 16546
rect 327736 3874 327764 236370
rect 328472 222154 328500 309470
rect 328564 227186 328592 316798
rect 328656 315654 328684 318106
rect 328644 315648 328696 315654
rect 328644 315590 328696 315596
rect 328644 315308 328696 315314
rect 328644 315250 328696 315256
rect 328656 309534 328684 315250
rect 328748 315042 328776 318242
rect 328828 318232 328880 318238
rect 328828 318174 328880 318180
rect 328736 315036 328788 315042
rect 328736 314978 328788 314984
rect 328840 312662 328868 318174
rect 328932 317937 328960 320039
rect 328918 317928 328974 317937
rect 328918 317863 328974 317872
rect 329024 313206 329052 321526
rect 329208 320090 329236 398550
rect 330482 398440 330538 398449
rect 330482 398375 330538 398384
rect 329288 391604 329340 391610
rect 329288 391546 329340 391552
rect 329116 320062 329236 320090
rect 329116 316538 329144 320062
rect 329194 319968 329250 319977
rect 329194 319903 329250 319912
rect 329208 319433 329236 319903
rect 329194 319424 329250 319433
rect 329194 319359 329250 319368
rect 329194 318336 329250 318345
rect 329194 318271 329250 318280
rect 329104 316532 329156 316538
rect 329104 316474 329156 316480
rect 329208 316402 329236 318271
rect 329300 316606 329328 391546
rect 329472 386096 329524 386102
rect 329378 386064 329434 386073
rect 329472 386038 329524 386044
rect 329378 385999 329434 386008
rect 329392 319784 329420 385999
rect 329484 321554 329512 386038
rect 329656 372156 329708 372162
rect 329656 372098 329708 372104
rect 329668 365702 329696 372098
rect 329748 366376 329800 366382
rect 329748 366318 329800 366324
rect 329656 365696 329708 365702
rect 329656 365638 329708 365644
rect 329656 359508 329708 359514
rect 329656 359450 329708 359456
rect 329484 321526 329604 321554
rect 329392 319756 329512 319784
rect 329484 318646 329512 319756
rect 329576 318714 329604 321526
rect 329668 318782 329696 359450
rect 329656 318776 329708 318782
rect 329760 318753 329788 366318
rect 330298 323776 330354 323785
rect 330298 323711 330354 323720
rect 330312 322969 330340 323711
rect 329838 322960 329894 322969
rect 329838 322895 329894 322904
rect 330298 322960 330354 322969
rect 330298 322895 330354 322904
rect 329656 318718 329708 318724
rect 329746 318744 329802 318753
rect 329564 318708 329616 318714
rect 329564 318650 329616 318656
rect 329472 318640 329524 318646
rect 329472 318582 329524 318588
rect 329378 318064 329434 318073
rect 329378 317999 329434 318008
rect 329392 316606 329420 317999
rect 329288 316600 329340 316606
rect 329288 316542 329340 316548
rect 329380 316600 329432 316606
rect 329380 316542 329432 316548
rect 329196 316396 329248 316402
rect 329196 316338 329248 316344
rect 329208 316305 329236 316338
rect 329194 316296 329250 316305
rect 329194 316231 329250 316240
rect 329392 316169 329420 316542
rect 329378 316160 329434 316169
rect 329378 316095 329434 316104
rect 329012 313200 329064 313206
rect 329012 313142 329064 313148
rect 328828 312656 328880 312662
rect 328828 312598 328880 312604
rect 329484 311894 329512 318582
rect 329576 317490 329604 318650
rect 329668 318617 329696 318718
rect 329746 318679 329802 318688
rect 329654 318608 329710 318617
rect 329654 318543 329710 318552
rect 329760 317665 329788 318679
rect 329746 317656 329802 317665
rect 329746 317591 329802 317600
rect 329564 317484 329616 317490
rect 329564 317426 329616 317432
rect 329392 311866 329512 311894
rect 329010 311400 329066 311409
rect 329010 311335 329066 311344
rect 329024 311137 329052 311335
rect 329010 311128 329066 311137
rect 329010 311063 329066 311072
rect 328644 309528 328696 309534
rect 328644 309470 328696 309476
rect 329392 307018 329420 311866
rect 329380 307012 329432 307018
rect 329380 306954 329432 306960
rect 329852 228993 329880 322895
rect 330206 321328 330262 321337
rect 330206 321263 330262 321272
rect 329932 320000 329984 320006
rect 329932 319942 329984 319948
rect 329944 319462 329972 319942
rect 329932 319456 329984 319462
rect 329932 319398 329984 319404
rect 330116 319456 330168 319462
rect 330116 319398 330168 319404
rect 329930 318064 329986 318073
rect 329930 317999 329986 318008
rect 329944 313886 329972 317999
rect 330024 313948 330076 313954
rect 330024 313890 330076 313896
rect 329932 313880 329984 313886
rect 329932 313822 329984 313828
rect 329932 313676 329984 313682
rect 329932 313618 329984 313624
rect 329944 232694 329972 313618
rect 330036 235958 330064 313890
rect 330128 313682 330156 319398
rect 330116 313676 330168 313682
rect 330116 313618 330168 313624
rect 330220 313274 330248 321263
rect 330208 313268 330260 313274
rect 330208 313210 330260 313216
rect 330116 312588 330168 312594
rect 330116 312530 330168 312536
rect 330128 237318 330156 312530
rect 330390 310448 330446 310457
rect 330390 310383 330446 310392
rect 330404 310185 330432 310383
rect 330390 310176 330446 310185
rect 330390 310111 330446 310120
rect 330496 305522 330524 398375
rect 331954 397352 332010 397361
rect 331954 397287 332010 397296
rect 330758 397216 330814 397225
rect 330758 397151 330814 397160
rect 330574 396536 330630 396545
rect 330574 396471 330630 396480
rect 330484 305516 330536 305522
rect 330484 305458 330536 305464
rect 330588 305386 330616 396471
rect 330668 386164 330720 386170
rect 330668 386106 330720 386112
rect 330576 305380 330628 305386
rect 330576 305322 330628 305328
rect 330680 304978 330708 386106
rect 330772 317218 330800 397151
rect 331864 395752 331916 395758
rect 331864 395694 331916 395700
rect 330944 395684 330996 395690
rect 330944 395626 330996 395632
rect 330852 387320 330904 387326
rect 330852 387262 330904 387268
rect 330760 317212 330812 317218
rect 330760 317154 330812 317160
rect 330864 311681 330892 387262
rect 330956 321337 330984 395626
rect 331036 383376 331088 383382
rect 331036 383318 331088 383324
rect 330942 321328 330998 321337
rect 330942 321263 330998 321272
rect 331048 317422 331076 383318
rect 331128 329112 331180 329118
rect 331128 329054 331180 329060
rect 331140 317898 331168 329054
rect 331218 327176 331274 327185
rect 331218 327111 331274 327120
rect 331128 317892 331180 317898
rect 331128 317834 331180 317840
rect 331036 317416 331088 317422
rect 331036 317358 331088 317364
rect 330850 311672 330906 311681
rect 330850 311607 330906 311616
rect 330758 310040 330814 310049
rect 330758 309975 330814 309984
rect 330772 309777 330800 309975
rect 330758 309768 330814 309777
rect 330758 309703 330814 309712
rect 330668 304972 330720 304978
rect 330668 304914 330720 304920
rect 330116 237312 330168 237318
rect 330116 237254 330168 237260
rect 330024 235952 330076 235958
rect 330024 235894 330076 235900
rect 329932 232688 329984 232694
rect 329932 232630 329984 232636
rect 331232 231849 331260 327111
rect 331678 320104 331734 320113
rect 331678 320039 331734 320048
rect 331310 318608 331366 318617
rect 331310 318543 331366 318552
rect 331324 234025 331352 318543
rect 331494 318200 331550 318209
rect 331494 318135 331550 318144
rect 331404 318096 331456 318102
rect 331404 318038 331456 318044
rect 331416 235278 331444 318038
rect 331404 235272 331456 235278
rect 331508 235249 331536 318135
rect 331692 317218 331720 320039
rect 331772 318776 331824 318782
rect 331772 318718 331824 318724
rect 331784 318102 331812 318718
rect 331772 318096 331824 318102
rect 331772 318038 331824 318044
rect 331680 317212 331732 317218
rect 331680 317154 331732 317160
rect 331692 316334 331720 317154
rect 331680 316328 331732 316334
rect 331680 316270 331732 316276
rect 331876 303346 331904 395694
rect 331968 311030 331996 397287
rect 332060 374746 332088 456894
rect 332232 449948 332284 449954
rect 332232 449890 332284 449896
rect 332140 394256 332192 394262
rect 332140 394198 332192 394204
rect 332048 374740 332100 374746
rect 332048 374682 332100 374688
rect 332048 347064 332100 347070
rect 332048 347006 332100 347012
rect 332060 318374 332088 347006
rect 332048 318368 332100 318374
rect 332048 318310 332100 318316
rect 332152 317354 332180 394198
rect 332244 373386 332272 449890
rect 333336 400580 333388 400586
rect 333336 400522 333388 400528
rect 333244 397044 333296 397050
rect 333244 396986 333296 396992
rect 332324 392896 332376 392902
rect 332324 392838 332376 392844
rect 332232 373380 332284 373386
rect 332232 373322 332284 373328
rect 332232 342916 332284 342922
rect 332232 342858 332284 342864
rect 332244 318578 332272 342858
rect 332336 319734 332364 392838
rect 332416 383308 332468 383314
rect 332416 383250 332468 383256
rect 332324 319728 332376 319734
rect 332324 319670 332376 319676
rect 332232 318572 332284 318578
rect 332232 318514 332284 318520
rect 332322 318200 332378 318209
rect 332322 318135 332378 318144
rect 332336 318102 332364 318135
rect 332324 318096 332376 318102
rect 332324 318038 332376 318044
rect 332140 317348 332192 317354
rect 332140 317290 332192 317296
rect 332048 316328 332100 316334
rect 332048 316270 332100 316276
rect 331956 311024 332008 311030
rect 331956 310966 332008 310972
rect 331864 303340 331916 303346
rect 331864 303282 331916 303288
rect 332060 236609 332088 316270
rect 332428 314673 332456 383250
rect 332784 371884 332836 371890
rect 332784 371826 332836 371832
rect 332600 371544 332652 371550
rect 332600 371486 332652 371492
rect 332612 371414 332640 371486
rect 332600 371408 332652 371414
rect 332600 371350 332652 371356
rect 332508 340196 332560 340202
rect 332508 340138 332560 340144
rect 332520 317694 332548 340138
rect 332508 317688 332560 317694
rect 332508 317630 332560 317636
rect 332414 314664 332470 314673
rect 332414 314599 332470 314608
rect 332612 309874 332640 371350
rect 332796 371278 332824 371826
rect 332784 371272 332836 371278
rect 332784 371214 332836 371220
rect 332690 317656 332746 317665
rect 332690 317591 332746 317600
rect 332600 309868 332652 309874
rect 332600 309810 332652 309816
rect 332600 250504 332652 250510
rect 332600 250446 332652 250452
rect 332046 236600 332102 236609
rect 332046 236535 332102 236544
rect 331404 235214 331456 235220
rect 331494 235240 331550 235249
rect 331494 235175 331550 235184
rect 331310 234016 331366 234025
rect 331310 233951 331366 233960
rect 331218 231840 331274 231849
rect 331218 231775 331274 231784
rect 329838 228984 329894 228993
rect 329838 228919 329894 228928
rect 328552 227180 328604 227186
rect 328552 227122 328604 227128
rect 328460 222148 328512 222154
rect 328460 222090 328512 222096
rect 327816 204876 327868 204882
rect 327816 204818 327868 204824
rect 327828 4078 327856 204818
rect 332612 203658 332640 250446
rect 332704 235385 332732 317591
rect 332796 309942 332824 371214
rect 333152 320952 333204 320958
rect 333152 320894 333204 320900
rect 333164 320754 333192 320894
rect 333152 320748 333204 320754
rect 333152 320690 333204 320696
rect 332874 319288 332930 319297
rect 332874 319223 332930 319232
rect 332784 309936 332836 309942
rect 332784 309878 332836 309884
rect 332784 307012 332836 307018
rect 332784 306954 332836 306960
rect 332690 235376 332746 235385
rect 332690 235311 332746 235320
rect 332796 231266 332824 306954
rect 332888 233209 332916 319223
rect 333256 300014 333284 396986
rect 333348 311166 333376 400522
rect 333428 397248 333480 397254
rect 333428 397190 333480 397196
rect 333336 311160 333388 311166
rect 333336 311102 333388 311108
rect 333440 309670 333468 397190
rect 333532 371550 333560 456962
rect 334624 454640 334676 454646
rect 334624 454582 334676 454588
rect 333888 400444 333940 400450
rect 333888 400386 333940 400392
rect 333900 400178 333928 400386
rect 333888 400172 333940 400178
rect 333888 400114 333940 400120
rect 334348 399968 334400 399974
rect 334348 399910 334400 399916
rect 333796 399288 333848 399294
rect 333796 399230 333848 399236
rect 333612 392964 333664 392970
rect 333612 392906 333664 392912
rect 333520 371544 333572 371550
rect 333520 371486 333572 371492
rect 333520 359576 333572 359582
rect 333520 359518 333572 359524
rect 333532 318442 333560 359518
rect 333520 318436 333572 318442
rect 333520 318378 333572 318384
rect 333624 316033 333652 392906
rect 333704 386028 333756 386034
rect 333704 385970 333756 385976
rect 333610 316024 333666 316033
rect 333610 315959 333666 315968
rect 333520 313268 333572 313274
rect 333520 313210 333572 313216
rect 333428 309664 333480 309670
rect 333428 309606 333480 309612
rect 333244 300008 333296 300014
rect 333244 299950 333296 299956
rect 333532 237289 333560 313210
rect 333716 312769 333744 385970
rect 333808 370598 333836 399230
rect 334360 395418 334388 399910
rect 334348 395412 334400 395418
rect 334348 395354 334400 395360
rect 334636 372366 334664 454582
rect 334728 404258 334756 457098
rect 334900 457088 334952 457094
rect 334900 457030 334952 457036
rect 334808 451648 334860 451654
rect 334808 451590 334860 451596
rect 334820 407046 334848 451590
rect 334912 420918 334940 457030
rect 336464 455864 336516 455870
rect 336464 455806 336516 455812
rect 335084 453484 335136 453490
rect 335084 453426 335136 453432
rect 334990 450256 335046 450265
rect 334990 450191 335046 450200
rect 334900 420912 334952 420918
rect 334900 420854 334952 420860
rect 334808 407040 334860 407046
rect 334808 406982 334860 406988
rect 334716 404252 334768 404258
rect 334716 404194 334768 404200
rect 334900 399764 334952 399770
rect 334900 399706 334952 399712
rect 334716 399356 334768 399362
rect 334716 399298 334768 399304
rect 334624 372360 334676 372366
rect 334624 372302 334676 372308
rect 333978 371920 334034 371929
rect 333978 371855 334034 371864
rect 333992 371346 334020 371855
rect 333980 371340 334032 371346
rect 333980 371282 334032 371288
rect 333796 370592 333848 370598
rect 333796 370534 333848 370540
rect 333992 364334 334020 371282
rect 334622 368792 334678 368801
rect 334622 368727 334678 368736
rect 333992 364306 334204 364334
rect 333796 356720 333848 356726
rect 333796 356662 333848 356668
rect 333808 317558 333836 356662
rect 334072 322244 334124 322250
rect 334072 322186 334124 322192
rect 334084 321554 334112 322186
rect 333992 321526 334112 321554
rect 333992 319977 334020 321526
rect 333978 319968 334034 319977
rect 333978 319903 334034 319912
rect 333886 319696 333942 319705
rect 333886 319631 333942 319640
rect 333900 319297 333928 319631
rect 333886 319288 333942 319297
rect 333886 319223 333942 319232
rect 333796 317552 333848 317558
rect 333796 317494 333848 317500
rect 333888 315240 333940 315246
rect 333888 315182 333940 315188
rect 333900 313274 333928 315182
rect 333888 313268 333940 313274
rect 333888 313210 333940 313216
rect 333702 312760 333758 312769
rect 333702 312695 333758 312704
rect 333518 237280 333574 237289
rect 333518 237215 333574 237224
rect 332874 233200 332930 233209
rect 332874 233135 332930 233144
rect 333992 233073 334020 319903
rect 334070 315480 334126 315489
rect 334070 315415 334126 315424
rect 333978 233064 334034 233073
rect 333978 232999 334034 233008
rect 334084 232626 334112 315415
rect 334176 291854 334204 364306
rect 334530 320648 334586 320657
rect 334530 320583 334586 320592
rect 334544 320385 334572 320583
rect 334530 320376 334586 320385
rect 334530 320311 334586 320320
rect 334256 312656 334308 312662
rect 334254 312624 334256 312633
rect 334308 312624 334310 312633
rect 334254 312559 334310 312568
rect 334164 291848 334216 291854
rect 334164 291790 334216 291796
rect 334268 237969 334296 312559
rect 334254 237960 334310 237969
rect 334254 237895 334310 237904
rect 334072 232620 334124 232626
rect 334072 232562 334124 232568
rect 332784 231260 332836 231266
rect 332784 231202 332836 231208
rect 332600 203652 332652 203658
rect 332600 203594 332652 203600
rect 332612 16574 332640 203594
rect 334636 20670 334664 368727
rect 334728 303142 334756 399298
rect 334808 397316 334860 397322
rect 334808 397258 334860 397264
rect 334820 304502 334848 397258
rect 334912 395554 334940 399706
rect 334900 395548 334952 395554
rect 334900 395490 334952 395496
rect 334898 395176 334954 395185
rect 334898 395111 334954 395120
rect 334912 309126 334940 395111
rect 335004 368393 335032 450191
rect 335096 372502 335124 453426
rect 336188 400512 336240 400518
rect 335910 400480 335966 400489
rect 336188 400454 336240 400460
rect 335910 400415 335966 400424
rect 335820 399832 335872 399838
rect 335820 399774 335872 399780
rect 335636 399696 335688 399702
rect 335636 399638 335688 399644
rect 335648 398206 335676 399638
rect 335636 398200 335688 398206
rect 335636 398142 335688 398148
rect 335832 395865 335860 399774
rect 335818 395856 335874 395865
rect 335818 395791 335874 395800
rect 335268 388884 335320 388890
rect 335268 388826 335320 388832
rect 335084 372496 335136 372502
rect 335084 372438 335136 372444
rect 334990 368384 335046 368393
rect 334990 368319 335046 368328
rect 334992 362228 335044 362234
rect 334992 362170 335044 362176
rect 335004 317762 335032 362170
rect 335176 333260 335228 333266
rect 335176 333202 335228 333208
rect 335084 323604 335136 323610
rect 335084 323546 335136 323552
rect 334992 317756 335044 317762
rect 334992 317698 335044 317704
rect 334990 317520 335046 317529
rect 334990 317455 335046 317464
rect 335004 317422 335032 317455
rect 334992 317416 335044 317422
rect 334992 317358 335044 317364
rect 334900 309120 334952 309126
rect 334900 309062 334952 309068
rect 334808 304496 334860 304502
rect 334808 304438 334860 304444
rect 334716 303136 334768 303142
rect 334716 303078 334768 303084
rect 335004 236706 335032 317358
rect 335096 297430 335124 323546
rect 335188 315489 335216 333202
rect 335280 322538 335308 388826
rect 335280 322510 335492 322538
rect 335464 320278 335492 322510
rect 335924 321554 335952 400415
rect 336096 395140 336148 395146
rect 336096 395082 336148 395088
rect 336004 395072 336056 395078
rect 336004 395014 336056 395020
rect 335556 321526 335952 321554
rect 335556 320414 335584 321526
rect 335544 320408 335596 320414
rect 335544 320350 335596 320356
rect 335452 320272 335504 320278
rect 335452 320214 335504 320220
rect 335360 319796 335412 319802
rect 335360 319738 335412 319744
rect 335372 318850 335400 319738
rect 335360 318844 335412 318850
rect 335360 318786 335412 318792
rect 335174 315480 335230 315489
rect 335174 315415 335230 315424
rect 335084 297424 335136 297430
rect 335084 297366 335136 297372
rect 334992 236700 335044 236706
rect 334992 236642 335044 236648
rect 335372 227118 335400 318786
rect 335464 229770 335492 320214
rect 335556 233889 335584 320350
rect 336016 300762 336044 395014
rect 336108 301442 336136 395082
rect 336200 307086 336228 400454
rect 336280 399424 336332 399430
rect 336280 399366 336332 399372
rect 336188 307080 336240 307086
rect 336188 307022 336240 307028
rect 336292 306882 336320 399366
rect 336372 396364 336424 396370
rect 336372 396306 336424 396312
rect 336280 306876 336332 306882
rect 336280 306818 336332 306824
rect 336384 305794 336412 396306
rect 336476 370870 336504 455806
rect 350724 454980 350776 454986
rect 350724 454922 350776 454928
rect 337936 454776 337988 454782
rect 337936 454718 337988 454724
rect 337474 454200 337530 454209
rect 337474 454135 337530 454144
rect 337384 451784 337436 451790
rect 337384 451726 337436 451732
rect 337396 406434 337424 451726
rect 337488 413982 337516 454135
rect 337658 454064 337714 454073
rect 337658 453999 337714 454008
rect 337672 419490 337700 453999
rect 337844 453620 337896 453626
rect 337844 453562 337896 453568
rect 337660 419484 337712 419490
rect 337660 419426 337712 419432
rect 337476 413976 337528 413982
rect 337476 413918 337528 413924
rect 337384 406428 337436 406434
rect 337384 406370 337436 406376
rect 336554 400344 336610 400353
rect 336554 400279 336610 400288
rect 336464 370864 336516 370870
rect 336464 370806 336516 370812
rect 336464 334620 336516 334626
rect 336464 334562 336516 334568
rect 336476 318850 336504 334562
rect 336464 318844 336516 318850
rect 336464 318786 336516 318792
rect 336568 316606 336596 400279
rect 337660 398880 337712 398886
rect 337660 398822 337712 398828
rect 337476 397180 337528 397186
rect 337476 397122 337528 397128
rect 336648 396908 336700 396914
rect 336648 396850 336700 396856
rect 336556 316600 336608 316606
rect 336556 316542 336608 316548
rect 336660 316402 336688 396850
rect 337384 391808 337436 391814
rect 337384 391750 337436 391756
rect 336924 326392 336976 326398
rect 336924 326334 336976 326340
rect 336738 321600 336794 321609
rect 336738 321535 336794 321544
rect 336648 316396 336700 316402
rect 336648 316338 336700 316344
rect 336372 305788 336424 305794
rect 336372 305730 336424 305736
rect 336096 301436 336148 301442
rect 336096 301378 336148 301384
rect 336004 300756 336056 300762
rect 336004 300698 336056 300704
rect 336188 300076 336240 300082
rect 336188 300018 336240 300024
rect 336200 298858 336228 300018
rect 336188 298852 336240 298858
rect 336188 298794 336240 298800
rect 336200 296714 336228 298794
rect 336016 296686 336228 296714
rect 335542 233880 335598 233889
rect 335542 233815 335598 233824
rect 335452 229764 335504 229770
rect 335452 229706 335504 229712
rect 335360 227112 335412 227118
rect 335360 227054 335412 227060
rect 336016 218754 336044 296686
rect 336752 227497 336780 321535
rect 336830 320376 336886 320385
rect 336830 320311 336886 320320
rect 336844 227633 336872 320311
rect 336936 320249 336964 326334
rect 337016 321088 337068 321094
rect 337016 321030 337068 321036
rect 336922 320240 336978 320249
rect 337028 320210 337056 321030
rect 336922 320175 336978 320184
rect 337016 320204 337068 320210
rect 336936 231198 336964 320175
rect 337016 320146 337068 320152
rect 337028 232558 337056 320146
rect 337396 297566 337424 391750
rect 337488 302802 337516 397122
rect 337568 397112 337620 397118
rect 337568 397054 337620 397060
rect 337580 309058 337608 397054
rect 337672 313954 337700 398822
rect 337752 397792 337804 397798
rect 337752 397734 337804 397740
rect 337764 314566 337792 397734
rect 337856 370666 337884 453562
rect 337948 372434 337976 454718
rect 338028 454708 338080 454714
rect 338028 454650 338080 454656
rect 338040 373454 338068 454650
rect 349988 454572 350040 454578
rect 349988 454514 350040 454520
rect 340788 454232 340840 454238
rect 340788 454174 340840 454180
rect 340512 454096 340564 454102
rect 340512 454038 340564 454044
rect 340144 452056 340196 452062
rect 340144 451998 340196 452004
rect 338764 451716 338816 451722
rect 338764 451658 338816 451664
rect 338776 409154 338804 451658
rect 339316 450084 339368 450090
rect 339316 450026 339368 450032
rect 338764 409148 338816 409154
rect 338764 409090 338816 409096
rect 338948 399152 339000 399158
rect 338948 399094 339000 399100
rect 338764 396024 338816 396030
rect 338764 395966 338816 395972
rect 338672 395276 338724 395282
rect 338672 395218 338724 395224
rect 338580 391672 338632 391678
rect 338580 391614 338632 391620
rect 338028 373448 338080 373454
rect 338028 373390 338080 373396
rect 337936 372428 337988 372434
rect 337936 372370 337988 372376
rect 337844 370660 337896 370666
rect 337844 370602 337896 370608
rect 337934 325136 337990 325145
rect 337934 325071 337990 325080
rect 337948 320385 337976 325071
rect 338210 321056 338266 321065
rect 338210 320991 338266 321000
rect 338118 320648 338174 320657
rect 338118 320583 338174 320592
rect 337934 320376 337990 320385
rect 337934 320311 337990 320320
rect 338132 320249 338160 320583
rect 338118 320240 338174 320249
rect 338118 320175 338174 320184
rect 337752 314560 337804 314566
rect 337752 314502 337804 314508
rect 337660 313948 337712 313954
rect 337660 313890 337712 313896
rect 337568 309052 337620 309058
rect 337568 308994 337620 309000
rect 337476 302796 337528 302802
rect 337476 302738 337528 302744
rect 337384 297560 337436 297566
rect 337384 297502 337436 297508
rect 337016 232552 337068 232558
rect 337016 232494 337068 232500
rect 336924 231192 336976 231198
rect 336924 231134 336976 231140
rect 336830 227624 336886 227633
rect 336830 227559 336886 227568
rect 336738 227488 336794 227497
rect 336738 227423 336794 227432
rect 338132 227050 338160 320175
rect 338224 319161 338252 320991
rect 338210 319152 338266 319161
rect 338266 319110 338436 319138
rect 338210 319087 338266 319096
rect 338210 316568 338266 316577
rect 338210 316503 338266 316512
rect 338120 227044 338172 227050
rect 338120 226986 338172 226992
rect 338224 226846 338252 316503
rect 338304 315580 338356 315586
rect 338304 315522 338356 315528
rect 338316 231130 338344 315522
rect 338408 238066 338436 319110
rect 338592 317966 338620 391614
rect 338580 317960 338632 317966
rect 338580 317902 338632 317908
rect 338684 317422 338712 395218
rect 338672 317416 338724 317422
rect 338672 317358 338724 317364
rect 338776 300150 338804 395966
rect 338856 393100 338908 393106
rect 338856 393042 338908 393048
rect 338764 300144 338816 300150
rect 338764 300086 338816 300092
rect 338868 298994 338896 393042
rect 338960 306950 338988 399094
rect 339222 397896 339278 397905
rect 339222 397831 339278 397840
rect 339132 397724 339184 397730
rect 339132 397666 339184 397672
rect 339040 396432 339092 396438
rect 339040 396374 339092 396380
rect 339052 308582 339080 396374
rect 339144 311234 339172 397666
rect 339236 315353 339264 397831
rect 339328 368558 339356 450026
rect 339406 449712 339462 449721
rect 339406 449647 339462 449656
rect 339420 368665 339448 449647
rect 340156 407794 340184 451998
rect 340328 451308 340380 451314
rect 340328 451250 340380 451256
rect 340234 448624 340290 448633
rect 340234 448559 340290 448568
rect 340248 411262 340276 448559
rect 340340 424386 340368 451250
rect 340328 424380 340380 424386
rect 340328 424322 340380 424328
rect 340236 411256 340288 411262
rect 340236 411198 340288 411204
rect 340144 407788 340196 407794
rect 340144 407730 340196 407736
rect 340052 399220 340104 399226
rect 340052 399162 340104 399168
rect 339960 395208 340012 395214
rect 339960 395150 340012 395156
rect 339972 385966 340000 395150
rect 339960 385960 340012 385966
rect 339960 385902 340012 385908
rect 339406 368656 339462 368665
rect 339406 368591 339462 368600
rect 339316 368552 339368 368558
rect 339316 368494 339368 368500
rect 339316 323672 339368 323678
rect 339316 323614 339368 323620
rect 339328 320249 339356 323614
rect 339960 322312 340012 322318
rect 339960 322254 340012 322260
rect 339972 321881 340000 322254
rect 339498 321872 339554 321881
rect 339498 321807 339554 321816
rect 339958 321872 340014 321881
rect 339958 321807 340014 321816
rect 339314 320240 339370 320249
rect 339314 320175 339370 320184
rect 339222 315344 339278 315353
rect 339222 315279 339278 315288
rect 339132 311228 339184 311234
rect 339132 311170 339184 311176
rect 339040 308576 339092 308582
rect 339040 308518 339092 308524
rect 338948 306944 339000 306950
rect 338948 306886 339000 306892
rect 338856 298988 338908 298994
rect 338856 298930 338908 298936
rect 338396 238060 338448 238066
rect 338396 238002 338448 238008
rect 338304 231124 338356 231130
rect 338304 231066 338356 231072
rect 338212 226840 338264 226846
rect 338212 226782 338264 226788
rect 339512 221474 339540 321807
rect 340064 321201 340092 399162
rect 340420 396840 340472 396846
rect 340420 396782 340472 396788
rect 340236 396160 340288 396166
rect 340236 396102 340288 396108
rect 340144 389156 340196 389162
rect 340144 389098 340196 389104
rect 340050 321192 340106 321201
rect 340050 321127 340106 321136
rect 339590 316704 339646 316713
rect 339590 316639 339646 316648
rect 339604 226778 339632 316639
rect 340156 295186 340184 389098
rect 340248 305658 340276 396102
rect 340328 395820 340380 395826
rect 340328 395762 340380 395768
rect 340340 310962 340368 395762
rect 340432 313274 340460 396782
rect 340524 370054 340552 454038
rect 340696 452668 340748 452674
rect 340696 452610 340748 452616
rect 340604 394324 340656 394330
rect 340604 394266 340656 394272
rect 340512 370048 340564 370054
rect 340512 369990 340564 369996
rect 340510 334656 340566 334665
rect 340510 334591 340566 334600
rect 340524 316713 340552 334591
rect 340510 316704 340566 316713
rect 340510 316639 340566 316648
rect 340616 314634 340644 394266
rect 340708 373318 340736 452610
rect 340800 374678 340828 454174
rect 341524 454164 341576 454170
rect 341524 454106 341576 454112
rect 340878 451752 340934 451761
rect 340878 451687 340934 451696
rect 340892 443698 340920 451687
rect 340972 451580 341024 451586
rect 340972 451522 341024 451528
rect 340984 445058 341012 451522
rect 340972 445052 341024 445058
rect 340972 444994 341024 445000
rect 340880 443692 340932 443698
rect 340880 443634 340932 443640
rect 340970 438288 341026 438297
rect 340970 438223 341026 438232
rect 340984 438190 341012 438223
rect 340972 438184 341024 438190
rect 340972 438126 341024 438132
rect 340970 436792 341026 436801
rect 340970 436727 340972 436736
rect 341024 436727 341026 436736
rect 340972 436698 341024 436704
rect 340970 428496 341026 428505
rect 340970 428431 340972 428440
rect 341024 428431 341026 428440
rect 340972 428402 341024 428408
rect 341536 412634 341564 454106
rect 347778 452704 347834 452713
rect 347778 452639 347834 452648
rect 347412 452192 347464 452198
rect 347412 452134 347464 452140
rect 345570 451888 345626 451897
rect 341800 451852 341852 451858
rect 345570 451823 345626 451832
rect 341800 451794 341852 451800
rect 341616 451512 341668 451518
rect 341616 451454 341668 451460
rect 341444 412606 341564 412634
rect 340970 405784 341026 405793
rect 340970 405719 341026 405728
rect 340984 405686 341012 405719
rect 340972 405680 341024 405686
rect 340972 405622 341024 405628
rect 340878 399256 340934 399265
rect 340878 399191 340934 399200
rect 340892 398857 340920 399191
rect 340878 398848 340934 398857
rect 340878 398783 340934 398792
rect 341062 398848 341118 398857
rect 341444 398834 341472 412606
rect 341628 405793 341656 451454
rect 341708 449404 341760 449410
rect 341708 449346 341760 449352
rect 341720 428505 341748 449346
rect 341812 436801 341840 451794
rect 345202 451480 345258 451489
rect 342260 451444 342312 451450
rect 345202 451415 345258 451424
rect 342260 451386 342312 451392
rect 341892 451308 341944 451314
rect 341892 451250 341944 451256
rect 341904 438297 341932 451250
rect 342168 450016 342220 450022
rect 342168 449958 342220 449964
rect 341890 438288 341946 438297
rect 341890 438223 341946 438232
rect 341798 436792 341854 436801
rect 341798 436727 341854 436736
rect 341706 428496 341762 428505
rect 341706 428431 341762 428440
rect 341614 405784 341670 405793
rect 341614 405719 341670 405728
rect 342074 403064 342130 403073
rect 342074 402999 342130 403008
rect 341982 402112 342038 402121
rect 341982 402047 342038 402056
rect 341892 400988 341944 400994
rect 341892 400930 341944 400936
rect 341706 400752 341762 400761
rect 341706 400687 341762 400696
rect 341720 400654 341748 400687
rect 341708 400648 341760 400654
rect 341708 400590 341760 400596
rect 341800 400444 341852 400450
rect 341800 400386 341852 400392
rect 341614 400072 341670 400081
rect 341614 400007 341670 400016
rect 341444 398806 341564 398834
rect 341062 398783 341118 398792
rect 341076 398313 341104 398783
rect 341062 398304 341118 398313
rect 341062 398239 341118 398248
rect 341430 398304 341486 398313
rect 341430 398239 341486 398248
rect 341156 397384 341208 397390
rect 341156 397326 341208 397332
rect 341168 392630 341196 397326
rect 341340 395888 341392 395894
rect 341340 395830 341392 395836
rect 341156 392624 341208 392630
rect 341156 392566 341208 392572
rect 340788 374672 340840 374678
rect 340788 374614 340840 374620
rect 340696 373312 340748 373318
rect 340696 373254 340748 373260
rect 340880 369844 340932 369850
rect 340880 369786 340932 369792
rect 340892 369238 340920 369786
rect 340880 369232 340932 369238
rect 340880 369174 340932 369180
rect 340878 325000 340934 325009
rect 340878 324935 340934 324944
rect 340604 314628 340656 314634
rect 340604 314570 340656 314576
rect 340420 313268 340472 313274
rect 340420 313210 340472 313216
rect 340328 310956 340380 310962
rect 340328 310898 340380 310904
rect 340236 305652 340288 305658
rect 340236 305594 340288 305600
rect 340144 295180 340196 295186
rect 340144 295122 340196 295128
rect 339592 226772 339644 226778
rect 339592 226714 339644 226720
rect 340892 223553 340920 324935
rect 341352 316878 341380 395830
rect 341340 316872 341392 316878
rect 341340 316814 341392 316820
rect 341444 315994 341472 398239
rect 341536 370734 341564 398806
rect 341524 370728 341576 370734
rect 341524 370670 341576 370676
rect 341522 368656 341578 368665
rect 341522 368591 341578 368600
rect 341432 315988 341484 315994
rect 341432 315930 341484 315936
rect 340878 223544 340934 223553
rect 340878 223479 340934 223488
rect 339500 221468 339552 221474
rect 339500 221410 339552 221416
rect 335360 218748 335412 218754
rect 335360 218690 335412 218696
rect 336004 218748 336056 218754
rect 336004 218690 336056 218696
rect 334624 20664 334676 20670
rect 334624 20606 334676 20612
rect 335372 16574 335400 218690
rect 338120 137352 338172 137358
rect 338120 137294 338172 137300
rect 337384 124976 337436 124982
rect 337384 124918 337436 124924
rect 332612 16546 332732 16574
rect 335372 16546 336320 16574
rect 330390 6896 330446 6905
rect 330390 6831 330446 6840
rect 327816 4072 327868 4078
rect 327816 4014 327868 4020
rect 329288 4072 329340 4078
rect 329288 4014 329340 4020
rect 329300 3874 329328 4014
rect 327724 3868 327776 3874
rect 327724 3810 327776 3816
rect 329196 3868 329248 3874
rect 329196 3810 329248 3816
rect 329288 3868 329340 3874
rect 329288 3810 329340 3816
rect 327644 3454 328040 3482
rect 327540 3392 327592 3398
rect 327540 3334 327592 3340
rect 328012 480 328040 3454
rect 329208 480 329236 3810
rect 330404 480 330432 6831
rect 331588 4140 331640 4146
rect 331588 4082 331640 4088
rect 331600 480 331628 4082
rect 332704 480 332732 16546
rect 333886 6760 333942 6769
rect 333886 6695 333942 6704
rect 333900 480 333928 6695
rect 335084 3392 335136 3398
rect 335084 3334 335136 3340
rect 335096 480 335124 3334
rect 336292 480 336320 16546
rect 337396 4078 337424 124918
rect 338132 16574 338160 137294
rect 338132 16546 338712 16574
rect 337474 6624 337530 6633
rect 337474 6559 337530 6568
rect 337384 4072 337436 4078
rect 337384 4014 337436 4020
rect 337488 480 337516 6559
rect 338684 480 338712 16546
rect 326774 354 326886 480
rect 326356 326 326886 354
rect 326774 -960 326886 326
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339512 354 339540 221410
rect 340880 167068 340932 167074
rect 340880 167010 340932 167016
rect 340892 3210 340920 167010
rect 341536 100706 341564 368591
rect 341628 304570 341656 400007
rect 341812 399430 341840 400386
rect 341904 399566 341932 400930
rect 341996 399566 342024 402047
rect 342088 400110 342116 402999
rect 342076 400104 342128 400110
rect 342076 400046 342128 400052
rect 342076 399628 342128 399634
rect 342076 399570 342128 399576
rect 341892 399560 341944 399566
rect 341892 399502 341944 399508
rect 341984 399560 342036 399566
rect 341984 399502 342036 399508
rect 341800 399424 341852 399430
rect 342088 399401 342116 399570
rect 341800 399366 341852 399372
rect 342074 399392 342130 399401
rect 342074 399327 342130 399336
rect 342076 398336 342128 398342
rect 342076 398278 342128 398284
rect 341892 398132 341944 398138
rect 341892 398074 341944 398080
rect 341708 396636 341760 396642
rect 341708 396578 341760 396584
rect 341616 304564 341668 304570
rect 341616 304506 341668 304512
rect 341720 302870 341748 396578
rect 341800 395956 341852 395962
rect 341800 395898 341852 395904
rect 341708 302864 341760 302870
rect 341708 302806 341760 302812
rect 341812 300490 341840 395898
rect 341904 307222 341932 398074
rect 341984 396704 342036 396710
rect 341984 396646 342036 396652
rect 341996 309806 342024 396646
rect 342088 312798 342116 398278
rect 342180 369238 342208 449958
rect 342272 447134 342300 451386
rect 345216 449970 345244 451415
rect 345584 449970 345612 451823
rect 345938 451616 345994 451625
rect 345938 451551 345994 451560
rect 345952 449970 345980 451551
rect 347424 449970 347452 452134
rect 347792 449970 347820 452639
rect 348148 451376 348200 451382
rect 348148 451318 348200 451324
rect 348160 449970 348188 451318
rect 349252 451308 349304 451314
rect 349252 451250 349304 451256
rect 349264 449970 349292 451250
rect 350000 449970 350028 454514
rect 350540 451920 350592 451926
rect 350540 451862 350592 451868
rect 350552 450242 350580 451862
rect 350552 450214 350626 450242
rect 345216 449942 345460 449970
rect 345584 449942 345828 449970
rect 345952 449942 346196 449970
rect 347424 449942 347668 449970
rect 347792 449942 348036 449970
rect 348160 449942 348404 449970
rect 349264 449942 349508 449970
rect 350000 449942 350244 449970
rect 350598 449956 350626 450214
rect 350736 449970 350764 454922
rect 352104 454844 352156 454850
rect 352104 454786 352156 454792
rect 351460 451784 351512 451790
rect 351460 451726 351512 451732
rect 351092 450016 351144 450022
rect 350736 449942 350980 449970
rect 351472 449970 351500 451726
rect 352116 449970 352144 454786
rect 353668 452124 353720 452130
rect 353668 452066 353720 452072
rect 352564 451716 352616 451722
rect 352564 451658 352616 451664
rect 352196 451376 352248 451382
rect 352196 451318 352248 451324
rect 351144 449964 351348 449970
rect 351092 449958 351348 449964
rect 351104 449942 351348 449958
rect 351472 449942 351716 449970
rect 352084 449942 352144 449970
rect 352208 449970 352236 451318
rect 352576 449970 352604 451658
rect 352930 451344 352986 451353
rect 352930 451279 352986 451288
rect 352944 449970 352972 451279
rect 353300 450696 353352 450702
rect 353300 450638 353352 450644
rect 353312 450022 353340 450638
rect 353300 450016 353352 450022
rect 352208 449942 352452 449970
rect 352576 449942 352820 449970
rect 352944 449942 353188 449970
rect 353300 449958 353352 449964
rect 353680 449970 353708 452066
rect 354864 451988 354916 451994
rect 354864 451930 354916 451936
rect 354128 450016 354180 450022
rect 353680 449942 353924 449970
rect 354876 449970 354904 451930
rect 355232 450696 355284 450702
rect 355232 450638 355284 450644
rect 355244 449970 355272 450638
rect 355336 450430 355364 484366
rect 356704 472660 356756 472666
rect 356704 472602 356756 472608
rect 356244 463004 356296 463010
rect 356244 462946 356296 462952
rect 355968 456816 356020 456822
rect 355968 456758 356020 456764
rect 355980 453558 356008 456758
rect 355416 453552 355468 453558
rect 355416 453494 355468 453500
rect 355968 453552 356020 453558
rect 355968 453494 356020 453500
rect 355324 450424 355376 450430
rect 355324 450366 355376 450372
rect 355428 449970 355456 453494
rect 356060 453280 356112 453286
rect 356060 453222 356112 453228
rect 355508 450424 355560 450430
rect 355508 450366 355560 450372
rect 354180 449964 354292 449970
rect 354128 449958 354292 449964
rect 354140 449942 354292 449958
rect 354660 449954 354812 449970
rect 354660 449948 354824 449954
rect 354660 449942 354772 449948
rect 354876 449942 355272 449970
rect 355396 449942 355456 449970
rect 355520 449970 355548 450366
rect 356072 450242 356100 453222
rect 356256 450906 356284 462946
rect 356716 455598 356744 472602
rect 358084 468512 358136 468518
rect 358084 468454 358136 468460
rect 357256 460284 357308 460290
rect 357256 460226 357308 460232
rect 356704 455592 356756 455598
rect 356704 455534 356756 455540
rect 356980 455592 357032 455598
rect 356980 455534 357032 455540
rect 356336 452668 356388 452674
rect 356336 452610 356388 452616
rect 356244 450900 356296 450906
rect 356244 450842 356296 450848
rect 356256 450566 356284 450842
rect 356244 450560 356296 450566
rect 356244 450502 356296 450508
rect 356072 450214 356146 450242
rect 355520 449942 355764 449970
rect 356118 449956 356146 450214
rect 356348 449970 356376 452610
rect 356704 450696 356756 450702
rect 356704 450638 356756 450644
rect 356716 450566 356744 450638
rect 356612 450560 356664 450566
rect 356612 450502 356664 450508
rect 356704 450560 356756 450566
rect 356704 450502 356756 450508
rect 356624 449970 356652 450502
rect 356992 449970 357020 455534
rect 357268 453286 357296 460226
rect 357624 454232 357676 454238
rect 357624 454174 357676 454180
rect 357348 453348 357400 453354
rect 357348 453290 357400 453296
rect 357256 453280 357308 453286
rect 357256 453222 357308 453228
rect 357360 452674 357388 453290
rect 357348 452668 357400 452674
rect 357348 452610 357400 452616
rect 357636 449970 357664 454174
rect 358096 453626 358124 468454
rect 358084 453620 358136 453626
rect 358084 453562 358136 453568
rect 358096 449970 358124 453562
rect 356348 449942 356500 449970
rect 356624 449942 356868 449970
rect 356992 449942 357236 449970
rect 357604 449942 357664 449970
rect 357972 449942 358124 449970
rect 354772 449890 354824 449896
rect 347272 449712 347328 449721
rect 347272 449647 347328 449656
rect 346536 449576 346592 449585
rect 342352 449540 342404 449546
rect 349632 449546 349876 449562
rect 346536 449511 346592 449520
rect 349620 449540 349876 449546
rect 342352 449482 342404 449488
rect 349672 449534 349876 449540
rect 349620 449482 349672 449488
rect 342364 448594 342392 449482
rect 344466 449440 344522 449449
rect 344112 449410 344356 449426
rect 344100 449404 344356 449410
rect 344152 449398 344356 449404
rect 345202 449440 345258 449449
rect 344522 449398 344724 449426
rect 345092 449398 345202 449426
rect 344466 449375 344522 449384
rect 349342 449440 349398 449449
rect 348528 449410 348772 449426
rect 345202 449375 345258 449384
rect 348516 449404 348772 449410
rect 344100 449346 344152 449352
rect 348568 449398 348772 449404
rect 349140 449398 349342 449426
rect 349342 449375 349398 449384
rect 353390 449440 353446 449449
rect 358082 449440 358138 449449
rect 353446 449398 353556 449426
rect 353390 449375 353446 449384
rect 358464 449426 358492 576846
rect 358636 456136 358688 456142
rect 358636 456078 358688 456084
rect 358648 451625 358676 456078
rect 359188 455932 359240 455938
rect 359188 455874 359240 455880
rect 359200 455462 359228 455874
rect 359188 455456 359240 455462
rect 359188 455398 359240 455404
rect 358728 454844 358780 454850
rect 358728 454786 358780 454792
rect 358740 454238 358768 454786
rect 358728 454232 358780 454238
rect 358728 454174 358780 454180
rect 359096 454028 359148 454034
rect 359096 453970 359148 453976
rect 359108 453490 359136 453970
rect 359096 453484 359148 453490
rect 359096 453426 359148 453432
rect 358634 451616 358690 451625
rect 358634 451551 358690 451560
rect 358544 451308 358596 451314
rect 358544 451250 358596 451256
rect 358556 449478 358584 451250
rect 358648 450242 358676 451551
rect 358648 450214 358722 450242
rect 358694 449956 358722 450214
rect 359108 449970 359136 453426
rect 359076 449942 359136 449970
rect 359200 449970 359228 455398
rect 359476 453914 359504 670686
rect 359556 643136 359608 643142
rect 359556 643078 359608 643084
rect 359568 454034 359596 643078
rect 359648 630692 359700 630698
rect 359648 630634 359700 630640
rect 359660 455938 359688 630634
rect 360844 511284 360896 511290
rect 360844 511226 360896 511232
rect 360856 460934 360884 511226
rect 360936 469872 360988 469878
rect 360936 469814 360988 469820
rect 360488 460906 360884 460934
rect 359648 455932 359700 455938
rect 359648 455874 359700 455880
rect 360488 455802 360516 460906
rect 360660 458856 360712 458862
rect 360660 458798 360712 458804
rect 360476 455796 360528 455802
rect 360476 455738 360528 455744
rect 359556 454028 359608 454034
rect 359556 453970 359608 453976
rect 359476 453886 359596 453914
rect 359568 451353 359596 453886
rect 360384 453484 360436 453490
rect 360384 453426 360436 453432
rect 359554 451344 359610 451353
rect 359554 451279 359610 451288
rect 359568 449970 359596 451279
rect 360152 449984 360208 449993
rect 359200 449942 359444 449970
rect 359568 449942 359812 449970
rect 360396 449970 360424 453426
rect 360488 450242 360516 455738
rect 360672 454714 360700 458798
rect 360660 454708 360712 454714
rect 360660 454650 360712 454656
rect 360488 450214 360562 450242
rect 360208 449942 360424 449970
rect 360534 449956 360562 450214
rect 360672 449970 360700 454650
rect 360948 454170 360976 469814
rect 362316 465724 362368 465730
rect 362316 465666 362368 465672
rect 362224 464364 362276 464370
rect 362224 464306 362276 464312
rect 361580 454708 361632 454714
rect 361580 454650 361632 454656
rect 360936 454164 360988 454170
rect 360936 454106 360988 454112
rect 360948 451274 360976 454106
rect 361592 454102 361620 454650
rect 361580 454096 361632 454102
rect 361580 454038 361632 454044
rect 361592 453370 361620 454038
rect 361592 453342 361804 453370
rect 361670 452568 361726 452577
rect 361670 452503 361726 452512
rect 361684 452169 361712 452503
rect 361670 452160 361726 452169
rect 361670 452095 361726 452104
rect 360948 451246 361068 451274
rect 361040 449970 361068 451246
rect 361684 449970 361712 452095
rect 360672 449942 360916 449970
rect 361040 449942 361284 449970
rect 361652 449942 361712 449970
rect 361776 449970 361804 453342
rect 362236 452577 362264 464306
rect 362328 460934 362356 465666
rect 363052 461644 363104 461650
rect 363052 461586 363104 461592
rect 363064 460934 363092 461586
rect 362328 460906 362540 460934
rect 363064 460906 363368 460934
rect 362316 456068 362368 456074
rect 362316 456010 362368 456016
rect 362222 452568 362278 452577
rect 362222 452503 362278 452512
rect 362224 451376 362276 451382
rect 362224 451318 362276 451324
rect 361776 449942 362020 449970
rect 360152 449919 360208 449928
rect 358138 449398 358492 449426
rect 358544 449472 358596 449478
rect 358544 449414 358596 449420
rect 362236 449410 362264 451318
rect 362328 450770 362356 456010
rect 362512 455734 362540 460906
rect 363236 460216 363288 460222
rect 363236 460158 363288 460164
rect 362500 455728 362552 455734
rect 362500 455670 362552 455676
rect 362316 450764 362368 450770
rect 362316 450706 362368 450712
rect 362328 450242 362356 450706
rect 362328 450214 362402 450242
rect 362374 449956 362402 450214
rect 362512 449970 362540 455670
rect 363248 454782 363276 460158
rect 363236 454776 363288 454782
rect 363236 454718 363288 454724
rect 363248 449970 363276 454718
rect 363340 454646 363368 460906
rect 363512 455932 363564 455938
rect 363512 455874 363564 455880
rect 363524 455666 363552 455874
rect 363512 455660 363564 455666
rect 363512 455602 363564 455608
rect 363328 454640 363380 454646
rect 363328 454582 363380 454588
rect 362512 449942 362756 449970
rect 363124 449942 363276 449970
rect 363340 449970 363368 454582
rect 363524 451274 363552 455602
rect 363616 454458 363644 698634
rect 363696 474020 363748 474026
rect 363696 473962 363748 473968
rect 363708 455938 363736 473962
rect 363696 455932 363748 455938
rect 363696 455874 363748 455880
rect 364352 455530 364380 700334
rect 364432 700324 364484 700330
rect 364432 700266 364484 700272
rect 364444 455870 364472 700266
rect 364996 698698 365024 703520
rect 397472 699718 397500 703520
rect 396724 699712 396776 699718
rect 396724 699654 396776 699660
rect 397460 699712 397512 699718
rect 397460 699654 397512 699660
rect 364984 698692 365036 698698
rect 364984 698634 365036 698640
rect 378784 696992 378836 696998
rect 378784 696934 378836 696940
rect 369860 683188 369912 683194
rect 369860 683130 369912 683136
rect 367744 590708 367796 590714
rect 367744 590650 367796 590656
rect 367756 468518 367784 590650
rect 367836 470620 367888 470626
rect 367836 470562 367888 470568
rect 367744 468512 367796 468518
rect 367744 468454 367796 468460
rect 367100 463752 367152 463758
rect 367100 463694 367152 463700
rect 365812 460964 365864 460970
rect 367112 460934 367140 463694
rect 365864 460912 366220 460934
rect 365812 460906 366220 460912
rect 367112 460906 367324 460934
rect 364432 455864 364484 455870
rect 364432 455806 364484 455812
rect 364340 455524 364392 455530
rect 364340 455466 364392 455472
rect 363616 454430 364012 454458
rect 363984 451314 364012 454430
rect 363972 451308 364024 451314
rect 363524 451246 363644 451274
rect 363972 451250 364024 451256
rect 363616 449970 363644 451246
rect 363984 449970 364012 451250
rect 364444 449970 364472 455806
rect 364708 455524 364760 455530
rect 364708 455466 364760 455472
rect 364720 449970 364748 455466
rect 365812 451444 365864 451450
rect 365812 451386 365864 451392
rect 365720 450832 365772 450838
rect 365720 450774 365772 450780
rect 365732 449970 365760 450774
rect 363340 449942 363492 449970
rect 363616 449942 363860 449970
rect 363984 449942 364228 449970
rect 364444 449942 364596 449970
rect 364720 449942 364964 449970
rect 365700 449942 365760 449970
rect 365824 449970 365852 451386
rect 366192 449970 366220 460906
rect 367192 454912 367244 454918
rect 367192 454854 367244 454860
rect 366548 450084 366600 450090
rect 366548 450026 366600 450032
rect 366560 449970 366588 450026
rect 367204 449970 367232 454854
rect 365824 449942 366068 449970
rect 366192 449942 366436 449970
rect 366560 449942 366804 449970
rect 367172 449942 367232 449970
rect 367296 449970 367324 460906
rect 367848 460290 367876 470562
rect 368572 467152 368624 467158
rect 368572 467094 368624 467100
rect 367836 460284 367888 460290
rect 367836 460226 367888 460232
rect 368018 452840 368074 452849
rect 368018 452775 368074 452784
rect 367652 450492 367704 450498
rect 367652 450434 367704 450440
rect 367664 449970 367692 450434
rect 368032 449970 368060 452775
rect 368584 452577 368612 467094
rect 368664 465112 368716 465118
rect 368664 465054 368716 465060
rect 368570 452568 368626 452577
rect 368570 452503 368626 452512
rect 368584 451489 368612 452503
rect 368570 451480 368626 451489
rect 368570 451415 368626 451424
rect 368676 449970 368704 465054
rect 369490 452568 369546 452577
rect 369490 452503 369546 452512
rect 369124 451376 369176 451382
rect 369124 451318 369176 451324
rect 367296 449942 367540 449970
rect 367664 449942 367908 449970
rect 368032 449942 368276 449970
rect 368644 449942 368704 449970
rect 369136 449970 369164 451318
rect 369504 449970 369532 452503
rect 369136 449942 369380 449970
rect 369504 449942 369748 449970
rect 369872 449478 369900 683130
rect 371424 632120 371476 632126
rect 371424 632062 371476 632068
rect 371436 460934 371464 632062
rect 372620 579692 372672 579698
rect 372620 579634 372672 579640
rect 371436 460906 371740 460934
rect 371330 454200 371386 454209
rect 371330 454135 371386 454144
rect 371240 453212 371292 453218
rect 371240 453154 371292 453160
rect 369952 453144 370004 453150
rect 369952 453086 370004 453092
rect 369964 451314 369992 453086
rect 371252 451926 371280 453154
rect 371240 451920 371292 451926
rect 371240 451862 371292 451868
rect 370228 451648 370280 451654
rect 370228 451590 370280 451596
rect 369952 451308 370004 451314
rect 369952 451250 370004 451256
rect 370088 450256 370144 450265
rect 370088 450191 370144 450200
rect 370102 449956 370130 450191
rect 370240 449970 370268 451590
rect 371344 449970 371372 454135
rect 371422 451752 371478 451761
rect 371422 451687 371478 451696
rect 370240 449942 370484 449970
rect 371220 449942 371372 449970
rect 371436 449970 371464 451687
rect 371436 449942 371588 449970
rect 371712 449562 371740 460906
rect 372632 452577 372660 579634
rect 376024 563100 376076 563106
rect 376024 563042 376076 563048
rect 374000 527196 374052 527202
rect 374000 527138 374052 527144
rect 373540 457156 373592 457162
rect 373540 457098 373592 457104
rect 372802 454064 372858 454073
rect 372802 453999 372858 454008
rect 372618 452568 372674 452577
rect 372618 452503 372674 452512
rect 372816 449970 372844 453999
rect 373400 450120 373456 450129
rect 373400 450055 373456 450064
rect 372692 449942 372844 449970
rect 373414 449956 373442 450055
rect 373552 449970 373580 457098
rect 374012 451489 374040 527138
rect 374092 474768 374144 474774
rect 374092 474710 374144 474716
rect 374104 452577 374132 474710
rect 375748 457088 375800 457094
rect 375748 457030 375800 457036
rect 374090 452568 374146 452577
rect 374090 452503 374146 452512
rect 373998 451480 374054 451489
rect 373998 451415 374054 451424
rect 374012 449970 374040 451415
rect 375380 451308 375432 451314
rect 375380 451250 375432 451256
rect 374506 450152 374558 450158
rect 374506 450094 374558 450100
rect 373552 449942 373796 449970
rect 374012 449942 374164 449970
rect 374518 449956 374546 450094
rect 375392 449970 375420 451250
rect 375760 449970 375788 457030
rect 376036 454850 376064 563042
rect 377404 536852 377456 536858
rect 377404 536794 377456 536800
rect 377416 463010 377444 536794
rect 377404 463004 377456 463010
rect 377404 462946 377456 462952
rect 378232 456952 378284 456958
rect 378232 456894 378284 456900
rect 376024 454844 376076 454850
rect 376024 454786 376076 454792
rect 377588 454504 377640 454510
rect 377588 454446 377640 454452
rect 376944 454368 376996 454374
rect 376944 454310 376996 454316
rect 376116 452940 376168 452946
rect 376116 452882 376168 452888
rect 376128 449970 376156 452882
rect 376760 452736 376812 452742
rect 376760 452678 376812 452684
rect 376772 449970 376800 452678
rect 375392 449942 375636 449970
rect 375760 449942 376004 449970
rect 376128 449942 376372 449970
rect 376740 449942 376800 449970
rect 376956 449970 376984 454310
rect 377220 452872 377272 452878
rect 377220 452814 377272 452820
rect 377232 449970 377260 452814
rect 377600 449970 377628 454446
rect 378244 449970 378272 456894
rect 378796 453490 378824 696934
rect 382924 616888 382976 616894
rect 382924 616830 382976 616836
rect 380164 457020 380216 457026
rect 380164 456962 380216 456968
rect 379796 454300 379848 454306
rect 379796 454242 379848 454248
rect 378784 453484 378836 453490
rect 378784 453426 378836 453432
rect 379060 451852 379112 451858
rect 379060 451794 379112 451800
rect 378690 451344 378746 451353
rect 378690 451279 378746 451288
rect 378324 450288 378376 450294
rect 378324 450230 378376 450236
rect 376956 449942 377108 449970
rect 377232 449942 377476 449970
rect 377600 449942 377844 449970
rect 378212 449942 378272 449970
rect 378336 449970 378364 450230
rect 378704 449970 378732 451279
rect 379072 449970 379100 451794
rect 379658 450220 379710 450226
rect 379658 450162 379710 450168
rect 378336 449942 378580 449970
rect 378704 449942 378948 449970
rect 379072 449942 379316 449970
rect 379670 449956 379698 450162
rect 379808 449970 379836 454242
rect 380176 449970 380204 456962
rect 381268 456884 381320 456890
rect 381268 456826 381320 456832
rect 380532 450628 380584 450634
rect 380532 450570 380584 450576
rect 380544 449970 380572 450570
rect 380900 450356 380952 450362
rect 380900 450298 380952 450304
rect 380912 449970 380940 450298
rect 381280 449970 381308 456826
rect 382936 456142 382964 616830
rect 392584 524476 392636 524482
rect 392584 524418 392636 524424
rect 392596 472666 392624 524418
rect 392584 472660 392636 472666
rect 392584 472602 392636 472608
rect 396736 461650 396764 699654
rect 412652 474026 412680 703582
rect 413480 703474 413508 703582
rect 413622 703520 413734 704960
rect 429212 703582 429700 703610
rect 413664 703474 413692 703520
rect 413480 703446 413692 703474
rect 412640 474020 412692 474026
rect 412640 473962 412692 473968
rect 396724 461644 396776 461650
rect 396724 461586 396776 461592
rect 429212 460222 429240 703582
rect 429672 703474 429700 703582
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 429856 703474 429884 703520
rect 429672 703446 429884 703474
rect 429200 460216 429252 460222
rect 429200 460158 429252 460164
rect 382924 456136 382976 456142
rect 382924 456078 382976 456084
rect 462332 456074 462360 703520
rect 478524 702434 478552 703520
rect 477512 702406 478552 702434
rect 477512 465730 477540 702406
rect 477500 465724 477552 465730
rect 477500 465666 477552 465672
rect 462320 456068 462372 456074
rect 462320 456010 462372 456016
rect 494072 454714 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 527192 469878 527220 703520
rect 543476 702434 543504 703520
rect 559668 702434 559696 703520
rect 542372 702406 543504 702434
rect 558932 702406 559696 702434
rect 527180 469872 527232 469878
rect 527180 469814 527232 469820
rect 542372 464370 542400 702406
rect 542360 464364 542412 464370
rect 542360 464306 542412 464312
rect 558932 458862 558960 702406
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580262 683904 580318 683913
rect 580262 683839 580318 683848
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 579986 630864 580042 630873
rect 579986 630799 580042 630808
rect 580000 630698 580028 630799
rect 579988 630692 580040 630698
rect 579988 630634 580040 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 580170 591016 580226 591025
rect 580170 590951 580226 590960
rect 580184 590714 580212 590951
rect 580172 590708 580224 590714
rect 580172 590650 580224 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 580170 564360 580226 564369
rect 580170 564295 580226 564304
rect 580184 563106 580212 564295
rect 580172 563100 580224 563106
rect 580172 563042 580224 563048
rect 579894 537840 579950 537849
rect 579894 537775 579950 537784
rect 579908 536858 579936 537775
rect 579896 536852 579948 536858
rect 579896 536794 579948 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580276 511290 580304 683839
rect 580354 511320 580410 511329
rect 580264 511284 580316 511290
rect 580354 511255 580410 511264
rect 580264 511226 580316 511232
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 580078 471472 580134 471481
rect 580078 471407 580134 471416
rect 580092 470626 580120 471407
rect 580080 470620 580132 470626
rect 580080 470562 580132 470568
rect 558920 458856 558972 458862
rect 558920 458798 558972 458804
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 494060 454708 494112 454714
rect 494060 454650 494112 454656
rect 382464 454436 382516 454442
rect 382464 454378 382516 454384
rect 381636 453008 381688 453014
rect 381636 452950 381688 452956
rect 381648 449970 381676 452950
rect 382476 449970 382504 454378
rect 580368 453354 580396 511255
rect 580356 453348 580408 453354
rect 580356 453290 580408 453296
rect 382740 453076 382792 453082
rect 382740 453018 382792 453024
rect 382556 451580 382608 451586
rect 382556 451522 382608 451528
rect 382568 450242 382596 451522
rect 382568 450214 382642 450242
rect 379808 449942 380052 449970
rect 380176 449942 380420 449970
rect 380544 449942 380788 449970
rect 380912 449942 381156 449970
rect 381280 449942 381524 449970
rect 381648 449942 381892 449970
rect 382260 449942 382504 449970
rect 382614 449956 382642 450214
rect 382752 449970 382780 453018
rect 383844 452804 383896 452810
rect 383844 452746 383896 452752
rect 383856 449970 383884 452746
rect 384580 452056 384632 452062
rect 384580 451998 384632 452004
rect 384592 449970 384620 451998
rect 385040 451920 385092 451926
rect 385040 451862 385092 451868
rect 385052 449970 385080 451862
rect 580264 450560 580316 450566
rect 580264 450502 580316 450508
rect 388444 450016 388496 450022
rect 382752 449942 382996 449970
rect 383856 449942 384100 449970
rect 384592 449942 384836 449970
rect 385052 449942 385204 449970
rect 388444 449958 388496 449964
rect 371928 449576 371984 449585
rect 371712 449534 371928 449562
rect 371928 449511 371984 449520
rect 370608 449478 370636 449509
rect 365076 449472 365128 449478
rect 369860 449472 369912 449478
rect 365128 449420 365332 449426
rect 365076 449414 365332 449420
rect 370596 449472 370648 449478
rect 369860 449414 369912 449420
rect 370594 449440 370596 449449
rect 370648 449440 370650 449449
rect 372066 449440 372122 449449
rect 362224 449404 362276 449410
rect 358082 449375 358138 449384
rect 348516 449346 348568 449352
rect 365088 449398 365332 449414
rect 370650 449398 370852 449426
rect 370594 449375 370650 449384
rect 372802 449440 372858 449449
rect 372122 449398 372324 449426
rect 372066 449375 372122 449384
rect 375010 449440 375066 449449
rect 372858 449398 373060 449426
rect 372802 449375 372858 449384
rect 383106 449440 383162 449449
rect 375066 449398 375268 449426
rect 375010 449375 375066 449384
rect 383842 449440 383898 449449
rect 383162 449398 383364 449426
rect 383732 449398 383842 449426
rect 383106 449375 383162 449384
rect 383842 449375 383898 449384
rect 384302 449440 384358 449449
rect 385682 449440 385738 449449
rect 384358 449398 384468 449426
rect 384302 449375 384358 449384
rect 385738 449398 385940 449426
rect 385682 449375 385738 449384
rect 362224 449346 362276 449352
rect 342444 449336 342496 449342
rect 342444 449278 342496 449284
rect 343960 449304 344016 449313
rect 342456 448662 342484 449278
rect 343960 449239 344016 449248
rect 346904 449304 346960 449313
rect 346904 449239 346960 449248
rect 368984 449304 369040 449313
rect 368984 449239 369040 449248
rect 374872 449304 374928 449313
rect 374872 449239 374928 449248
rect 385544 449304 385600 449313
rect 385544 449239 385600 449248
rect 342444 448656 342496 448662
rect 342444 448598 342496 448604
rect 342352 448588 342404 448594
rect 342352 448530 342404 448536
rect 342272 447106 342484 447134
rect 342456 439521 342484 447106
rect 342442 439512 342498 439521
rect 342442 439447 342498 439456
rect 388456 422294 388484 449958
rect 389824 449948 389876 449954
rect 389824 449890 389876 449896
rect 389836 431934 389864 449890
rect 389824 431928 389876 431934
rect 389824 431870 389876 431876
rect 580172 431928 580224 431934
rect 580172 431870 580224 431876
rect 580184 431633 580212 431870
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 388456 422266 389036 422294
rect 389008 405686 389036 422266
rect 580276 418305 580304 450502
rect 580262 418296 580318 418305
rect 580262 418231 580318 418240
rect 388996 405680 389048 405686
rect 388996 405622 389048 405628
rect 580172 405680 580224 405686
rect 580172 405622 580224 405628
rect 580184 404977 580212 405622
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580722 400888 580778 400897
rect 580722 400823 580778 400832
rect 342260 400444 342312 400450
rect 342260 400386 342312 400392
rect 342272 400246 342300 400386
rect 387524 400376 387576 400382
rect 387524 400318 387576 400324
rect 342260 400240 342312 400246
rect 342260 400182 342312 400188
rect 342260 400104 342312 400110
rect 342260 400046 342312 400052
rect 342272 399634 342300 400046
rect 342502 399956 342530 400044
rect 342364 399928 342530 399956
rect 342364 399752 342392 399928
rect 342594 399888 342622 400044
rect 342548 399860 342622 399888
rect 342364 399724 342484 399752
rect 342260 399628 342312 399634
rect 342260 399570 342312 399576
rect 342260 399424 342312 399430
rect 342260 399366 342312 399372
rect 342272 395457 342300 399366
rect 342258 395448 342314 395457
rect 342258 395383 342314 395392
rect 342456 389910 342484 399724
rect 342548 398206 342576 399860
rect 342686 399752 342714 400044
rect 342640 399724 342714 399752
rect 342778 399752 342806 400044
rect 342870 399906 342898 400044
rect 342858 399900 342910 399906
rect 342858 399842 342910 399848
rect 342962 399838 342990 400044
rect 343054 399906 343082 400044
rect 343042 399900 343094 399906
rect 343042 399842 343094 399848
rect 342950 399832 343002 399838
rect 343146 399786 343174 400044
rect 342950 399774 343002 399780
rect 343054 399758 343174 399786
rect 342778 399724 342852 399752
rect 342536 398200 342588 398206
rect 342536 398142 342588 398148
rect 342640 396074 342668 399724
rect 342720 398200 342772 398206
rect 342824 398177 342852 399724
rect 343054 399684 343082 399758
rect 343238 399684 343266 400044
rect 343330 399906 343358 400044
rect 343318 399900 343370 399906
rect 343318 399842 343370 399848
rect 343422 399786 343450 400044
rect 343514 399838 343542 400044
rect 343008 399656 343082 399684
rect 343192 399656 343266 399684
rect 343376 399758 343450 399786
rect 343502 399832 343554 399838
rect 343502 399774 343554 399780
rect 342720 398142 342772 398148
rect 342810 398168 342866 398177
rect 342548 396046 342668 396074
rect 342548 396012 342576 396046
rect 342548 395984 342668 396012
rect 342536 394596 342588 394602
rect 342536 394538 342588 394544
rect 342444 389904 342496 389910
rect 342444 389846 342496 389852
rect 342258 389192 342314 389201
rect 342258 389127 342314 389136
rect 342272 388618 342300 389127
rect 342548 388754 342576 394538
rect 342536 388748 342588 388754
rect 342536 388690 342588 388696
rect 342260 388612 342312 388618
rect 342260 388554 342312 388560
rect 342640 377466 342668 395984
rect 342732 380254 342760 398142
rect 342810 398103 342866 398112
rect 342904 394868 342956 394874
rect 342904 394810 342956 394816
rect 342720 380248 342772 380254
rect 342720 380190 342772 380196
rect 342628 377460 342680 377466
rect 342628 377402 342680 377408
rect 342168 369232 342220 369238
rect 342168 369174 342220 369180
rect 342350 325272 342406 325281
rect 342350 325207 342406 325216
rect 342364 320346 342392 325207
rect 342352 320340 342404 320346
rect 342352 320282 342404 320288
rect 342076 312792 342128 312798
rect 342076 312734 342128 312740
rect 342260 311160 342312 311166
rect 342260 311102 342312 311108
rect 341984 309800 342036 309806
rect 341984 309742 342036 309748
rect 341892 307216 341944 307222
rect 341892 307158 341944 307164
rect 341800 300484 341852 300490
rect 341800 300426 341852 300432
rect 342272 203590 342300 311102
rect 342364 219337 342392 320282
rect 342916 295254 342944 394810
rect 343008 394602 343036 399656
rect 343088 397452 343140 397458
rect 343088 397394 343140 397400
rect 342996 394596 343048 394602
rect 342996 394538 343048 394544
rect 342996 393508 343048 393514
rect 342996 393450 343048 393456
rect 343008 297498 343036 393450
rect 343100 392086 343128 397394
rect 343192 393922 343220 399656
rect 343376 396817 343404 399758
rect 343502 399696 343554 399702
rect 343502 399638 343554 399644
rect 343606 399650 343634 400044
rect 343698 399770 343726 400044
rect 343790 399838 343818 400044
rect 343882 399906 343910 400044
rect 343974 399906 344002 400044
rect 343870 399900 343922 399906
rect 343870 399842 343922 399848
rect 343962 399900 344014 399906
rect 343962 399842 344014 399848
rect 344066 399838 344094 400044
rect 344158 399906 344186 400044
rect 344146 399900 344198 399906
rect 344146 399842 344198 399848
rect 343778 399832 343830 399838
rect 343778 399774 343830 399780
rect 344054 399832 344106 399838
rect 344250 399786 344278 400044
rect 344342 399906 344370 400044
rect 344330 399900 344382 399906
rect 344330 399842 344382 399848
rect 344054 399774 344106 399780
rect 343686 399764 343738 399770
rect 343962 399764 344014 399770
rect 343686 399706 343738 399712
rect 343882 399724 343962 399752
rect 343882 399650 343910 399724
rect 343962 399706 344014 399712
rect 344204 399758 344278 399786
rect 343514 398834 343542 399638
rect 343606 399622 343680 399650
rect 343514 398806 343588 398834
rect 343456 398744 343508 398750
rect 343456 398686 343508 398692
rect 343362 396808 343418 396817
rect 343362 396743 343418 396752
rect 343364 396568 343416 396574
rect 343364 396510 343416 396516
rect 343376 395486 343404 396510
rect 343364 395480 343416 395486
rect 343364 395422 343416 395428
rect 343468 394074 343496 398686
rect 343560 395962 343588 398806
rect 343652 398478 343680 399622
rect 343836 399622 343910 399650
rect 344008 399628 344060 399634
rect 343640 398472 343692 398478
rect 343640 398414 343692 398420
rect 343836 398410 343864 399622
rect 344008 399570 344060 399576
rect 344100 399628 344152 399634
rect 344100 399570 344152 399576
rect 343916 399560 343968 399566
rect 343916 399502 343968 399508
rect 343824 398404 343876 398410
rect 343824 398346 343876 398352
rect 343928 398002 343956 399502
rect 344020 399265 344048 399570
rect 344006 399256 344062 399265
rect 344006 399191 344062 399200
rect 344112 398290 344140 399570
rect 344020 398262 344140 398290
rect 343916 397996 343968 398002
rect 343916 397938 343968 397944
rect 343732 397860 343784 397866
rect 343732 397802 343784 397808
rect 343640 396500 343692 396506
rect 343640 396442 343692 396448
rect 343548 395956 343600 395962
rect 343548 395898 343600 395904
rect 343652 394369 343680 396442
rect 343638 394360 343694 394369
rect 343638 394295 343694 394304
rect 343376 394046 343496 394074
rect 343180 393916 343232 393922
rect 343180 393858 343232 393864
rect 343180 393100 343232 393106
rect 343180 393042 343232 393048
rect 343088 392080 343140 392086
rect 343088 392022 343140 392028
rect 343088 388748 343140 388754
rect 343088 388690 343140 388696
rect 343100 304434 343128 388690
rect 343192 308514 343220 393042
rect 343270 383480 343326 383489
rect 343270 383415 343326 383424
rect 343180 308508 343232 308514
rect 343180 308450 343232 308456
rect 343088 304428 343140 304434
rect 343088 304370 343140 304376
rect 343284 300286 343312 383415
rect 343376 319598 343404 394046
rect 343456 393916 343508 393922
rect 343456 393858 343508 393864
rect 343468 387433 343496 393858
rect 343744 391241 343772 397802
rect 343824 397588 343876 397594
rect 343824 397530 343876 397536
rect 343836 392562 343864 397530
rect 344020 397390 344048 398262
rect 344100 398200 344152 398206
rect 344100 398142 344152 398148
rect 344008 397384 344060 397390
rect 344008 397326 344060 397332
rect 343916 395412 343968 395418
rect 343916 395354 343968 395360
rect 343824 392556 343876 392562
rect 343824 392498 343876 392504
rect 343730 391232 343786 391241
rect 343730 391167 343786 391176
rect 343454 387424 343510 387433
rect 343454 387359 343510 387368
rect 343548 383512 343600 383518
rect 343548 383454 343600 383460
rect 343456 383444 343508 383450
rect 343456 383386 343508 383392
rect 343364 319592 343416 319598
rect 343364 319534 343416 319540
rect 343468 311166 343496 383386
rect 343560 312526 343588 383454
rect 343928 319258 343956 395354
rect 344112 392494 344140 398142
rect 344204 395865 344232 399758
rect 344434 399752 344462 400044
rect 344388 399724 344462 399752
rect 344284 399696 344336 399702
rect 344284 399638 344336 399644
rect 344296 398682 344324 399638
rect 344284 398676 344336 398682
rect 344284 398618 344336 398624
rect 344284 398336 344336 398342
rect 344284 398278 344336 398284
rect 344190 395856 344246 395865
rect 344190 395791 344246 395800
rect 344192 395616 344244 395622
rect 344192 395558 344244 395564
rect 344100 392488 344152 392494
rect 344100 392430 344152 392436
rect 344100 387184 344152 387190
rect 344100 387126 344152 387132
rect 343916 319252 343968 319258
rect 343916 319194 343968 319200
rect 344112 312905 344140 387126
rect 344204 387025 344232 395558
rect 344190 387016 344246 387025
rect 344190 386951 344246 386960
rect 344098 312896 344154 312905
rect 344098 312831 344154 312840
rect 343548 312520 343600 312526
rect 343548 312462 343600 312468
rect 343456 311160 343508 311166
rect 343456 311102 343508 311108
rect 343272 300280 343324 300286
rect 343272 300222 343324 300228
rect 342996 297492 343048 297498
rect 342996 297434 343048 297440
rect 342904 295248 342956 295254
rect 342904 295190 342956 295196
rect 344296 295118 344324 398278
rect 344388 395418 344416 399724
rect 344526 399650 344554 400044
rect 344618 399752 344646 400044
rect 344710 399906 344738 400044
rect 344698 399900 344750 399906
rect 344698 399842 344750 399848
rect 344802 399786 344830 400044
rect 344894 399906 344922 400044
rect 344882 399900 344934 399906
rect 344882 399842 344934 399848
rect 344756 399758 344830 399786
rect 344618 399724 344692 399752
rect 344480 399622 344554 399650
rect 344480 398993 344508 399622
rect 344560 399560 344612 399566
rect 344560 399502 344612 399508
rect 344572 399344 344600 399502
rect 344664 399480 344692 399724
rect 344756 399634 344784 399758
rect 344986 399752 345014 400044
rect 344940 399724 345014 399752
rect 344836 399696 344888 399702
rect 344836 399638 344888 399644
rect 344744 399628 344796 399634
rect 344744 399570 344796 399576
rect 344664 399452 344784 399480
rect 344572 399316 344692 399344
rect 344560 399220 344612 399226
rect 344560 399162 344612 399168
rect 344466 398984 344522 398993
rect 344466 398919 344522 398928
rect 344468 398676 344520 398682
rect 344468 398618 344520 398624
rect 344480 398546 344508 398618
rect 344468 398540 344520 398546
rect 344468 398482 344520 398488
rect 344572 398274 344600 399162
rect 344664 398993 344692 399316
rect 344650 398984 344706 398993
rect 344650 398919 344706 398928
rect 344652 398812 344704 398818
rect 344756 398800 344784 399452
rect 344704 398772 344784 398800
rect 344652 398754 344704 398760
rect 344560 398268 344612 398274
rect 344560 398210 344612 398216
rect 344376 395412 344428 395418
rect 344376 395354 344428 395360
rect 344652 393644 344704 393650
rect 344652 393586 344704 393592
rect 344664 392714 344692 393586
rect 344480 392686 344692 392714
rect 344376 390788 344428 390794
rect 344376 390730 344428 390736
rect 344388 301714 344416 390730
rect 344376 301708 344428 301714
rect 344376 301650 344428 301656
rect 344480 299062 344508 392686
rect 344560 392556 344612 392562
rect 344560 392498 344612 392504
rect 344572 307290 344600 392498
rect 344744 392488 344796 392494
rect 344744 392430 344796 392436
rect 344650 388240 344706 388249
rect 344650 388175 344706 388184
rect 344560 307284 344612 307290
rect 344560 307226 344612 307232
rect 344664 300218 344692 388175
rect 344756 310146 344784 392430
rect 344848 387394 344876 399638
rect 344940 392698 344968 399724
rect 345078 399650 345106 400044
rect 345170 399752 345198 400044
rect 345262 399906 345290 400044
rect 345250 399900 345302 399906
rect 345250 399842 345302 399848
rect 345354 399752 345382 400044
rect 345446 399786 345474 400044
rect 345538 399906 345566 400044
rect 345526 399900 345578 399906
rect 345526 399842 345578 399848
rect 345446 399758 345520 399786
rect 345170 399724 345244 399752
rect 345032 399622 345106 399650
rect 345032 396137 345060 399622
rect 345112 398744 345164 398750
rect 345112 398686 345164 398692
rect 345124 398138 345152 398686
rect 345112 398132 345164 398138
rect 345112 398074 345164 398080
rect 345018 396128 345074 396137
rect 345018 396063 345074 396072
rect 345216 395944 345244 399724
rect 345032 395916 345244 395944
rect 345308 399724 345382 399752
rect 345032 395622 345060 395916
rect 345308 395876 345336 399724
rect 345388 399628 345440 399634
rect 345388 399570 345440 399576
rect 345400 397372 345428 399570
rect 345492 398682 345520 399758
rect 345630 399752 345658 400044
rect 345722 399838 345750 400044
rect 345814 399906 345842 400044
rect 345802 399900 345854 399906
rect 345802 399842 345854 399848
rect 345710 399832 345762 399838
rect 345710 399774 345762 399780
rect 345906 399752 345934 400044
rect 345584 399724 345658 399752
rect 345860 399724 345934 399752
rect 345998 399752 346026 400044
rect 346090 399906 346118 400044
rect 346078 399900 346130 399906
rect 346078 399842 346130 399848
rect 346182 399838 346210 400044
rect 346274 399906 346302 400044
rect 346262 399900 346314 399906
rect 346262 399842 346314 399848
rect 346170 399832 346222 399838
rect 346170 399774 346222 399780
rect 346366 399752 346394 400044
rect 346458 399906 346486 400044
rect 346550 399906 346578 400044
rect 346446 399900 346498 399906
rect 346446 399842 346498 399848
rect 346538 399900 346590 399906
rect 346538 399842 346590 399848
rect 346492 399764 346544 399770
rect 345998 399724 346072 399752
rect 346366 399724 346440 399752
rect 345480 398676 345532 398682
rect 345480 398618 345532 398624
rect 345400 397344 345520 397372
rect 345124 395848 345336 395876
rect 345020 395616 345072 395622
rect 345020 395558 345072 395564
rect 344928 392692 344980 392698
rect 344928 392634 344980 392640
rect 345124 391105 345152 395848
rect 345296 395616 345348 395622
rect 345296 395558 345348 395564
rect 345204 395412 345256 395418
rect 345204 395354 345256 395360
rect 345110 391096 345166 391105
rect 345110 391031 345166 391040
rect 344928 388952 344980 388958
rect 344928 388894 344980 388900
rect 344836 387388 344888 387394
rect 344836 387330 344888 387336
rect 344940 315722 344968 388894
rect 345216 387258 345244 395354
rect 345308 388686 345336 395558
rect 345388 395004 345440 395010
rect 345388 394946 345440 394952
rect 345400 388929 345428 394946
rect 345386 388920 345442 388929
rect 345386 388855 345442 388864
rect 345296 388680 345348 388686
rect 345296 388622 345348 388628
rect 345204 387252 345256 387258
rect 345204 387194 345256 387200
rect 345492 320793 345520 397344
rect 345584 395622 345612 399724
rect 345756 399628 345808 399634
rect 345756 399570 345808 399576
rect 345664 399356 345716 399362
rect 345664 399298 345716 399304
rect 345676 399265 345704 399298
rect 345662 399256 345718 399265
rect 345662 399191 345718 399200
rect 345664 397928 345716 397934
rect 345664 397870 345716 397876
rect 345676 397730 345704 397870
rect 345664 397724 345716 397730
rect 345664 397666 345716 397672
rect 345664 397384 345716 397390
rect 345664 397326 345716 397332
rect 345676 396166 345704 397326
rect 345664 396160 345716 396166
rect 345664 396102 345716 396108
rect 345572 395616 345624 395622
rect 345572 395558 345624 395564
rect 345664 395616 345716 395622
rect 345664 395558 345716 395564
rect 345676 395282 345704 395558
rect 345768 395418 345796 399570
rect 345860 398041 345888 399724
rect 345940 399628 345992 399634
rect 345940 399570 345992 399576
rect 345846 398032 345902 398041
rect 345846 397967 345902 397976
rect 345848 397724 345900 397730
rect 345848 397666 345900 397672
rect 345860 396098 345888 397666
rect 345952 396574 345980 399570
rect 345940 396568 345992 396574
rect 345940 396510 345992 396516
rect 346044 396216 346072 399724
rect 346124 399628 346176 399634
rect 346124 399570 346176 399576
rect 346308 399628 346360 399634
rect 346308 399570 346360 399576
rect 346136 396778 346164 399570
rect 346214 398984 346270 398993
rect 346214 398919 346216 398928
rect 346268 398919 346270 398928
rect 346216 398890 346268 398896
rect 346216 398676 346268 398682
rect 346216 398618 346268 398624
rect 346228 397730 346256 398618
rect 346216 397724 346268 397730
rect 346216 397666 346268 397672
rect 346124 396772 346176 396778
rect 346124 396714 346176 396720
rect 345952 396188 346072 396216
rect 345848 396092 345900 396098
rect 345848 396034 345900 396040
rect 345848 395956 345900 395962
rect 345848 395898 345900 395904
rect 345756 395412 345808 395418
rect 345756 395354 345808 395360
rect 345664 395276 345716 395282
rect 345664 395218 345716 395224
rect 345860 395078 345888 395898
rect 345848 395072 345900 395078
rect 345848 395014 345900 395020
rect 345952 394890 345980 396188
rect 346032 396092 346084 396098
rect 346032 396034 346084 396040
rect 345584 394862 345980 394890
rect 345584 329118 345612 394862
rect 346044 392714 346072 396034
rect 346122 395448 346178 395457
rect 346122 395383 346178 395392
rect 345860 392686 346072 392714
rect 345664 391740 345716 391746
rect 345664 391682 345716 391688
rect 345572 329112 345624 329118
rect 345572 329054 345624 329060
rect 345478 320784 345534 320793
rect 345478 320719 345534 320728
rect 344928 315716 344980 315722
rect 344928 315658 344980 315664
rect 344744 310140 344796 310146
rect 344744 310082 344796 310088
rect 345676 300354 345704 391682
rect 345756 389904 345808 389910
rect 345756 389846 345808 389852
rect 345768 307154 345796 389846
rect 345860 381721 345888 392686
rect 345940 392080 345992 392086
rect 345940 392022 345992 392028
rect 345846 381712 345902 381721
rect 345846 381647 345902 381656
rect 345848 379568 345900 379574
rect 345848 379510 345900 379516
rect 345756 307148 345808 307154
rect 345756 307090 345808 307096
rect 345664 300348 345716 300354
rect 345664 300290 345716 300296
rect 344652 300212 344704 300218
rect 344652 300154 344704 300160
rect 345860 299130 345888 379510
rect 345952 319394 345980 392022
rect 346032 387252 346084 387258
rect 346032 387194 346084 387200
rect 345940 319388 345992 319394
rect 345940 319330 345992 319336
rect 345940 316804 345992 316810
rect 345940 316746 345992 316752
rect 345848 299124 345900 299130
rect 345848 299066 345900 299072
rect 344468 299056 344520 299062
rect 344468 298998 344520 299004
rect 344284 295112 344336 295118
rect 344284 295054 344336 295060
rect 345952 247722 345980 316746
rect 346044 309602 346072 387194
rect 346136 320929 346164 395383
rect 346320 395010 346348 399570
rect 346412 399430 346440 399724
rect 346642 399752 346670 400044
rect 346734 399945 346762 400044
rect 346720 399936 346776 399945
rect 346720 399871 346776 399880
rect 346826 399820 346854 400044
rect 346918 399906 346946 400044
rect 346906 399900 346958 399906
rect 346906 399842 346958 399848
rect 346780 399809 346854 399820
rect 346492 399706 346544 399712
rect 346596 399724 346670 399752
rect 346766 399800 346854 399809
rect 346822 399792 346854 399800
rect 347010 399786 347038 400044
rect 347102 399945 347130 400044
rect 347088 399936 347144 399945
rect 347088 399871 347144 399880
rect 346964 399758 347038 399786
rect 346964 399752 346992 399758
rect 347194 399752 347222 400044
rect 347286 399838 347314 400044
rect 347274 399832 347326 399838
rect 347274 399774 347326 399780
rect 346766 399735 346822 399744
rect 346872 399724 346992 399752
rect 347148 399724 347222 399752
rect 347378 399752 347406 400044
rect 347470 399906 347498 400044
rect 347458 399900 347510 399906
rect 347458 399842 347510 399848
rect 347562 399786 347590 400044
rect 347654 399906 347682 400044
rect 347642 399900 347694 399906
rect 347642 399842 347694 399848
rect 347746 399786 347774 400044
rect 347838 399945 347866 400044
rect 347824 399936 347880 399945
rect 347824 399871 347880 399880
rect 347562 399758 347636 399786
rect 347378 399724 347452 399752
rect 346400 399424 346452 399430
rect 346400 399366 346452 399372
rect 346400 398812 346452 398818
rect 346400 398754 346452 398760
rect 346412 398138 346440 398754
rect 346400 398132 346452 398138
rect 346400 398074 346452 398080
rect 346504 395078 346532 399706
rect 346596 397866 346624 399724
rect 346768 399628 346820 399634
rect 346768 399570 346820 399576
rect 346674 398984 346730 398993
rect 346674 398919 346676 398928
rect 346728 398919 346730 398928
rect 346676 398890 346728 398896
rect 346584 397860 346636 397866
rect 346584 397802 346636 397808
rect 346584 397724 346636 397730
rect 346584 397666 346636 397672
rect 346596 397526 346624 397666
rect 346584 397520 346636 397526
rect 346584 397462 346636 397468
rect 346780 396506 346808 399570
rect 346872 399401 346900 399724
rect 347044 399696 347096 399702
rect 347044 399638 347096 399644
rect 346952 399628 347004 399634
rect 346952 399570 347004 399576
rect 346858 399392 346914 399401
rect 346858 399327 346914 399336
rect 346964 398256 346992 399570
rect 346872 398228 346992 398256
rect 346768 396500 346820 396506
rect 346768 396442 346820 396448
rect 346872 395298 346900 398228
rect 347056 398154 347084 399638
rect 346964 398126 347084 398154
rect 346964 397458 346992 398126
rect 347044 398064 347096 398070
rect 347044 398006 347096 398012
rect 346952 397452 347004 397458
rect 346952 397394 347004 397400
rect 346596 395270 346900 395298
rect 346492 395072 346544 395078
rect 346398 395040 346454 395049
rect 346308 395004 346360 395010
rect 346492 395014 346544 395020
rect 346398 394975 346454 394984
rect 346308 394946 346360 394952
rect 346214 388512 346270 388521
rect 346214 388447 346270 388456
rect 346228 371890 346256 388447
rect 346412 387122 346440 394975
rect 346492 392420 346544 392426
rect 346492 392362 346544 392368
rect 346400 387116 346452 387122
rect 346400 387058 346452 387064
rect 346216 371884 346268 371890
rect 346216 371826 346268 371832
rect 346122 320920 346178 320929
rect 346122 320855 346178 320864
rect 346504 319190 346532 392362
rect 346492 319184 346544 319190
rect 346492 319126 346544 319132
rect 346596 318986 346624 395270
rect 346676 395072 346728 395078
rect 346676 395014 346728 395020
rect 346768 395072 346820 395078
rect 346768 395014 346820 395020
rect 346688 385898 346716 395014
rect 346780 389162 346808 395014
rect 347056 392544 347084 398006
rect 346964 392516 347084 392544
rect 346768 389156 346820 389162
rect 346768 389098 346820 389104
rect 346676 385892 346728 385898
rect 346676 385834 346728 385840
rect 346584 318980 346636 318986
rect 346584 318922 346636 318928
rect 346032 309596 346084 309602
rect 346032 309538 346084 309544
rect 346964 296682 346992 392516
rect 347148 392426 347176 399724
rect 347320 399628 347372 399634
rect 347320 399570 347372 399576
rect 347226 399528 347282 399537
rect 347226 399463 347228 399472
rect 347280 399463 347282 399472
rect 347228 399434 347280 399440
rect 347226 397760 347282 397769
rect 347226 397695 347282 397704
rect 347136 392420 347188 392426
rect 347136 392362 347188 392368
rect 347240 391490 347268 397695
rect 347332 395049 347360 399570
rect 347424 398721 347452 399724
rect 347504 399696 347556 399702
rect 347504 399638 347556 399644
rect 347410 398712 347466 398721
rect 347410 398647 347466 398656
rect 347516 395729 347544 399638
rect 347502 395720 347558 395729
rect 347502 395655 347558 395664
rect 347608 395078 347636 399758
rect 347700 399758 347774 399786
rect 347700 399514 347728 399758
rect 347930 399752 347958 400044
rect 348022 399906 348050 400044
rect 348010 399900 348062 399906
rect 348010 399842 348062 399848
rect 348114 399838 348142 400044
rect 348206 399838 348234 400044
rect 348298 399906 348326 400044
rect 348286 399900 348338 399906
rect 348286 399842 348338 399848
rect 348390 399838 348418 400044
rect 348482 399945 348510 400044
rect 348468 399936 348524 399945
rect 348468 399871 348524 399880
rect 348102 399832 348154 399838
rect 348102 399774 348154 399780
rect 348194 399832 348246 399838
rect 348194 399774 348246 399780
rect 348378 399832 348430 399838
rect 348574 399786 348602 400044
rect 348378 399774 348430 399780
rect 348528 399758 348602 399786
rect 347930 399724 348004 399752
rect 347872 399628 347924 399634
rect 347872 399570 347924 399576
rect 347700 399486 347820 399514
rect 347688 399424 347740 399430
rect 347688 399366 347740 399372
rect 347700 398070 347728 399366
rect 347688 398064 347740 398070
rect 347688 398006 347740 398012
rect 347792 396681 347820 399486
rect 347884 398177 347912 399570
rect 347870 398168 347926 398177
rect 347870 398103 347926 398112
rect 347872 397588 347924 397594
rect 347872 397530 347924 397536
rect 347778 396672 347834 396681
rect 347778 396607 347834 396616
rect 347596 395072 347648 395078
rect 347318 395040 347374 395049
rect 347884 395026 347912 397530
rect 347596 395014 347648 395020
rect 347318 394975 347374 394984
rect 347792 394998 347912 395026
rect 347688 394392 347740 394398
rect 347688 394334 347740 394340
rect 347056 391462 347268 391490
rect 346952 296676 347004 296682
rect 346952 296618 347004 296624
rect 347056 295322 347084 391462
rect 347700 389178 347728 394334
rect 347792 393718 347820 394998
rect 347870 394904 347926 394913
rect 347870 394839 347926 394848
rect 347780 393712 347832 393718
rect 347780 393654 347832 393660
rect 347240 389150 347728 389178
rect 347136 388612 347188 388618
rect 347136 388554 347188 388560
rect 347148 304366 347176 388554
rect 347136 304360 347188 304366
rect 347136 304302 347188 304308
rect 347240 299198 347268 389150
rect 347412 388680 347464 388686
rect 347412 388622 347464 388628
rect 347320 387388 347372 387394
rect 347320 387330 347372 387336
rect 347332 305998 347360 387330
rect 347424 310078 347452 388622
rect 347884 388482 347912 394839
rect 347976 393854 348004 399724
rect 348240 399696 348292 399702
rect 348292 399656 348464 399684
rect 348240 399638 348292 399644
rect 348148 399628 348200 399634
rect 348148 399570 348200 399576
rect 348056 399492 348108 399498
rect 348056 399434 348108 399440
rect 347964 393848 348016 393854
rect 347964 393790 348016 393796
rect 347964 393712 348016 393718
rect 347964 393654 348016 393660
rect 347872 388476 347924 388482
rect 347872 388418 347924 388424
rect 347502 383344 347558 383353
rect 347502 383279 347558 383288
rect 347412 310072 347464 310078
rect 347412 310014 347464 310020
rect 347516 309738 347544 383279
rect 347976 319122 348004 393654
rect 348068 380186 348096 399434
rect 348160 397526 348188 399570
rect 348332 398472 348384 398478
rect 348332 398414 348384 398420
rect 348148 397520 348200 397526
rect 348148 397462 348200 397468
rect 348344 397361 348372 398414
rect 348330 397352 348386 397361
rect 348330 397287 348386 397296
rect 348146 395448 348202 395457
rect 348146 395383 348202 395392
rect 348160 383042 348188 395383
rect 348240 395276 348292 395282
rect 348240 395218 348292 395224
rect 348252 384334 348280 395218
rect 348332 393848 348384 393854
rect 348332 393790 348384 393796
rect 348240 384328 348292 384334
rect 348240 384270 348292 384276
rect 348148 383036 348200 383042
rect 348148 382978 348200 382984
rect 348056 380180 348108 380186
rect 348056 380122 348108 380128
rect 347964 319116 348016 319122
rect 347964 319058 348016 319064
rect 347596 315376 347648 315382
rect 347596 315318 347648 315324
rect 347504 309732 347556 309738
rect 347504 309674 347556 309680
rect 347320 305992 347372 305998
rect 347320 305934 347372 305940
rect 347228 299192 347280 299198
rect 347228 299134 347280 299140
rect 347044 295316 347096 295322
rect 347044 295258 347096 295264
rect 347608 253230 347636 315318
rect 348344 299402 348372 393790
rect 348436 388793 348464 399656
rect 348528 397458 348556 399758
rect 348666 399684 348694 400044
rect 348758 399752 348786 400044
rect 348850 399820 348878 400044
rect 348942 399945 348970 400044
rect 348928 399936 348984 399945
rect 348928 399871 348984 399880
rect 348850 399792 348924 399820
rect 348758 399724 348832 399752
rect 348620 399656 348694 399684
rect 348620 397633 348648 399656
rect 348700 399356 348752 399362
rect 348700 399298 348752 399304
rect 348606 397624 348662 397633
rect 348606 397559 348662 397568
rect 348608 397520 348660 397526
rect 348608 397462 348660 397468
rect 348516 397452 348568 397458
rect 348516 397394 348568 397400
rect 348516 396772 348568 396778
rect 348516 396714 348568 396720
rect 348422 388784 348478 388793
rect 348422 388719 348478 388728
rect 348422 387560 348478 387569
rect 348422 387495 348478 387504
rect 348436 306066 348464 387495
rect 348528 379409 348556 396714
rect 348620 383246 348648 397462
rect 348712 392086 348740 399298
rect 348804 395282 348832 399724
rect 348896 397594 348924 399792
rect 349034 399684 349062 400044
rect 348988 399656 349062 399684
rect 348884 397588 348936 397594
rect 348884 397530 348936 397536
rect 348884 397452 348936 397458
rect 348884 397394 348936 397400
rect 348792 395276 348844 395282
rect 348792 395218 348844 395224
rect 348700 392080 348752 392086
rect 348700 392022 348752 392028
rect 348896 390554 348924 397394
rect 348988 390794 349016 399656
rect 349126 399616 349154 400044
rect 349218 399684 349246 400044
rect 349310 399945 349338 400044
rect 349296 399936 349352 399945
rect 349296 399871 349352 399880
rect 349402 399752 349430 400044
rect 349356 399724 349430 399752
rect 349218 399656 349292 399684
rect 349080 399588 349154 399616
rect 349080 394398 349108 399588
rect 349160 399016 349212 399022
rect 349160 398958 349212 398964
rect 349172 398857 349200 398958
rect 349158 398848 349214 398857
rect 349158 398783 349214 398792
rect 349160 398404 349212 398410
rect 349160 398346 349212 398352
rect 349172 398138 349200 398346
rect 349160 398132 349212 398138
rect 349160 398074 349212 398080
rect 349264 396930 349292 399656
rect 349172 396902 349292 396930
rect 349172 394874 349200 396902
rect 349250 396808 349306 396817
rect 349250 396743 349306 396752
rect 349160 394868 349212 394874
rect 349160 394810 349212 394816
rect 349068 394392 349120 394398
rect 349068 394334 349120 394340
rect 348976 390788 349028 390794
rect 348976 390730 349028 390736
rect 348896 390526 349016 390554
rect 348608 383240 348660 383246
rect 348608 383182 348660 383188
rect 348608 383036 348660 383042
rect 348608 382978 348660 382984
rect 348514 379400 348570 379409
rect 348514 379335 348570 379344
rect 348516 377460 348568 377466
rect 348516 377402 348568 377408
rect 348424 306060 348476 306066
rect 348424 306002 348476 306008
rect 348332 299396 348384 299402
rect 348332 299338 348384 299344
rect 348528 297362 348556 377402
rect 348620 302938 348648 382978
rect 348700 378072 348752 378078
rect 348700 378014 348752 378020
rect 348608 302932 348660 302938
rect 348608 302874 348660 302880
rect 348712 301646 348740 378014
rect 348792 377596 348844 377602
rect 348792 377538 348844 377544
rect 348700 301640 348752 301646
rect 348700 301582 348752 301588
rect 348804 301578 348832 377538
rect 348884 315512 348936 315518
rect 348884 315454 348936 315460
rect 348792 301572 348844 301578
rect 348792 301514 348844 301520
rect 348516 297356 348568 297362
rect 348516 297298 348568 297304
rect 348896 272542 348924 315454
rect 348988 299266 349016 390526
rect 349264 389174 349292 396743
rect 349356 393378 349384 399724
rect 349494 399684 349522 400044
rect 349586 399906 349614 400044
rect 349678 399906 349706 400044
rect 349770 399906 349798 400044
rect 349574 399900 349626 399906
rect 349574 399842 349626 399848
rect 349666 399900 349718 399906
rect 349666 399842 349718 399848
rect 349758 399900 349810 399906
rect 349758 399842 349810 399848
rect 349862 399786 349890 400044
rect 349954 399906 349982 400044
rect 349942 399900 349994 399906
rect 349942 399842 349994 399848
rect 350046 399838 350074 400044
rect 349724 399758 349890 399786
rect 350034 399832 350086 399838
rect 350034 399774 350086 399780
rect 349494 399656 349568 399684
rect 349436 399560 349488 399566
rect 349436 399502 349488 399508
rect 349448 393650 349476 399502
rect 349436 393644 349488 393650
rect 349436 393586 349488 393592
rect 349344 393372 349396 393378
rect 349344 393314 349396 393320
rect 349436 393372 349488 393378
rect 349436 393314 349488 393320
rect 349264 389146 349384 389174
rect 349356 388550 349384 389146
rect 349344 388544 349396 388550
rect 349344 388486 349396 388492
rect 349448 378865 349476 393314
rect 349540 388657 349568 399656
rect 349620 399492 349672 399498
rect 349620 399434 349672 399440
rect 349632 393378 349660 399434
rect 349620 393372 349672 393378
rect 349620 393314 349672 393320
rect 349620 390516 349672 390522
rect 349620 390458 349672 390464
rect 349526 388648 349582 388657
rect 349526 388583 349582 388592
rect 349434 378856 349490 378865
rect 349434 378791 349490 378800
rect 349632 322017 349660 390458
rect 349724 389026 349752 399758
rect 349804 399696 349856 399702
rect 350138 399684 350166 400044
rect 350230 399752 350258 400044
rect 350322 399906 350350 400044
rect 350310 399900 350362 399906
rect 350310 399842 350362 399848
rect 350414 399838 350442 400044
rect 350402 399832 350454 399838
rect 350402 399774 350454 399780
rect 350506 399752 350534 400044
rect 350598 399906 350626 400044
rect 350586 399900 350638 399906
rect 350586 399842 350638 399848
rect 350690 399838 350718 400044
rect 350782 399906 350810 400044
rect 350874 399945 350902 400044
rect 350860 399936 350916 399945
rect 350770 399900 350822 399906
rect 350860 399871 350916 399880
rect 350770 399842 350822 399848
rect 350966 399838 350994 400044
rect 351058 399906 351086 400044
rect 351150 399906 351178 400044
rect 351242 399906 351270 400044
rect 351046 399900 351098 399906
rect 351046 399842 351098 399848
rect 351138 399900 351190 399906
rect 351138 399842 351190 399848
rect 351230 399900 351282 399906
rect 351230 399842 351282 399848
rect 350678 399832 350730 399838
rect 350678 399774 350730 399780
rect 350954 399832 351006 399838
rect 351334 399786 351362 400044
rect 351426 399906 351454 400044
rect 351414 399900 351466 399906
rect 351414 399842 351466 399848
rect 350954 399774 351006 399780
rect 350816 399764 350868 399770
rect 350230 399724 350304 399752
rect 350506 399724 350580 399752
rect 349804 399638 349856 399644
rect 350092 399656 350166 399684
rect 349816 397905 349844 399638
rect 349988 399492 350040 399498
rect 349988 399434 350040 399440
rect 349896 399424 349948 399430
rect 349896 399366 349948 399372
rect 349802 397896 349858 397905
rect 349802 397831 349858 397840
rect 349908 396778 349936 399366
rect 350000 398449 350028 399434
rect 349986 398440 350042 398449
rect 349986 398375 350042 398384
rect 349986 398304 350042 398313
rect 349986 398239 350042 398248
rect 350000 397633 350028 398239
rect 349986 397624 350042 397633
rect 349986 397559 350042 397568
rect 349896 396772 349948 396778
rect 349896 396714 349948 396720
rect 349986 395448 350042 395457
rect 349986 395383 350042 395392
rect 349712 389020 349764 389026
rect 349712 388962 349764 388968
rect 349804 387116 349856 387122
rect 349804 387058 349856 387064
rect 349618 322008 349674 322017
rect 349618 321943 349674 321952
rect 349816 305930 349844 387058
rect 349896 383240 349948 383246
rect 349896 383182 349948 383188
rect 349804 305924 349856 305930
rect 349804 305866 349856 305872
rect 349908 303006 349936 383182
rect 350000 378729 350028 395383
rect 350092 390522 350120 399656
rect 350276 399616 350304 399724
rect 350448 399628 350500 399634
rect 350276 399588 350350 399616
rect 350322 399548 350350 399588
rect 350448 399570 350500 399576
rect 350322 399520 350396 399548
rect 350264 399424 350316 399430
rect 350264 399366 350316 399372
rect 350172 397452 350224 397458
rect 350172 397394 350224 397400
rect 350184 396642 350212 397394
rect 350172 396636 350224 396642
rect 350172 396578 350224 396584
rect 350080 390516 350132 390522
rect 350080 390458 350132 390464
rect 350080 386572 350132 386578
rect 350080 386514 350132 386520
rect 349986 378720 350042 378729
rect 349986 378655 350042 378664
rect 349986 377632 350042 377641
rect 349986 377567 350042 377576
rect 349896 303000 349948 303006
rect 349896 302942 349948 302948
rect 348976 299260 349028 299266
rect 348976 299202 349028 299208
rect 350000 298926 350028 377567
rect 350092 317150 350120 386514
rect 350172 377528 350224 377534
rect 350172 377470 350224 377476
rect 350080 317144 350132 317150
rect 350080 317086 350132 317092
rect 350184 312730 350212 377470
rect 350276 342922 350304 399366
rect 350368 391814 350396 399520
rect 350460 398682 350488 399570
rect 350448 398676 350500 398682
rect 350448 398618 350500 398624
rect 350552 394754 350580 399724
rect 350816 399706 350868 399712
rect 351104 399758 351362 399786
rect 350724 399696 350776 399702
rect 350724 399638 350776 399644
rect 350632 399628 350684 399634
rect 350632 399570 350684 399576
rect 350460 394726 350580 394754
rect 350460 393174 350488 394726
rect 350644 394694 350672 399570
rect 350736 396817 350764 399638
rect 350828 397594 350856 399706
rect 350908 399696 350960 399702
rect 350908 399638 350960 399644
rect 350920 399480 350948 399638
rect 350920 399452 351040 399480
rect 350908 399356 350960 399362
rect 350908 399298 350960 399304
rect 350816 397588 350868 397594
rect 350816 397530 350868 397536
rect 350722 396808 350778 396817
rect 350722 396743 350778 396752
rect 350552 394666 350672 394694
rect 350448 393168 350500 393174
rect 350448 393110 350500 393116
rect 350356 391808 350408 391814
rect 350356 391750 350408 391756
rect 350552 389842 350580 394666
rect 350816 394392 350868 394398
rect 350816 394334 350868 394340
rect 350828 394126 350856 394334
rect 350816 394120 350868 394126
rect 350816 394062 350868 394068
rect 350816 393984 350868 393990
rect 350816 393926 350868 393932
rect 350724 393780 350776 393786
rect 350724 393722 350776 393728
rect 350630 393544 350686 393553
rect 350630 393479 350632 393488
rect 350684 393479 350686 393488
rect 350632 393450 350684 393456
rect 350540 389836 350592 389842
rect 350540 389778 350592 389784
rect 350736 356726 350764 393722
rect 350828 362234 350856 393926
rect 350920 373425 350948 399298
rect 351012 394210 351040 399452
rect 351104 397905 351132 399758
rect 351518 399752 351546 400044
rect 351610 399945 351638 400044
rect 351596 399936 351652 399945
rect 351702 399906 351730 400044
rect 351596 399871 351652 399880
rect 351690 399900 351742 399906
rect 351690 399842 351742 399848
rect 351644 399764 351696 399770
rect 351518 399724 351592 399752
rect 351184 399696 351236 399702
rect 351184 399638 351236 399644
rect 351196 399362 351224 399638
rect 351276 399628 351328 399634
rect 351460 399628 351512 399634
rect 351328 399588 351408 399616
rect 351276 399570 351328 399576
rect 351274 399528 351330 399537
rect 351274 399463 351330 399472
rect 351288 399362 351316 399463
rect 351184 399356 351236 399362
rect 351184 399298 351236 399304
rect 351276 399356 351328 399362
rect 351276 399298 351328 399304
rect 351184 399220 351236 399226
rect 351184 399162 351236 399168
rect 351196 398274 351224 399162
rect 351184 398268 351236 398274
rect 351184 398210 351236 398216
rect 351090 397896 351146 397905
rect 351090 397831 351146 397840
rect 351276 397588 351328 397594
rect 351276 397530 351328 397536
rect 351184 397520 351236 397526
rect 351184 397462 351236 397468
rect 351012 394182 351132 394210
rect 351000 394120 351052 394126
rect 351000 394062 351052 394068
rect 351012 379137 351040 394062
rect 351104 393854 351132 394182
rect 351092 393848 351144 393854
rect 351092 393790 351144 393796
rect 350998 379128 351054 379137
rect 350998 379063 351054 379072
rect 350906 373416 350962 373425
rect 350906 373351 350962 373360
rect 350816 362228 350868 362234
rect 350816 362170 350868 362176
rect 350724 356720 350776 356726
rect 350724 356662 350776 356668
rect 350264 342916 350316 342922
rect 350264 342858 350316 342864
rect 350264 336048 350316 336054
rect 350264 335990 350316 335996
rect 350172 312724 350224 312730
rect 350172 312666 350224 312672
rect 349988 298920 350040 298926
rect 349988 298862 350040 298868
rect 350276 286550 350304 335990
rect 351196 306270 351224 397462
rect 351288 393718 351316 397530
rect 351380 393990 351408 399588
rect 351460 399570 351512 399576
rect 351368 393984 351420 393990
rect 351368 393926 351420 393932
rect 351276 393712 351328 393718
rect 351276 393654 351328 393660
rect 351368 388476 351420 388482
rect 351368 388418 351420 388424
rect 351276 388204 351328 388210
rect 351276 388146 351328 388152
rect 351184 306264 351236 306270
rect 351184 306206 351236 306212
rect 351288 301850 351316 388146
rect 351380 314022 351408 388418
rect 351472 379273 351500 399570
rect 351458 379264 351514 379273
rect 351458 379199 351514 379208
rect 351564 347070 351592 399724
rect 351644 399706 351696 399712
rect 351656 394126 351684 399706
rect 351794 399684 351822 400044
rect 351748 399656 351822 399684
rect 351886 399684 351914 400044
rect 351978 399752 352006 400044
rect 352070 399906 352098 400044
rect 352058 399900 352110 399906
rect 352058 399842 352110 399848
rect 352162 399752 352190 400044
rect 352254 399906 352282 400044
rect 352242 399900 352294 399906
rect 352242 399842 352294 399848
rect 351978 399724 352052 399752
rect 352162 399724 352236 399752
rect 351886 399656 351960 399684
rect 351644 394120 351696 394126
rect 351644 394062 351696 394068
rect 351644 393848 351696 393854
rect 351644 393790 351696 393796
rect 351552 347064 351604 347070
rect 351552 347006 351604 347012
rect 351656 340202 351684 393790
rect 351748 393786 351776 399656
rect 351828 398676 351880 398682
rect 351828 398618 351880 398624
rect 351840 398041 351868 398618
rect 351826 398032 351882 398041
rect 351826 397967 351882 397976
rect 351932 397594 351960 399656
rect 352024 398342 352052 399724
rect 352104 399424 352156 399430
rect 352104 399366 352156 399372
rect 352012 398336 352064 398342
rect 352012 398278 352064 398284
rect 352012 398064 352064 398070
rect 352012 398006 352064 398012
rect 351920 397588 351972 397594
rect 351920 397530 351972 397536
rect 352024 394233 352052 398006
rect 352010 394224 352066 394233
rect 352010 394159 352066 394168
rect 351736 393780 351788 393786
rect 351736 393722 351788 393728
rect 352116 359582 352144 399366
rect 352208 398410 352236 399724
rect 352346 399684 352374 400044
rect 352438 399906 352466 400044
rect 352426 399900 352478 399906
rect 352426 399842 352478 399848
rect 352300 399656 352374 399684
rect 352300 398449 352328 399656
rect 352530 399616 352558 400044
rect 352622 399684 352650 400044
rect 352714 399786 352742 400044
rect 352806 399906 352834 400044
rect 352794 399900 352846 399906
rect 352794 399842 352846 399848
rect 352714 399758 352788 399786
rect 352622 399656 352696 399684
rect 352530 399588 352604 399616
rect 352380 399560 352432 399566
rect 352380 399502 352432 399508
rect 352286 398440 352342 398449
rect 352196 398404 352248 398410
rect 352286 398375 352342 398384
rect 352196 398346 352248 398352
rect 352288 398268 352340 398274
rect 352288 398210 352340 398216
rect 352196 397588 352248 397594
rect 352196 397530 352248 397536
rect 352208 377369 352236 397530
rect 352300 384441 352328 398210
rect 352392 397526 352420 399502
rect 352472 399424 352524 399430
rect 352472 399366 352524 399372
rect 352380 397520 352432 397526
rect 352380 397462 352432 397468
rect 352286 384432 352342 384441
rect 352286 384367 352342 384376
rect 352194 377360 352250 377369
rect 352194 377295 352250 377304
rect 352104 359576 352156 359582
rect 352104 359518 352156 359524
rect 351644 340196 351696 340202
rect 351644 340138 351696 340144
rect 352484 319054 352512 399366
rect 352576 396545 352604 399588
rect 352668 398274 352696 399656
rect 352656 398268 352708 398274
rect 352656 398210 352708 398216
rect 352656 397996 352708 398002
rect 352656 397938 352708 397944
rect 352562 396536 352618 396545
rect 352562 396471 352618 396480
rect 352668 393972 352696 397938
rect 352760 397866 352788 399758
rect 352898 399752 352926 400044
rect 352990 399906 353018 400044
rect 352978 399900 353030 399906
rect 352978 399842 353030 399848
rect 353082 399752 353110 400044
rect 352852 399724 352926 399752
rect 353036 399724 353110 399752
rect 352748 397860 352800 397866
rect 352748 397802 352800 397808
rect 352748 397520 352800 397526
rect 352748 397462 352800 397468
rect 352576 393944 352696 393972
rect 352472 319048 352524 319054
rect 352472 318990 352524 318996
rect 351460 315444 351512 315450
rect 351460 315386 351512 315392
rect 351368 314016 351420 314022
rect 351368 313958 351420 313964
rect 351276 301844 351328 301850
rect 351276 301786 351328 301792
rect 349252 286544 349304 286550
rect 349252 286486 349304 286492
rect 350264 286544 350316 286550
rect 350264 286486 350316 286492
rect 349264 286346 349292 286486
rect 349252 286340 349304 286346
rect 349252 286282 349304 286288
rect 348884 272536 348936 272542
rect 348884 272478 348936 272484
rect 347596 253224 347648 253230
rect 347596 253166 347648 253172
rect 345940 247716 345992 247722
rect 345940 247658 345992 247664
rect 342350 219328 342406 219337
rect 342350 219263 342406 219272
rect 342260 203584 342312 203590
rect 342260 203526 342312 203532
rect 341524 100700 341576 100706
rect 341524 100642 341576 100648
rect 340970 72448 341026 72457
rect 340970 72383 341026 72392
rect 340984 3398 341012 72383
rect 342272 16574 342300 203526
rect 345020 148436 345072 148442
rect 345020 148378 345072 148384
rect 343638 113792 343694 113801
rect 343638 113727 343694 113736
rect 343652 16574 343680 113727
rect 345032 16574 345060 148378
rect 347780 105596 347832 105602
rect 347780 105538 347832 105544
rect 347792 16574 347820 105538
rect 342272 16546 342944 16574
rect 343652 16546 344600 16574
rect 345032 16546 345336 16574
rect 347792 16546 348096 16574
rect 340972 3392 341024 3398
rect 340972 3334 341024 3340
rect 342168 3392 342220 3398
rect 342168 3334 342220 3340
rect 340892 3182 341012 3210
rect 340984 480 341012 3182
rect 342180 480 342208 3334
rect 339838 354 339950 480
rect 339512 326 339950 354
rect 339838 -960 339950 326
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 354 342944 16546
rect 344572 480 344600 16546
rect 343334 354 343446 480
rect 342916 326 343446 354
rect 343334 -960 343446 326
rect 344530 -960 344642 480
rect 345308 354 345336 16546
rect 346952 3936 347004 3942
rect 346952 3878 347004 3884
rect 346964 480 346992 3878
rect 348068 480 348096 16546
rect 349160 4004 349212 4010
rect 349160 3946 349212 3952
rect 349172 1986 349200 3946
rect 349264 3398 349292 286282
rect 351472 251870 351500 315386
rect 352576 301782 352604 393944
rect 352656 393644 352708 393650
rect 352656 393586 352708 393592
rect 352668 303074 352696 393586
rect 352760 306134 352788 397462
rect 352852 394398 352880 399724
rect 352932 399628 352984 399634
rect 352932 399570 352984 399576
rect 352944 399537 352972 399570
rect 352930 399528 352986 399537
rect 352930 399463 352986 399472
rect 352932 397860 352984 397866
rect 352932 397802 352984 397808
rect 352840 394392 352892 394398
rect 352840 394334 352892 394340
rect 352840 392624 352892 392630
rect 352840 392566 352892 392572
rect 352852 308650 352880 392566
rect 352944 319326 352972 397802
rect 353036 397497 353064 399724
rect 353174 399684 353202 400044
rect 353266 399945 353294 400044
rect 353252 399936 353308 399945
rect 353252 399871 353308 399880
rect 353358 399820 353386 400044
rect 353128 399656 353202 399684
rect 353312 399792 353386 399820
rect 353022 397488 353078 397497
rect 353022 397423 353078 397432
rect 353128 392329 353156 399656
rect 353206 399528 353262 399537
rect 353206 399463 353262 399472
rect 353220 399362 353248 399463
rect 353208 399356 353260 399362
rect 353208 399298 353260 399304
rect 353312 397497 353340 399792
rect 353450 399752 353478 400044
rect 353404 399724 353478 399752
rect 353404 398993 353432 399724
rect 353542 399650 353570 400044
rect 353634 399752 353662 400044
rect 353726 399820 353754 400044
rect 353818 399945 353846 400044
rect 353804 399936 353860 399945
rect 353910 399906 353938 400044
rect 353804 399871 353860 399880
rect 353898 399900 353950 399906
rect 353898 399842 353950 399848
rect 353726 399792 353800 399820
rect 353772 399786 353800 399792
rect 353772 399758 353892 399786
rect 353634 399724 353708 399752
rect 353496 399622 353570 399650
rect 353390 398984 353446 398993
rect 353390 398919 353446 398928
rect 353392 398268 353444 398274
rect 353392 398210 353444 398216
rect 353298 397488 353354 397497
rect 353298 397423 353354 397432
rect 353404 394210 353432 398210
rect 353496 395214 353524 399622
rect 353576 399492 353628 399498
rect 353576 399434 353628 399440
rect 353588 399265 353616 399434
rect 353574 399256 353630 399265
rect 353574 399191 353630 399200
rect 353484 395208 353536 395214
rect 353484 395150 353536 395156
rect 353680 394398 353708 399724
rect 353760 399696 353812 399702
rect 353760 399638 353812 399644
rect 353772 395146 353800 399638
rect 353760 395140 353812 395146
rect 353760 395082 353812 395088
rect 353668 394392 353720 394398
rect 353668 394334 353720 394340
rect 353312 394182 353432 394210
rect 353114 392320 353170 392329
rect 353114 392255 353170 392264
rect 353312 390289 353340 394182
rect 353392 393984 353444 393990
rect 353392 393926 353444 393932
rect 353298 390280 353354 390289
rect 353298 390215 353354 390224
rect 353404 321026 353432 393926
rect 353576 393712 353628 393718
rect 353864 393666 353892 399758
rect 354002 399752 354030 400044
rect 354094 399906 354122 400044
rect 354082 399900 354134 399906
rect 354082 399842 354134 399848
rect 354186 399752 354214 400044
rect 354278 399906 354306 400044
rect 354370 399945 354398 400044
rect 354356 399936 354412 399945
rect 354266 399900 354318 399906
rect 354356 399871 354412 399880
rect 354266 399842 354318 399848
rect 354462 399786 354490 400044
rect 353576 393654 353628 393660
rect 353588 379574 353616 393654
rect 353772 393638 353892 393666
rect 353956 399724 354030 399752
rect 354140 399724 354214 399752
rect 354324 399758 354490 399786
rect 353772 391513 353800 393638
rect 353956 393530 353984 399724
rect 354036 399628 354088 399634
rect 354036 399570 354088 399576
rect 353864 393502 353984 393530
rect 353864 391785 353892 393502
rect 353944 393372 353996 393378
rect 353944 393314 353996 393320
rect 353850 391776 353906 391785
rect 353850 391711 353906 391720
rect 353758 391504 353814 391513
rect 353758 391439 353814 391448
rect 353576 379568 353628 379574
rect 353576 379510 353628 379516
rect 353392 321020 353444 321026
rect 353392 320962 353444 320968
rect 352932 319320 352984 319326
rect 352932 319262 352984 319268
rect 352840 308644 352892 308650
rect 352840 308586 352892 308592
rect 352748 306128 352800 306134
rect 352748 306070 352800 306076
rect 353956 305454 353984 393314
rect 354048 391649 354076 399570
rect 354140 393990 354168 399724
rect 354220 399424 354272 399430
rect 354220 399366 354272 399372
rect 354232 395321 354260 399366
rect 354324 395593 354352 399758
rect 354404 399696 354456 399702
rect 354554 399684 354582 400044
rect 354404 399638 354456 399644
rect 354508 399656 354582 399684
rect 354310 395584 354366 395593
rect 354310 395519 354366 395528
rect 354218 395312 354274 395321
rect 354218 395247 354274 395256
rect 354416 394694 354444 399638
rect 354232 394666 354444 394694
rect 354128 393984 354180 393990
rect 354128 393926 354180 393932
rect 354034 391640 354090 391649
rect 354034 391575 354090 391584
rect 354232 391202 354260 394666
rect 354508 394482 354536 399656
rect 354646 399616 354674 400044
rect 354738 399752 354766 400044
rect 354830 399945 354858 400044
rect 354816 399936 354872 399945
rect 354816 399871 354872 399880
rect 354922 399820 354950 400044
rect 354876 399792 354950 399820
rect 354738 399724 354812 399752
rect 354600 399588 354674 399616
rect 354600 397526 354628 399588
rect 354784 399430 354812 399724
rect 354772 399424 354824 399430
rect 354772 399366 354824 399372
rect 354876 399242 354904 399792
rect 355014 399752 355042 400044
rect 354784 399214 354904 399242
rect 354968 399724 355042 399752
rect 354784 398546 354812 399214
rect 354968 399106 354996 399724
rect 355106 399684 355134 400044
rect 355198 399752 355226 400044
rect 355290 399945 355318 400044
rect 355276 399936 355332 399945
rect 355276 399871 355332 399880
rect 355382 399752 355410 400044
rect 355474 399906 355502 400044
rect 355462 399900 355514 399906
rect 355462 399842 355514 399848
rect 355566 399752 355594 400044
rect 355198 399724 355272 399752
rect 354876 399078 354996 399106
rect 355060 399656 355134 399684
rect 354772 398540 354824 398546
rect 354772 398482 354824 398488
rect 354588 397520 354640 397526
rect 354588 397462 354640 397468
rect 354416 394454 354536 394482
rect 354416 391354 354444 394454
rect 354496 394392 354548 394398
rect 354496 394334 354548 394340
rect 354588 394392 354640 394398
rect 354588 394334 354640 394340
rect 354324 391326 354444 391354
rect 354220 391196 354272 391202
rect 354220 391138 354272 391144
rect 354034 390280 354090 390289
rect 354034 390215 354090 390224
rect 354220 390244 354272 390250
rect 354048 310010 354076 390215
rect 354220 390186 354272 390192
rect 354128 389836 354180 389842
rect 354128 389778 354180 389784
rect 354140 315586 354168 389778
rect 354232 318034 354260 390186
rect 354324 389745 354352 391326
rect 354404 391196 354456 391202
rect 354404 391138 354456 391144
rect 354310 389736 354366 389745
rect 354310 389671 354366 389680
rect 354220 318028 354272 318034
rect 354220 317970 354272 317976
rect 354128 315580 354180 315586
rect 354128 315522 354180 315528
rect 354036 310004 354088 310010
rect 354036 309946 354088 309952
rect 353944 305448 353996 305454
rect 353944 305390 353996 305396
rect 354416 304910 354444 391138
rect 354508 383110 354536 394334
rect 354600 393378 354628 394334
rect 354588 393372 354640 393378
rect 354588 393314 354640 393320
rect 354496 383104 354548 383110
rect 354496 383046 354548 383052
rect 354876 319666 354904 399078
rect 354954 396672 355010 396681
rect 354954 396607 355010 396616
rect 354968 387394 354996 396607
rect 355060 388210 355088 399656
rect 355244 399566 355272 399724
rect 355336 399724 355410 399752
rect 355520 399724 355594 399752
rect 355232 399560 355284 399566
rect 355232 399502 355284 399508
rect 355336 399344 355364 399724
rect 355416 399560 355468 399566
rect 355416 399502 355468 399508
rect 355244 399316 355364 399344
rect 355244 389174 355272 399316
rect 355322 399256 355378 399265
rect 355322 399191 355378 399200
rect 355336 398274 355364 399191
rect 355324 398268 355376 398274
rect 355324 398210 355376 398216
rect 355428 398206 355456 399502
rect 355416 398200 355468 398206
rect 355416 398142 355468 398148
rect 355520 397746 355548 399724
rect 355658 399684 355686 400044
rect 355750 399906 355778 400044
rect 355738 399900 355790 399906
rect 355738 399842 355790 399848
rect 355842 399752 355870 400044
rect 355612 399656 355686 399684
rect 355796 399724 355870 399752
rect 355612 398002 355640 399656
rect 355692 399560 355744 399566
rect 355692 399502 355744 399508
rect 355704 398857 355732 399502
rect 355690 398848 355746 398857
rect 355690 398783 355746 398792
rect 355600 397996 355652 398002
rect 355600 397938 355652 397944
rect 355520 397718 355732 397746
rect 355508 396228 355560 396234
rect 355508 396170 355560 396176
rect 355416 393984 355468 393990
rect 355416 393926 355468 393932
rect 355324 393372 355376 393378
rect 355324 393314 355376 393320
rect 355152 389146 355272 389174
rect 355048 388204 355100 388210
rect 355048 388146 355100 388152
rect 354956 387388 355008 387394
rect 354956 387330 355008 387336
rect 354864 319660 354916 319666
rect 354864 319602 354916 319608
rect 354404 304904 354456 304910
rect 354404 304846 354456 304852
rect 355152 304638 355180 389146
rect 355336 305833 355364 393314
rect 355428 310350 355456 393926
rect 355520 311438 355548 396170
rect 355600 396092 355652 396098
rect 355600 396034 355652 396040
rect 355612 380225 355640 396034
rect 355704 386578 355732 397718
rect 355692 386572 355744 386578
rect 355692 386514 355744 386520
rect 355598 380216 355654 380225
rect 355598 380151 355654 380160
rect 355508 311432 355560 311438
rect 355508 311374 355560 311380
rect 355416 310344 355468 310350
rect 355416 310286 355468 310292
rect 355796 306202 355824 399724
rect 355934 399684 355962 400044
rect 355888 399656 355962 399684
rect 356026 399684 356054 400044
rect 356118 399838 356146 400044
rect 356106 399832 356158 399838
rect 356106 399774 356158 399780
rect 356210 399786 356238 400044
rect 356302 399906 356330 400044
rect 356290 399900 356342 399906
rect 356290 399842 356342 399848
rect 356394 399786 356422 400044
rect 356486 399906 356514 400044
rect 356578 399906 356606 400044
rect 356670 399945 356698 400044
rect 356656 399936 356712 399945
rect 356474 399900 356526 399906
rect 356474 399842 356526 399848
rect 356566 399900 356618 399906
rect 356762 399906 356790 400044
rect 356656 399871 356712 399880
rect 356750 399900 356802 399906
rect 356566 399842 356618 399848
rect 356750 399842 356802 399848
rect 356854 399786 356882 400044
rect 356946 399838 356974 400044
rect 356210 399758 356284 399786
rect 356152 399696 356204 399702
rect 356026 399656 356100 399684
rect 355888 394618 355916 399656
rect 355968 399560 356020 399566
rect 355968 399502 356020 399508
rect 355980 397225 356008 399502
rect 355966 397216 356022 397225
rect 355966 397151 356022 397160
rect 355888 394590 356008 394618
rect 355876 394460 355928 394466
rect 355876 394402 355928 394408
rect 355888 393378 355916 394402
rect 355980 393689 356008 394590
rect 356072 393990 356100 399656
rect 356152 399638 356204 399644
rect 356164 397322 356192 399638
rect 356256 398070 356284 399758
rect 356348 399758 356422 399786
rect 356520 399764 356572 399770
rect 356244 398064 356296 398070
rect 356244 398006 356296 398012
rect 356348 397848 356376 399758
rect 356520 399706 356572 399712
rect 356624 399758 356882 399786
rect 356934 399832 356986 399838
rect 356934 399774 356986 399780
rect 356428 399696 356480 399702
rect 356428 399638 356480 399644
rect 356256 397820 356376 397848
rect 356152 397316 356204 397322
rect 356152 397258 356204 397264
rect 356256 396370 356284 397820
rect 356336 397724 356388 397730
rect 356336 397666 356388 397672
rect 356244 396364 356296 396370
rect 356244 396306 356296 396312
rect 356060 393984 356112 393990
rect 356060 393926 356112 393932
rect 355966 393680 356022 393689
rect 355966 393615 356022 393624
rect 355876 393372 355928 393378
rect 355876 393314 355928 393320
rect 356348 390250 356376 397666
rect 356440 394505 356468 399638
rect 356532 397934 356560 399706
rect 356520 397928 356572 397934
rect 356520 397870 356572 397876
rect 356624 397662 356652 399758
rect 356796 399696 356848 399702
rect 357038 399684 357066 400044
rect 357130 399945 357158 400044
rect 357116 399936 357172 399945
rect 357116 399871 357172 399880
rect 357222 399752 357250 400044
rect 357314 399906 357342 400044
rect 357406 399906 357434 400044
rect 357302 399900 357354 399906
rect 357302 399842 357354 399848
rect 357394 399900 357446 399906
rect 357394 399842 357446 399848
rect 357498 399786 357526 400044
rect 357452 399758 357526 399786
rect 357590 399786 357618 400044
rect 357682 399906 357710 400044
rect 357670 399900 357722 399906
rect 357670 399842 357722 399848
rect 357774 399838 357802 400044
rect 357866 399945 357894 400044
rect 357852 399936 357908 399945
rect 357958 399906 357986 400044
rect 357852 399871 357908 399880
rect 357946 399900 357998 399906
rect 357946 399842 357998 399848
rect 357762 399832 357814 399838
rect 357590 399758 357664 399786
rect 358050 399786 358078 400044
rect 358142 399906 358170 400044
rect 358130 399900 358182 399906
rect 358130 399842 358182 399848
rect 357762 399774 357814 399780
rect 357222 399724 357388 399752
rect 356796 399638 356848 399644
rect 356992 399656 357066 399684
rect 356702 398168 356758 398177
rect 356702 398103 356758 398112
rect 356612 397656 356664 397662
rect 356612 397598 356664 397604
rect 356612 397520 356664 397526
rect 356612 397462 356664 397468
rect 356624 397390 356652 397462
rect 356612 397384 356664 397390
rect 356612 397326 356664 397332
rect 356716 397236 356744 398103
rect 356808 397662 356836 399638
rect 356796 397656 356848 397662
rect 356796 397598 356848 397604
rect 356888 397588 356940 397594
rect 356888 397530 356940 397536
rect 356796 397316 356848 397322
rect 356796 397258 356848 397264
rect 356624 397208 356744 397236
rect 356426 394496 356482 394505
rect 356426 394431 356482 394440
rect 356336 390244 356388 390250
rect 356336 390186 356388 390192
rect 356624 314226 356652 397208
rect 356808 395298 356836 397258
rect 356716 395270 356836 395298
rect 356612 314220 356664 314226
rect 356612 314162 356664 314168
rect 355784 306196 355836 306202
rect 355784 306138 355836 306144
rect 355322 305824 355378 305833
rect 355322 305759 355378 305768
rect 355140 304632 355192 304638
rect 355140 304574 355192 304580
rect 356716 303210 356744 395270
rect 356796 395208 356848 395214
rect 356796 395150 356848 395156
rect 356808 307494 356836 395150
rect 356900 393825 356928 397530
rect 356992 396098 357020 399656
rect 357164 399628 357216 399634
rect 357164 399570 357216 399576
rect 357072 398404 357124 398410
rect 357072 398346 357124 398352
rect 356980 396092 357032 396098
rect 356980 396034 357032 396040
rect 357084 394694 357112 398346
rect 357176 398070 357204 399570
rect 357256 399492 357308 399498
rect 357256 399434 357308 399440
rect 357164 398064 357216 398070
rect 357164 398006 357216 398012
rect 357164 397656 357216 397662
rect 357164 397598 357216 397604
rect 356992 394666 357112 394694
rect 356886 393816 356942 393825
rect 356886 393751 356942 393760
rect 356888 391196 356940 391202
rect 356888 391138 356940 391144
rect 356900 310214 356928 391138
rect 356992 311710 357020 394666
rect 357072 393780 357124 393786
rect 357072 393722 357124 393728
rect 357084 318782 357112 393722
rect 357176 389174 357204 397598
rect 357268 396710 357296 399434
rect 357360 398478 357388 399724
rect 357348 398472 357400 398478
rect 357348 398414 357400 398420
rect 357348 398064 357400 398070
rect 357348 398006 357400 398012
rect 357360 397594 357388 398006
rect 357348 397588 357400 397594
rect 357348 397530 357400 397536
rect 357348 397384 357400 397390
rect 357348 397326 357400 397332
rect 357256 396704 357308 396710
rect 357256 396646 357308 396652
rect 357360 391202 357388 397326
rect 357452 396438 357480 399758
rect 357636 399752 357664 399758
rect 358004 399758 358078 399786
rect 357636 399724 357710 399752
rect 357682 399684 357710 399724
rect 357682 399656 357756 399684
rect 357532 399628 357584 399634
rect 357532 399570 357584 399576
rect 357440 396432 357492 396438
rect 357440 396374 357492 396380
rect 357544 392465 357572 399570
rect 357624 399560 357676 399566
rect 357624 399502 357676 399508
rect 357636 398410 357664 399502
rect 357624 398404 357676 398410
rect 357624 398346 357676 398352
rect 357624 398268 357676 398274
rect 357624 398210 357676 398216
rect 357530 392456 357586 392465
rect 357530 392391 357586 392400
rect 357348 391196 357400 391202
rect 357348 391138 357400 391144
rect 357636 390554 357664 398210
rect 357728 395418 357756 399656
rect 357808 399628 357860 399634
rect 357808 399570 357860 399576
rect 357820 398954 357848 399570
rect 357808 398948 357860 398954
rect 357808 398890 357860 398896
rect 358004 398528 358032 399758
rect 358234 399752 358262 400044
rect 358326 399838 358354 400044
rect 358418 399945 358446 400044
rect 358404 399936 358460 399945
rect 358404 399871 358460 399880
rect 358314 399832 358366 399838
rect 358314 399774 358366 399780
rect 358188 399724 358262 399752
rect 358188 399090 358216 399724
rect 358360 399696 358412 399702
rect 358510 399650 358538 400044
rect 358602 399752 358630 400044
rect 358694 399906 358722 400044
rect 358682 399900 358734 399906
rect 358682 399842 358734 399848
rect 358602 399724 358676 399752
rect 358360 399638 358412 399644
rect 358268 399628 358320 399634
rect 358268 399570 358320 399576
rect 358176 399084 358228 399090
rect 358176 399026 358228 399032
rect 357820 398500 358032 398528
rect 358176 398540 358228 398546
rect 357716 395412 357768 395418
rect 357716 395354 357768 395360
rect 357820 394694 357848 398500
rect 358176 398482 358228 398488
rect 357992 398404 358044 398410
rect 357992 398346 358044 398352
rect 358004 397497 358032 398346
rect 357990 397488 358046 397497
rect 357990 397423 358046 397432
rect 357900 395412 357952 395418
rect 357900 395354 357952 395360
rect 357544 390526 357664 390554
rect 357728 394666 357848 394694
rect 357544 389174 357572 390526
rect 357176 389146 357296 389174
rect 357268 378078 357296 389146
rect 357452 389146 357572 389174
rect 357256 378072 357308 378078
rect 357256 378014 357308 378020
rect 357452 320890 357480 389146
rect 357624 387524 357676 387530
rect 357624 387466 357676 387472
rect 357636 381585 357664 387466
rect 357728 387122 357756 394666
rect 357912 390554 357940 395354
rect 358188 394058 358216 398482
rect 358280 396234 358308 399570
rect 358372 396760 358400 399638
rect 358464 399622 358538 399650
rect 358464 397390 358492 399622
rect 358452 397384 358504 397390
rect 358452 397326 358504 397332
rect 358372 396732 358492 396760
rect 358358 396672 358414 396681
rect 358358 396607 358414 396616
rect 358268 396228 358320 396234
rect 358268 396170 358320 396176
rect 358268 396092 358320 396098
rect 358268 396034 358320 396040
rect 358176 394052 358228 394058
rect 358176 393994 358228 394000
rect 358176 393848 358228 393854
rect 358176 393790 358228 393796
rect 358188 390554 358216 393790
rect 357820 390526 357940 390554
rect 358096 390526 358216 390554
rect 357820 387297 357848 390526
rect 357806 387288 357862 387297
rect 357806 387223 357862 387232
rect 357716 387116 357768 387122
rect 357716 387058 357768 387064
rect 357622 381576 357678 381585
rect 357622 381511 357678 381520
rect 357440 320884 357492 320890
rect 357440 320826 357492 320832
rect 357072 318776 357124 318782
rect 357072 318718 357124 318724
rect 356980 311704 357032 311710
rect 356980 311646 357032 311652
rect 356888 310208 356940 310214
rect 356888 310150 356940 310156
rect 356796 307488 356848 307494
rect 356796 307430 356848 307436
rect 358096 307358 358124 390526
rect 358280 389174 358308 396034
rect 358188 389146 358308 389174
rect 358188 311574 358216 389146
rect 358372 372570 358400 396607
rect 358360 372564 358412 372570
rect 358360 372506 358412 372512
rect 358176 311568 358228 311574
rect 358176 311510 358228 311516
rect 358084 307352 358136 307358
rect 358084 307294 358136 307300
rect 356704 303204 356756 303210
rect 356704 303146 356756 303152
rect 352656 303068 352708 303074
rect 352656 303010 352708 303016
rect 358464 302122 358492 396732
rect 358542 395312 358598 395321
rect 358542 395247 358598 395256
rect 358556 387530 358584 395247
rect 358648 395214 358676 399724
rect 358786 399684 358814 400044
rect 358878 399786 358906 400044
rect 358970 399906 358998 400044
rect 358958 399900 359010 399906
rect 358958 399842 359010 399848
rect 358878 399758 358952 399786
rect 358786 399656 358860 399684
rect 358728 399492 358780 399498
rect 358728 399434 358780 399440
rect 358636 395208 358688 395214
rect 358636 395150 358688 395156
rect 358544 387524 358596 387530
rect 358544 387466 358596 387472
rect 358740 312866 358768 399434
rect 358832 398274 358860 399656
rect 358820 398268 358872 398274
rect 358820 398210 358872 398216
rect 358820 398132 358872 398138
rect 358820 398074 358872 398080
rect 358832 397633 358860 398074
rect 358818 397624 358874 397633
rect 358818 397559 358874 397568
rect 358924 397254 358952 399758
rect 359062 399752 359090 400044
rect 359154 399906 359182 400044
rect 359246 399906 359274 400044
rect 359142 399900 359194 399906
rect 359142 399842 359194 399848
rect 359234 399900 359286 399906
rect 359234 399842 359286 399848
rect 359338 399752 359366 400044
rect 359430 399820 359458 400044
rect 359522 399945 359550 400044
rect 359508 399936 359564 399945
rect 359508 399871 359564 399880
rect 359614 399820 359642 400044
rect 359706 399838 359734 400044
rect 359430 399792 359504 399820
rect 359062 399724 359136 399752
rect 359338 399724 359412 399752
rect 359004 399628 359056 399634
rect 359004 399570 359056 399576
rect 359016 399265 359044 399570
rect 359002 399256 359058 399265
rect 359002 399191 359058 399200
rect 359004 398948 359056 398954
rect 359004 398890 359056 398896
rect 358912 397248 358964 397254
rect 358912 397190 358964 397196
rect 359016 395298 359044 398890
rect 359108 396098 359136 399724
rect 359280 399628 359332 399634
rect 359280 399570 359332 399576
rect 359188 399560 359240 399566
rect 359186 399528 359188 399537
rect 359240 399528 359242 399537
rect 359186 399463 359242 399472
rect 359292 397032 359320 399570
rect 359384 397866 359412 399724
rect 359372 397860 359424 397866
rect 359372 397802 359424 397808
rect 359476 397322 359504 399792
rect 359568 399792 359642 399820
rect 359694 399832 359746 399838
rect 359568 399752 359596 399792
rect 359798 399809 359826 400044
rect 359890 399906 359918 400044
rect 359982 399906 360010 400044
rect 360074 399945 360102 400044
rect 360060 399936 360116 399945
rect 359878 399900 359930 399906
rect 359878 399842 359930 399848
rect 359970 399900 360022 399906
rect 360060 399871 360116 399880
rect 359970 399842 360022 399848
rect 359694 399774 359746 399780
rect 359784 399800 359840 399809
rect 359568 399724 359642 399752
rect 359784 399735 359840 399744
rect 360016 399764 360068 399770
rect 359614 399616 359642 399724
rect 360166 399752 360194 400044
rect 360258 399906 360286 400044
rect 360350 399906 360378 400044
rect 360442 399906 360470 400044
rect 360534 399906 360562 400044
rect 360246 399900 360298 399906
rect 360246 399842 360298 399848
rect 360338 399900 360390 399906
rect 360338 399842 360390 399848
rect 360430 399900 360482 399906
rect 360430 399842 360482 399848
rect 360522 399900 360574 399906
rect 360522 399842 360574 399848
rect 360016 399706 360068 399712
rect 360120 399724 360194 399752
rect 359568 399588 359642 399616
rect 359740 399628 359792 399634
rect 359568 399430 359596 399588
rect 359740 399570 359792 399576
rect 359648 399492 359700 399498
rect 359648 399434 359700 399440
rect 359556 399424 359608 399430
rect 359556 399366 359608 399372
rect 359556 399220 359608 399226
rect 359556 399162 359608 399168
rect 359568 398954 359596 399162
rect 359556 398948 359608 398954
rect 359556 398890 359608 398896
rect 359464 397316 359516 397322
rect 359464 397258 359516 397264
rect 359292 397004 359412 397032
rect 359278 396536 359334 396545
rect 359278 396471 359334 396480
rect 359096 396092 359148 396098
rect 359096 396034 359148 396040
rect 359016 395270 359228 395298
rect 359002 395040 359058 395049
rect 359002 394975 359058 394984
rect 359016 377602 359044 394975
rect 359096 392692 359148 392698
rect 359096 392634 359148 392640
rect 359108 383518 359136 392634
rect 359096 383512 359148 383518
rect 359096 383454 359148 383460
rect 359004 377596 359056 377602
rect 359004 377538 359056 377544
rect 358728 312860 358780 312866
rect 358728 312802 358780 312808
rect 359200 306338 359228 395270
rect 359188 306332 359240 306338
rect 359188 306274 359240 306280
rect 358452 302116 358504 302122
rect 358452 302058 358504 302064
rect 359292 301986 359320 396471
rect 359384 303414 359412 397004
rect 359464 396772 359516 396778
rect 359464 396714 359516 396720
rect 359476 318306 359504 396714
rect 359556 394120 359608 394126
rect 359556 394062 359608 394068
rect 359568 393786 359596 394062
rect 359556 393780 359608 393786
rect 359556 393722 359608 393728
rect 359660 393650 359688 399434
rect 359752 399022 359780 399570
rect 359924 399560 359976 399566
rect 359924 399502 359976 399508
rect 359740 399016 359792 399022
rect 359740 398958 359792 398964
rect 359740 396500 359792 396506
rect 359740 396442 359792 396448
rect 359648 393644 359700 393650
rect 359648 393586 359700 393592
rect 359752 390554 359780 396442
rect 359936 393922 359964 399502
rect 359924 393916 359976 393922
rect 359924 393858 359976 393864
rect 360028 392698 360056 399706
rect 360120 396506 360148 399724
rect 360626 399684 360654 400044
rect 360718 399838 360746 400044
rect 360706 399832 360758 399838
rect 360706 399774 360758 399780
rect 360810 399684 360838 400044
rect 360902 399809 360930 400044
rect 360888 399800 360944 399809
rect 360888 399735 360944 399744
rect 360994 399752 361022 400044
rect 361086 399906 361114 400044
rect 361074 399900 361126 399906
rect 361074 399842 361126 399848
rect 361178 399752 361206 400044
rect 361270 399906 361298 400044
rect 361362 399906 361390 400044
rect 361454 399906 361482 400044
rect 361546 399945 361574 400044
rect 361532 399936 361588 399945
rect 361258 399900 361310 399906
rect 361258 399842 361310 399848
rect 361350 399900 361402 399906
rect 361350 399842 361402 399848
rect 361442 399900 361494 399906
rect 361638 399906 361666 400044
rect 361532 399871 361588 399880
rect 361626 399900 361678 399906
rect 361442 399842 361494 399848
rect 361626 399842 361678 399848
rect 361488 399764 361540 399770
rect 360994 399724 361068 399752
rect 361178 399724 361252 399752
rect 360580 399656 360654 399684
rect 360764 399656 360838 399684
rect 360200 399628 360252 399634
rect 360200 399570 360252 399576
rect 360212 397526 360240 399570
rect 360476 399560 360528 399566
rect 360476 399502 360528 399508
rect 360384 399492 360436 399498
rect 360384 399434 360436 399440
rect 360292 399356 360344 399362
rect 360292 399298 360344 399304
rect 360304 399022 360332 399298
rect 360292 399016 360344 399022
rect 360292 398958 360344 398964
rect 360200 397520 360252 397526
rect 360200 397462 360252 397468
rect 360292 396704 360344 396710
rect 360292 396646 360344 396652
rect 360108 396500 360160 396506
rect 360108 396442 360160 396448
rect 360016 392692 360068 392698
rect 360016 392634 360068 392640
rect 359660 390526 359780 390554
rect 359660 389174 359688 390526
rect 360304 389174 360332 396646
rect 359568 389146 359688 389174
rect 360212 389146 360332 389174
rect 359568 320958 359596 389146
rect 360212 383042 360240 389146
rect 360200 383036 360252 383042
rect 360200 382978 360252 382984
rect 359556 320952 359608 320958
rect 359556 320894 359608 320900
rect 359464 318300 359516 318306
rect 359464 318242 359516 318248
rect 360200 316736 360252 316742
rect 360200 316678 360252 316684
rect 360212 316130 360240 316678
rect 360200 316124 360252 316130
rect 360200 316066 360252 316072
rect 359372 303408 359424 303414
rect 359372 303350 359424 303356
rect 359280 301980 359332 301986
rect 359280 301922 359332 301928
rect 352564 301776 352616 301782
rect 352564 301718 352616 301724
rect 357440 258120 357492 258126
rect 357440 258062 357492 258068
rect 351460 251864 351512 251870
rect 351460 251806 351512 251812
rect 356060 145648 356112 145654
rect 356060 145590 356112 145596
rect 351920 136060 351972 136066
rect 351920 136002 351972 136008
rect 351932 16574 351960 136002
rect 354678 64152 354734 64161
rect 354678 64087 354734 64096
rect 354692 16574 354720 64087
rect 356072 16574 356100 145590
rect 357452 16574 357480 258062
rect 359464 145716 359516 145722
rect 359464 145658 359516 145664
rect 351932 16546 352880 16574
rect 354692 16546 355272 16574
rect 356072 16546 356376 16574
rect 357452 16546 357572 16574
rect 351642 3768 351698 3777
rect 351642 3703 351698 3712
rect 349252 3392 349304 3398
rect 349252 3334 349304 3340
rect 350448 3392 350500 3398
rect 350448 3334 350500 3340
rect 349172 1958 349292 1986
rect 349264 480 349292 1958
rect 350460 480 350488 3334
rect 351656 480 351684 3703
rect 352852 480 352880 16546
rect 354034 3768 354090 3777
rect 354034 3703 354090 3712
rect 354048 480 354076 3703
rect 355244 480 355272 16546
rect 356348 480 356376 16546
rect 357544 480 357572 16546
rect 358726 9480 358782 9489
rect 358726 9415 358782 9424
rect 358740 480 358768 9415
rect 359476 3398 359504 145658
rect 360212 16574 360240 316066
rect 360396 303278 360424 399434
rect 360488 398818 360516 399502
rect 360476 398812 360528 398818
rect 360476 398754 360528 398760
rect 360476 397248 360528 397254
rect 360476 397190 360528 397196
rect 360488 383178 360516 397190
rect 360580 396692 360608 399656
rect 360660 398744 360712 398750
rect 360660 398686 360712 398692
rect 360672 398342 360700 398686
rect 360660 398336 360712 398342
rect 360660 398278 360712 398284
rect 360764 397458 360792 399656
rect 361040 399294 361068 399724
rect 361120 399628 361172 399634
rect 361120 399570 361172 399576
rect 361028 399288 361080 399294
rect 361028 399230 361080 399236
rect 360844 398812 360896 398818
rect 360844 398754 360896 398760
rect 360752 397452 360804 397458
rect 360752 397394 360804 397400
rect 360580 396664 360792 396692
rect 360568 396568 360620 396574
rect 360568 396510 360620 396516
rect 360580 388686 360608 396510
rect 360660 390788 360712 390794
rect 360660 390730 360712 390736
rect 360568 388680 360620 388686
rect 360568 388622 360620 388628
rect 360476 383172 360528 383178
rect 360476 383114 360528 383120
rect 360672 307698 360700 390730
rect 360660 307692 360712 307698
rect 360660 307634 360712 307640
rect 360384 303272 360436 303278
rect 360384 303214 360436 303220
rect 360764 302054 360792 396664
rect 360856 395758 360884 398754
rect 361132 396692 361160 399570
rect 361224 397254 361252 399724
rect 361730 399752 361758 400044
rect 361822 399906 361850 400044
rect 361810 399900 361862 399906
rect 361810 399842 361862 399848
rect 361914 399786 361942 400044
rect 362006 399945 362034 400044
rect 361992 399936 362048 399945
rect 361992 399871 362048 399880
rect 362098 399820 362126 400044
rect 361488 399706 361540 399712
rect 361684 399724 361758 399752
rect 361868 399758 361942 399786
rect 362052 399792 362126 399820
rect 361396 399696 361448 399702
rect 361396 399638 361448 399644
rect 361304 399560 361356 399566
rect 361304 399502 361356 399508
rect 361212 397248 361264 397254
rect 361212 397190 361264 397196
rect 361132 396664 361252 396692
rect 360844 395752 360896 395758
rect 360844 395694 360896 395700
rect 361120 395412 361172 395418
rect 361120 395354 361172 395360
rect 360844 393780 360896 393786
rect 360844 393722 360896 393728
rect 360856 308718 360884 393722
rect 361132 389174 361160 395354
rect 360948 389146 361160 389174
rect 360948 318238 360976 389146
rect 361224 388482 361252 396664
rect 361316 390794 361344 399502
rect 361408 396574 361436 399638
rect 361500 398857 361528 399706
rect 361580 399696 361632 399702
rect 361580 399638 361632 399644
rect 361486 398848 361542 398857
rect 361486 398783 361542 398792
rect 361488 398744 361540 398750
rect 361488 398686 361540 398692
rect 361500 397769 361528 398686
rect 361486 397760 361542 397769
rect 361486 397695 361542 397704
rect 361592 396710 361620 399638
rect 361580 396704 361632 396710
rect 361580 396646 361632 396652
rect 361396 396568 361448 396574
rect 361684 396522 361712 399724
rect 361764 399628 361816 399634
rect 361764 399570 361816 399576
rect 361396 396510 361448 396516
rect 361592 396494 361712 396522
rect 361592 392834 361620 396494
rect 361672 396432 361724 396438
rect 361672 396374 361724 396380
rect 361580 392828 361632 392834
rect 361580 392770 361632 392776
rect 361304 390788 361356 390794
rect 361304 390730 361356 390736
rect 361212 388476 361264 388482
rect 361212 388418 361264 388424
rect 360936 318232 360988 318238
rect 360936 318174 360988 318180
rect 361396 316124 361448 316130
rect 361396 316066 361448 316072
rect 361408 315994 361436 316066
rect 361396 315988 361448 315994
rect 361396 315930 361448 315936
rect 361684 311506 361712 396374
rect 361776 319530 361804 399570
rect 361868 383246 361896 399758
rect 362052 397798 362080 399792
rect 362190 399752 362218 400044
rect 362144 399724 362218 399752
rect 362040 397792 362092 397798
rect 362040 397734 362092 397740
rect 362040 396704 362092 396710
rect 362040 396646 362092 396652
rect 361856 383240 361908 383246
rect 361856 383182 361908 383188
rect 361764 319524 361816 319530
rect 361764 319466 361816 319472
rect 361672 311500 361724 311506
rect 361672 311442 361724 311448
rect 360844 308712 360896 308718
rect 360844 308654 360896 308660
rect 360752 302048 360804 302054
rect 360752 301990 360804 301996
rect 362052 300422 362080 396646
rect 362144 395146 362172 399724
rect 362282 399650 362310 400044
rect 362374 399752 362402 400044
rect 362466 399906 362494 400044
rect 362454 399900 362506 399906
rect 362454 399842 362506 399848
rect 362558 399752 362586 400044
rect 362374 399724 362448 399752
rect 362282 399622 362356 399650
rect 362328 398546 362356 399622
rect 362420 398614 362448 399724
rect 362512 399724 362586 399752
rect 362408 398608 362460 398614
rect 362408 398550 362460 398556
rect 362316 398540 362368 398546
rect 362316 398482 362368 398488
rect 362224 398268 362276 398274
rect 362224 398210 362276 398216
rect 362132 395140 362184 395146
rect 362132 395082 362184 395088
rect 362236 311370 362264 398210
rect 362512 396710 362540 399724
rect 362650 399684 362678 400044
rect 362742 399838 362770 400044
rect 362834 399906 362862 400044
rect 362926 399906 362954 400044
rect 363018 399906 363046 400044
rect 362822 399900 362874 399906
rect 362822 399842 362874 399848
rect 362914 399900 362966 399906
rect 362914 399842 362966 399848
rect 363006 399900 363058 399906
rect 363006 399842 363058 399848
rect 362730 399832 362782 399838
rect 363110 399786 363138 400044
rect 363202 399838 363230 400044
rect 363294 399945 363322 400044
rect 363280 399936 363336 399945
rect 363280 399871 363336 399880
rect 362730 399774 362782 399780
rect 362960 399764 363012 399770
rect 362960 399706 363012 399712
rect 363064 399758 363138 399786
rect 363190 399832 363242 399838
rect 363190 399774 363242 399780
rect 362868 399696 362920 399702
rect 362650 399656 362724 399684
rect 362592 399560 362644 399566
rect 362592 399502 362644 399508
rect 362500 396704 362552 396710
rect 362500 396646 362552 396652
rect 362604 396438 362632 399502
rect 362696 396778 362724 399656
rect 362788 399656 362868 399684
rect 362684 396772 362736 396778
rect 362684 396714 362736 396720
rect 362592 396432 362644 396438
rect 362592 396374 362644 396380
rect 362788 393145 362816 399656
rect 362868 399638 362920 399644
rect 362972 399158 363000 399706
rect 363064 399362 363092 399758
rect 363144 399696 363196 399702
rect 363386 399684 363414 400044
rect 363478 399838 363506 400044
rect 363570 399906 363598 400044
rect 363662 399945 363690 400044
rect 363648 399936 363704 399945
rect 363558 399900 363610 399906
rect 363754 399906 363782 400044
rect 363648 399871 363704 399880
rect 363742 399900 363794 399906
rect 363558 399842 363610 399848
rect 363742 399842 363794 399848
rect 363846 399838 363874 400044
rect 363938 399906 363966 400044
rect 363926 399900 363978 399906
rect 363926 399842 363978 399848
rect 363466 399832 363518 399838
rect 363466 399774 363518 399780
rect 363834 399832 363886 399838
rect 364030 399786 364058 400044
rect 364122 399906 364150 400044
rect 364214 399945 364242 400044
rect 364200 399936 364256 399945
rect 364110 399900 364162 399906
rect 364306 399906 364334 400044
rect 364398 399906 364426 400044
rect 364200 399871 364256 399880
rect 364294 399900 364346 399906
rect 364110 399842 364162 399848
rect 364294 399842 364346 399848
rect 364386 399900 364438 399906
rect 364386 399842 364438 399848
rect 363834 399774 363886 399780
rect 363696 399764 363748 399770
rect 363696 399706 363748 399712
rect 363984 399758 364058 399786
rect 364156 399764 364208 399770
rect 363604 399696 363656 399702
rect 363144 399638 363196 399644
rect 363340 399656 363414 399684
rect 363524 399656 363604 399684
rect 363052 399356 363104 399362
rect 363052 399298 363104 399304
rect 362960 399152 363012 399158
rect 362960 399094 363012 399100
rect 362868 398608 362920 398614
rect 362868 398550 362920 398556
rect 362880 398041 362908 398550
rect 362866 398032 362922 398041
rect 362866 397967 362922 397976
rect 362868 397860 362920 397866
rect 362868 397802 362920 397808
rect 362880 396030 362908 397802
rect 362868 396024 362920 396030
rect 362868 395966 362920 395972
rect 363156 394694 363184 399638
rect 363236 399628 363288 399634
rect 363236 399570 363288 399576
rect 363064 394666 363184 394694
rect 363248 394670 363276 399570
rect 362774 393136 362830 393145
rect 362774 393071 362830 393080
rect 363064 392630 363092 394666
rect 363236 394664 363288 394670
rect 363236 394606 363288 394612
rect 363340 394602 363368 399656
rect 363420 399356 363472 399362
rect 363420 399298 363472 399304
rect 363144 394596 363196 394602
rect 363144 394538 363196 394544
rect 363328 394596 363380 394602
rect 363328 394538 363380 394544
rect 363156 392766 363184 394538
rect 363234 394496 363290 394505
rect 363234 394431 363290 394440
rect 363144 392760 363196 392766
rect 363144 392702 363196 392708
rect 363052 392624 363104 392630
rect 363052 392566 363104 392572
rect 363248 377534 363276 394431
rect 363236 377528 363288 377534
rect 363236 377470 363288 377476
rect 362224 311364 362276 311370
rect 362224 311306 362276 311312
rect 362040 300416 362092 300422
rect 362040 300358 362092 300364
rect 363432 297634 363460 399298
rect 363524 393854 363552 399656
rect 363604 399638 363656 399644
rect 363604 399560 363656 399566
rect 363604 399502 363656 399508
rect 363616 396642 363644 399502
rect 363708 397730 363736 399706
rect 363880 399628 363932 399634
rect 363880 399570 363932 399576
rect 363788 399492 363840 399498
rect 363788 399434 363840 399440
rect 363696 397724 363748 397730
rect 363696 397666 363748 397672
rect 363604 396636 363656 396642
rect 363604 396578 363656 396584
rect 363696 396364 363748 396370
rect 363696 396306 363748 396312
rect 363512 393848 363564 393854
rect 363708 393802 363736 396306
rect 363512 393790 363564 393796
rect 363616 393774 363736 393802
rect 363512 393508 363564 393514
rect 363512 393450 363564 393456
rect 363524 385830 363552 393450
rect 363512 385824 363564 385830
rect 363512 385766 363564 385772
rect 363616 308854 363644 393774
rect 363696 393712 363748 393718
rect 363696 393654 363748 393660
rect 363708 322318 363736 393654
rect 363696 322312 363748 322318
rect 363696 322254 363748 322260
rect 363604 308848 363656 308854
rect 363604 308790 363656 308796
rect 363800 307630 363828 399434
rect 363892 314158 363920 399570
rect 363984 393514 364012 399758
rect 364490 399752 364518 400044
rect 364582 399906 364610 400044
rect 364570 399900 364622 399906
rect 364570 399842 364622 399848
rect 364490 399724 364564 399752
rect 364156 399706 364208 399712
rect 364168 399537 364196 399706
rect 364340 399560 364392 399566
rect 364154 399528 364210 399537
rect 364064 399492 364116 399498
rect 364340 399502 364392 399508
rect 364432 399560 364484 399566
rect 364432 399502 364484 399508
rect 364154 399463 364210 399472
rect 364064 399434 364116 399440
rect 364076 395593 364104 399434
rect 364248 399152 364300 399158
rect 364248 399094 364300 399100
rect 364260 398954 364288 399094
rect 364248 398948 364300 398954
rect 364248 398890 364300 398896
rect 364156 397724 364208 397730
rect 364156 397666 364208 397672
rect 364062 395584 364118 395593
rect 364062 395519 364118 395528
rect 364168 393718 364196 397666
rect 364248 396636 364300 396642
rect 364248 396578 364300 396584
rect 364156 393712 364208 393718
rect 364156 393654 364208 393660
rect 363972 393508 364024 393514
rect 363972 393450 364024 393456
rect 364260 393038 364288 396578
rect 364248 393032 364300 393038
rect 364248 392974 364300 392980
rect 364352 392737 364380 399502
rect 364444 397186 364472 399502
rect 364432 397180 364484 397186
rect 364432 397122 364484 397128
rect 364536 395321 364564 399724
rect 364674 399650 364702 400044
rect 364766 399945 364794 400044
rect 364752 399936 364808 399945
rect 364858 399906 364886 400044
rect 364752 399871 364808 399880
rect 364846 399900 364898 399906
rect 364846 399842 364898 399848
rect 364950 399786 364978 400044
rect 364904 399758 364978 399786
rect 364800 399696 364852 399702
rect 364674 399622 364748 399650
rect 364800 399638 364852 399644
rect 364616 399560 364668 399566
rect 364616 399502 364668 399508
rect 364522 395312 364578 395321
rect 364522 395247 364578 395256
rect 364522 395040 364578 395049
rect 364522 394975 364578 394984
rect 364338 392728 364394 392737
rect 364338 392663 364394 392672
rect 364536 318170 364564 394975
rect 364628 373561 364656 399502
rect 364720 395185 364748 399622
rect 364706 395176 364762 395185
rect 364706 395111 364762 395120
rect 364708 394664 364760 394670
rect 364708 394606 364760 394612
rect 364614 373552 364670 373561
rect 364614 373487 364670 373496
rect 364524 318164 364576 318170
rect 364524 318106 364576 318112
rect 363880 314152 363932 314158
rect 363880 314094 363932 314100
rect 363788 307624 363840 307630
rect 363788 307566 363840 307572
rect 364720 303482 364748 394606
rect 364812 390554 364840 399638
rect 364904 395962 364932 399758
rect 365042 399684 365070 400044
rect 365134 399809 365162 400044
rect 365226 399838 365254 400044
rect 365318 399945 365346 400044
rect 365304 399936 365360 399945
rect 365304 399871 365360 399880
rect 365410 399838 365438 400044
rect 365214 399832 365266 399838
rect 365120 399800 365176 399809
rect 365214 399774 365266 399780
rect 365398 399832 365450 399838
rect 365398 399774 365450 399780
rect 365120 399735 365176 399744
rect 365502 399752 365530 400044
rect 365594 399906 365622 400044
rect 365686 399906 365714 400044
rect 365778 399906 365806 400044
rect 365582 399900 365634 399906
rect 365582 399842 365634 399848
rect 365674 399900 365726 399906
rect 365674 399842 365726 399848
rect 365766 399900 365818 399906
rect 365766 399842 365818 399848
rect 365870 399838 365898 400044
rect 365962 399838 365990 400044
rect 365858 399832 365910 399838
rect 365858 399774 365910 399780
rect 365950 399832 366002 399838
rect 366054 399809 366082 400044
rect 365950 399774 366002 399780
rect 366040 399800 366096 399809
rect 365502 399724 365576 399752
rect 366146 399786 366174 400044
rect 366238 399906 366266 400044
rect 366226 399900 366278 399906
rect 366226 399842 366278 399848
rect 366330 399786 366358 400044
rect 366422 399906 366450 400044
rect 366410 399900 366462 399906
rect 366410 399842 366462 399848
rect 366146 399758 366266 399786
rect 366330 399758 366404 399786
rect 366040 399735 366096 399744
rect 365260 399696 365312 399702
rect 365042 399656 365116 399684
rect 365088 399537 365116 399656
rect 365260 399638 365312 399644
rect 365168 399560 365220 399566
rect 365074 399528 365130 399537
rect 365168 399502 365220 399508
rect 365074 399463 365130 399472
rect 364984 397384 365036 397390
rect 364984 397326 365036 397332
rect 364892 395956 364944 395962
rect 364892 395898 364944 395904
rect 364812 390526 364932 390554
rect 364904 308446 364932 390526
rect 364892 308440 364944 308446
rect 364892 308382 364944 308388
rect 364708 303476 364760 303482
rect 364708 303418 364760 303424
rect 364996 297702 365024 397326
rect 365180 396001 365208 399502
rect 365166 395992 365222 396001
rect 365166 395927 365222 395936
rect 365272 390554 365300 399638
rect 365352 399560 365404 399566
rect 365352 399502 365404 399508
rect 365364 396370 365392 399502
rect 365352 396364 365404 396370
rect 365352 396306 365404 396312
rect 365548 391746 365576 399724
rect 365812 399696 365864 399702
rect 365812 399638 365864 399644
rect 365904 399696 365956 399702
rect 365904 399638 365956 399644
rect 366088 399696 366140 399702
rect 366238 399684 366266 399758
rect 366238 399656 366312 399684
rect 366088 399638 366140 399644
rect 365720 399628 365772 399634
rect 365720 399570 365772 399576
rect 365732 399242 365760 399570
rect 365640 399214 365760 399242
rect 365640 393786 365668 399214
rect 365824 397866 365852 399638
rect 365812 397860 365864 397866
rect 365812 397802 365864 397808
rect 365812 397588 365864 397594
rect 365812 397530 365864 397536
rect 365720 395140 365772 395146
rect 365720 395082 365772 395088
rect 365628 393780 365680 393786
rect 365628 393722 365680 393728
rect 365536 391740 365588 391746
rect 365536 391682 365588 391688
rect 365180 390526 365300 390554
rect 365180 313002 365208 390526
rect 365168 312996 365220 313002
rect 365168 312938 365220 312944
rect 365732 303550 365760 395082
rect 365824 308786 365852 397530
rect 365916 393990 365944 399638
rect 365996 399424 366048 399430
rect 365996 399366 366048 399372
rect 365904 393984 365956 393990
rect 365904 393926 365956 393932
rect 366008 389174 366036 399366
rect 365916 389146 366036 389174
rect 365916 385694 365944 389146
rect 365904 385688 365956 385694
rect 365904 385630 365956 385636
rect 365812 308780 365864 308786
rect 365812 308722 365864 308728
rect 365720 303544 365772 303550
rect 365720 303486 365772 303492
rect 366100 298110 366128 399638
rect 366180 399560 366232 399566
rect 366180 399502 366232 399508
rect 366192 389910 366220 399502
rect 366284 397390 366312 399656
rect 366272 397384 366324 397390
rect 366376 397361 366404 399758
rect 366514 399752 366542 400044
rect 366468 399724 366542 399752
rect 366468 397390 366496 399724
rect 366606 399684 366634 400044
rect 366698 399906 366726 400044
rect 366790 399906 366818 400044
rect 366882 399906 366910 400044
rect 366686 399900 366738 399906
rect 366686 399842 366738 399848
rect 366778 399900 366830 399906
rect 366778 399842 366830 399848
rect 366870 399900 366922 399906
rect 366870 399842 366922 399848
rect 366974 399752 367002 400044
rect 367066 399906 367094 400044
rect 367054 399900 367106 399906
rect 367054 399842 367106 399848
rect 367158 399752 367186 400044
rect 367250 399945 367278 400044
rect 367236 399936 367292 399945
rect 367236 399871 367292 399880
rect 367342 399786 367370 400044
rect 367434 399906 367462 400044
rect 367422 399900 367474 399906
rect 367422 399842 367474 399848
rect 367526 399838 367554 400044
rect 367618 399945 367646 400044
rect 367604 399936 367660 399945
rect 367604 399871 367660 399880
rect 366560 399656 366634 399684
rect 366928 399724 367002 399752
rect 367112 399724 367186 399752
rect 367296 399758 367370 399786
rect 367514 399832 367566 399838
rect 367710 399820 367738 400044
rect 367802 399906 367830 400044
rect 367790 399900 367842 399906
rect 367790 399842 367842 399848
rect 367514 399774 367566 399780
rect 367664 399792 367738 399820
rect 366560 398818 366588 399656
rect 366824 399628 366876 399634
rect 366824 399570 366876 399576
rect 366640 399492 366692 399498
rect 366640 399434 366692 399440
rect 366548 398812 366600 398818
rect 366548 398754 366600 398760
rect 366546 398712 366602 398721
rect 366546 398647 366548 398656
rect 366600 398647 366602 398656
rect 366548 398618 366600 398624
rect 366548 397656 366600 397662
rect 366548 397598 366600 397604
rect 366456 397384 366508 397390
rect 366272 397326 366324 397332
rect 366362 397352 366418 397361
rect 366456 397326 366508 397332
rect 366362 397287 366418 397296
rect 366456 394732 366508 394738
rect 366456 394674 366508 394680
rect 366272 393984 366324 393990
rect 366272 393926 366324 393932
rect 366180 389904 366232 389910
rect 366180 389846 366232 389852
rect 366284 383217 366312 393926
rect 366270 383208 366326 383217
rect 366270 383143 366326 383152
rect 366468 308922 366496 394674
rect 366560 315994 366588 397598
rect 366652 397361 366680 399434
rect 366732 397384 366784 397390
rect 366638 397352 366694 397361
rect 366732 397326 366784 397332
rect 366638 397287 366694 397296
rect 366744 394330 366772 397326
rect 366836 397050 366864 399570
rect 366824 397044 366876 397050
rect 366824 396986 366876 396992
rect 366732 394324 366784 394330
rect 366732 394266 366784 394272
rect 366928 393718 366956 399724
rect 367112 399650 367140 399724
rect 367020 399622 367140 399650
rect 367192 399628 367244 399634
rect 367020 397390 367048 399622
rect 367192 399570 367244 399576
rect 367100 399560 367152 399566
rect 367100 399502 367152 399508
rect 367008 397384 367060 397390
rect 367008 397326 367060 397332
rect 367112 394738 367140 399502
rect 367204 397361 367232 399570
rect 367190 397352 367246 397361
rect 367190 397287 367246 397296
rect 367190 395992 367246 396001
rect 367190 395927 367246 395936
rect 367100 394732 367152 394738
rect 367100 394674 367152 394680
rect 366916 393712 366968 393718
rect 366916 393654 366968 393660
rect 367204 393650 367232 395927
rect 367296 393990 367324 399758
rect 367376 399696 367428 399702
rect 367376 399638 367428 399644
rect 367468 399696 367520 399702
rect 367468 399638 367520 399644
rect 367284 393984 367336 393990
rect 367284 393926 367336 393932
rect 367388 393802 367416 399638
rect 367480 398177 367508 399638
rect 367466 398168 367522 398177
rect 367466 398103 367522 398112
rect 367664 395350 367692 399792
rect 367894 399752 367922 400044
rect 367986 399906 368014 400044
rect 367974 399900 368026 399906
rect 367974 399842 368026 399848
rect 368078 399838 368106 400044
rect 368170 399838 368198 400044
rect 368066 399832 368118 399838
rect 368066 399774 368118 399780
rect 368158 399832 368210 399838
rect 368158 399774 368210 399780
rect 367848 399724 367922 399752
rect 367744 399696 367796 399702
rect 367744 399638 367796 399644
rect 367652 395344 367704 395350
rect 367652 395286 367704 395292
rect 367388 393774 367692 393802
rect 367468 393712 367520 393718
rect 367468 393654 367520 393660
rect 367192 393644 367244 393650
rect 367192 393586 367244 393592
rect 367376 392556 367428 392562
rect 367376 392498 367428 392504
rect 367388 377466 367416 392498
rect 367376 377460 367428 377466
rect 367376 377402 367428 377408
rect 366548 315988 366600 315994
rect 366548 315930 366600 315936
rect 366456 308916 366508 308922
rect 366456 308858 366508 308864
rect 366088 298104 366140 298110
rect 366088 298046 366140 298052
rect 367480 297770 367508 393654
rect 367560 393644 367612 393650
rect 367560 393586 367612 393592
rect 367572 300830 367600 393586
rect 367560 300824 367612 300830
rect 367560 300766 367612 300772
rect 367664 300558 367692 393774
rect 367756 392562 367784 399638
rect 367848 398041 367876 399724
rect 368020 399696 368072 399702
rect 368020 399638 368072 399644
rect 368032 399208 368060 399638
rect 368112 399628 368164 399634
rect 368262 399616 368290 400044
rect 368354 399906 368382 400044
rect 368342 399900 368394 399906
rect 368342 399842 368394 399848
rect 368446 399838 368474 400044
rect 368538 399838 368566 400044
rect 368630 399906 368658 400044
rect 368722 399945 368750 400044
rect 368708 399936 368764 399945
rect 368618 399900 368670 399906
rect 368708 399871 368764 399880
rect 368618 399842 368670 399848
rect 368434 399832 368486 399838
rect 368434 399774 368486 399780
rect 368526 399832 368578 399838
rect 368814 399786 368842 400044
rect 368526 399774 368578 399780
rect 368112 399570 368164 399576
rect 368216 399588 368290 399616
rect 368768 399758 368842 399786
rect 367940 399180 368060 399208
rect 367834 398032 367890 398041
rect 367834 397967 367890 397976
rect 367836 397928 367888 397934
rect 367836 397870 367888 397876
rect 367744 392556 367796 392562
rect 367744 392498 367796 392504
rect 367848 389174 367876 397870
rect 367940 394262 367968 399180
rect 368124 399140 368152 399570
rect 368032 399112 368152 399140
rect 368032 395690 368060 399112
rect 368216 399072 368244 399588
rect 368572 399560 368624 399566
rect 368572 399502 368624 399508
rect 368296 399492 368348 399498
rect 368296 399434 368348 399440
rect 368480 399492 368532 399498
rect 368480 399434 368532 399440
rect 368124 399044 368244 399072
rect 368124 396982 368152 399044
rect 368308 398120 368336 399434
rect 368216 398092 368336 398120
rect 368112 396976 368164 396982
rect 368112 396918 368164 396924
rect 368020 395684 368072 395690
rect 368020 395626 368072 395632
rect 367928 394256 367980 394262
rect 367928 394198 367980 394204
rect 367928 393984 367980 393990
rect 367928 393926 367980 393932
rect 367756 389146 367876 389174
rect 367756 383450 367784 389146
rect 367744 383444 367796 383450
rect 367744 383386 367796 383392
rect 367940 308310 367968 393926
rect 368216 391950 368244 398092
rect 368294 398032 368350 398041
rect 368294 397967 368350 397976
rect 368204 391944 368256 391950
rect 368204 391886 368256 391892
rect 368308 308990 368336 397967
rect 368492 392850 368520 399434
rect 368584 393990 368612 399502
rect 368664 399492 368716 399498
rect 368664 399434 368716 399440
rect 368676 398585 368704 399434
rect 368662 398576 368718 398585
rect 368662 398511 368718 398520
rect 368768 397984 368796 399758
rect 368906 399752 368934 400044
rect 368998 399906 369026 400044
rect 368986 399900 369038 399906
rect 368986 399842 369038 399848
rect 369090 399752 369118 400044
rect 369182 399945 369210 400044
rect 369168 399936 369224 399945
rect 369168 399871 369224 399880
rect 369274 399786 369302 400044
rect 369228 399770 369302 399786
rect 368906 399724 368980 399752
rect 368848 399628 368900 399634
rect 368848 399570 368900 399576
rect 368676 397956 368796 397984
rect 368676 397730 368704 397956
rect 368754 397896 368810 397905
rect 368754 397831 368810 397840
rect 368664 397724 368716 397730
rect 368664 397666 368716 397672
rect 368572 393984 368624 393990
rect 368572 393926 368624 393932
rect 368492 392822 368612 392850
rect 368478 392728 368534 392737
rect 368478 392663 368534 392672
rect 368492 392018 368520 392663
rect 368480 392012 368532 392018
rect 368480 391954 368532 391960
rect 368584 391610 368612 392822
rect 368768 392034 368796 397831
rect 368676 392006 368796 392034
rect 368572 391604 368624 391610
rect 368572 391546 368624 391552
rect 368676 321094 368704 392006
rect 368756 390788 368808 390794
rect 368756 390730 368808 390736
rect 368768 336054 368796 390730
rect 368860 377505 368888 399570
rect 368952 398886 368980 399724
rect 369044 399724 369118 399752
rect 369216 399764 369302 399770
rect 368940 398880 368992 398886
rect 368940 398822 368992 398828
rect 368940 398676 368992 398682
rect 368940 398618 368992 398624
rect 368846 377496 368902 377505
rect 368846 377431 368902 377440
rect 368756 336048 368808 336054
rect 368756 335990 368808 335996
rect 368664 321088 368716 321094
rect 368664 321030 368716 321036
rect 368296 308984 368348 308990
rect 368296 308926 368348 308932
rect 367928 308304 367980 308310
rect 367928 308246 367980 308252
rect 367652 300552 367704 300558
rect 367652 300494 367704 300500
rect 368952 298042 368980 398618
rect 369044 397934 369072 399724
rect 369268 399758 369302 399764
rect 369216 399706 369268 399712
rect 369366 399684 369394 400044
rect 369458 399906 369486 400044
rect 369550 399945 369578 400044
rect 369536 399936 369592 399945
rect 369446 399900 369498 399906
rect 369536 399871 369592 399880
rect 369446 399842 369498 399848
rect 369642 399752 369670 400044
rect 369734 399945 369762 400044
rect 369720 399936 369776 399945
rect 369720 399871 369776 399880
rect 369826 399838 369854 400044
rect 369918 399906 369946 400044
rect 370010 399906 370038 400044
rect 369906 399900 369958 399906
rect 369906 399842 369958 399848
rect 369998 399900 370050 399906
rect 369998 399842 370050 399848
rect 370102 399838 370130 400044
rect 370194 399906 370222 400044
rect 370182 399900 370234 399906
rect 370182 399842 370234 399848
rect 369814 399832 369866 399838
rect 369814 399774 369866 399780
rect 370090 399832 370142 399838
rect 370286 399809 370314 400044
rect 370378 399945 370406 400044
rect 370364 399936 370420 399945
rect 370364 399871 370420 399880
rect 370090 399774 370142 399780
rect 370272 399800 370328 399809
rect 369596 399724 369670 399752
rect 370470 399786 370498 400044
rect 370562 399838 370590 400044
rect 370654 399945 370682 400044
rect 370640 399936 370696 399945
rect 370640 399871 370696 399880
rect 370272 399735 370328 399744
rect 370424 399758 370498 399786
rect 370550 399832 370602 399838
rect 370746 399820 370774 400044
rect 370550 399774 370602 399780
rect 370700 399792 370774 399820
rect 369366 399656 369440 399684
rect 369124 399628 369176 399634
rect 369124 399570 369176 399576
rect 369032 397928 369084 397934
rect 369032 397870 369084 397876
rect 369136 397526 369164 399570
rect 369412 399514 369440 399656
rect 369412 399486 369532 399514
rect 369400 399424 369452 399430
rect 369400 399366 369452 399372
rect 369308 398880 369360 398886
rect 369308 398822 369360 398828
rect 369124 397520 369176 397526
rect 369124 397462 369176 397468
rect 369030 395720 369086 395729
rect 369030 395655 369086 395664
rect 369044 303618 369072 395655
rect 369124 393984 369176 393990
rect 369124 393926 369176 393932
rect 369032 303612 369084 303618
rect 369032 303554 369084 303560
rect 369136 298858 369164 393926
rect 369124 298852 369176 298858
rect 369124 298794 369176 298800
rect 368940 298036 368992 298042
rect 368940 297978 368992 297984
rect 369320 297838 369348 398822
rect 369412 391921 369440 399366
rect 369504 397458 369532 399486
rect 369492 397452 369544 397458
rect 369492 397394 369544 397400
rect 369398 391912 369454 391921
rect 369398 391847 369454 391856
rect 369596 390794 369624 399724
rect 369860 399628 369912 399634
rect 369860 399570 369912 399576
rect 369676 399492 369728 399498
rect 369676 399434 369728 399440
rect 369688 398274 369716 399434
rect 369872 399265 369900 399570
rect 369952 399560 370004 399566
rect 369952 399502 370004 399508
rect 370320 399560 370372 399566
rect 370320 399502 370372 399508
rect 369858 399256 369914 399265
rect 369858 399191 369914 399200
rect 369768 398540 369820 398546
rect 369768 398482 369820 398488
rect 369676 398268 369728 398274
rect 369676 398210 369728 398216
rect 369780 396074 369808 398482
rect 369860 397384 369912 397390
rect 369860 397326 369912 397332
rect 369688 396046 369808 396074
rect 369584 390788 369636 390794
rect 369584 390730 369636 390736
rect 369688 389174 369716 396046
rect 369872 389174 369900 397326
rect 369964 395418 369992 399502
rect 370136 399492 370188 399498
rect 370136 399434 370188 399440
rect 370042 398712 370098 398721
rect 370042 398647 370098 398656
rect 369952 395412 370004 395418
rect 369952 395354 370004 395360
rect 369688 389146 369808 389174
rect 369872 389146 369992 389174
rect 369780 385762 369808 389146
rect 369768 385756 369820 385762
rect 369768 385698 369820 385704
rect 369964 300694 369992 389146
rect 370056 388754 370084 398647
rect 370148 397118 370176 399434
rect 370228 399288 370280 399294
rect 370228 399230 370280 399236
rect 370240 398449 370268 399230
rect 370226 398440 370282 398449
rect 370226 398375 370282 398384
rect 370136 397112 370188 397118
rect 370136 397054 370188 397060
rect 370228 394052 370280 394058
rect 370228 393994 370280 394000
rect 370136 393984 370188 393990
rect 370136 393926 370188 393932
rect 370148 388958 370176 393926
rect 370136 388952 370188 388958
rect 370136 388894 370188 388900
rect 370240 388890 370268 393994
rect 370228 388884 370280 388890
rect 370228 388826 370280 388832
rect 370044 388748 370096 388754
rect 370044 388690 370096 388696
rect 370332 312934 370360 399502
rect 370424 397662 370452 399758
rect 370596 399696 370648 399702
rect 370596 399638 370648 399644
rect 370504 399628 370556 399634
rect 370504 399570 370556 399576
rect 370516 399537 370544 399570
rect 370502 399528 370558 399537
rect 370502 399463 370558 399472
rect 370608 398585 370636 399638
rect 370700 399362 370728 399792
rect 370838 399752 370866 400044
rect 370792 399724 370866 399752
rect 370688 399356 370740 399362
rect 370688 399298 370740 399304
rect 370686 399256 370742 399265
rect 370686 399191 370742 399200
rect 370594 398576 370650 398585
rect 370594 398511 370650 398520
rect 370594 398440 370650 398449
rect 370594 398375 370650 398384
rect 370412 397656 370464 397662
rect 370412 397598 370464 397604
rect 370504 394732 370556 394738
rect 370504 394674 370556 394680
rect 370320 312928 370372 312934
rect 370320 312870 370372 312876
rect 370516 304706 370544 394674
rect 370608 393990 370636 398375
rect 370700 395894 370728 399191
rect 370792 397769 370820 399724
rect 370930 399684 370958 400044
rect 371022 399911 371050 400044
rect 371008 399902 371064 399911
rect 371008 399837 371064 399846
rect 371114 399786 371142 400044
rect 370884 399656 370958 399684
rect 371068 399758 371142 399786
rect 370778 397760 370834 397769
rect 370778 397695 370834 397704
rect 370780 397520 370832 397526
rect 370780 397462 370832 397468
rect 370688 395888 370740 395894
rect 370688 395830 370740 395836
rect 370596 393984 370648 393990
rect 370596 393926 370648 393932
rect 370686 393952 370742 393961
rect 370686 393887 370742 393896
rect 370596 393848 370648 393854
rect 370596 393790 370648 393796
rect 370608 307426 370636 393790
rect 370700 308825 370728 393887
rect 370792 393854 370820 397462
rect 370884 394058 370912 399656
rect 370964 399356 371016 399362
rect 370964 399298 371016 399304
rect 370976 395826 371004 399298
rect 371068 397905 371096 399758
rect 371206 399650 371234 400044
rect 371298 399752 371326 400044
rect 371390 399906 371418 400044
rect 371482 399945 371510 400044
rect 371468 399936 371524 399945
rect 371378 399900 371430 399906
rect 371468 399871 371524 399880
rect 371378 399842 371430 399848
rect 371298 399724 371372 399752
rect 371206 399622 371280 399650
rect 371146 399528 371202 399537
rect 371146 399463 371202 399472
rect 371160 398410 371188 399463
rect 371148 398404 371200 398410
rect 371148 398346 371200 398352
rect 371054 397896 371110 397905
rect 371054 397831 371110 397840
rect 370964 395820 371016 395826
rect 370964 395762 371016 395768
rect 371252 394738 371280 399622
rect 371344 399378 371372 399724
rect 371574 399684 371602 400044
rect 371666 399945 371694 400044
rect 371652 399936 371708 399945
rect 371652 399871 371708 399880
rect 371758 399820 371786 400044
rect 371712 399792 371786 399820
rect 371574 399656 371648 399684
rect 371344 399350 371464 399378
rect 371330 399256 371386 399265
rect 371330 399191 371386 399200
rect 371240 394732 371292 394738
rect 371240 394674 371292 394680
rect 371240 394256 371292 394262
rect 371240 394198 371292 394204
rect 370872 394052 370924 394058
rect 370872 393994 370924 394000
rect 370780 393848 370832 393854
rect 370780 393790 370832 393796
rect 371252 391406 371280 394198
rect 371240 391400 371292 391406
rect 371240 391342 371292 391348
rect 371344 391270 371372 399191
rect 371332 391264 371384 391270
rect 371332 391206 371384 391212
rect 371436 311778 371464 399350
rect 371516 399356 371568 399362
rect 371516 399298 371568 399304
rect 371528 394262 371556 399298
rect 371516 394256 371568 394262
rect 371516 394198 371568 394204
rect 371516 394052 371568 394058
rect 371516 393994 371568 394000
rect 371424 311772 371476 311778
rect 371424 311714 371476 311720
rect 371528 311302 371556 393994
rect 371620 313138 371648 399656
rect 371712 399362 371740 399792
rect 371850 399752 371878 400044
rect 371942 399906 371970 400044
rect 372034 399911 372062 400044
rect 371930 399900 371982 399906
rect 371930 399842 371982 399848
rect 372020 399902 372076 399911
rect 372020 399837 372076 399846
rect 372126 399786 372154 400044
rect 371804 399724 371878 399752
rect 371976 399764 372028 399770
rect 371700 399356 371752 399362
rect 371700 399298 371752 399304
rect 371698 399256 371754 399265
rect 371698 399191 371754 399200
rect 371712 319462 371740 399191
rect 371804 395350 371832 399724
rect 371976 399706 372028 399712
rect 372080 399758 372154 399786
rect 371988 399650 372016 399706
rect 371896 399622 372016 399650
rect 371792 395344 371844 395350
rect 371792 395286 371844 395292
rect 371896 394058 371924 399622
rect 371884 394052 371936 394058
rect 371884 393994 371936 394000
rect 371792 393984 371844 393990
rect 371792 393926 371844 393932
rect 371804 333266 371832 393926
rect 371792 333260 371844 333266
rect 371792 333202 371844 333208
rect 371700 319456 371752 319462
rect 371700 319398 371752 319404
rect 371608 313132 371660 313138
rect 371608 313074 371660 313080
rect 371516 311296 371568 311302
rect 371516 311238 371568 311244
rect 370686 308816 370742 308825
rect 370686 308751 370742 308760
rect 370596 307420 370648 307426
rect 370596 307362 370648 307368
rect 370504 304700 370556 304706
rect 370504 304642 370556 304648
rect 372080 301918 372108 399758
rect 372218 399650 372246 400044
rect 372310 399786 372338 400044
rect 372402 399906 372430 400044
rect 372390 399900 372442 399906
rect 372390 399842 372442 399848
rect 372494 399786 372522 400044
rect 372586 399906 372614 400044
rect 372678 399911 372706 400044
rect 372574 399900 372626 399906
rect 372574 399842 372626 399848
rect 372664 399902 372720 399911
rect 372664 399837 372720 399846
rect 372310 399758 372384 399786
rect 372172 399622 372246 399650
rect 372172 305862 372200 399622
rect 372252 399084 372304 399090
rect 372252 399026 372304 399032
rect 372264 398954 372292 399026
rect 372252 398948 372304 398954
rect 372252 398890 372304 398896
rect 372250 398712 372306 398721
rect 372250 398647 372306 398656
rect 372264 398274 372292 398647
rect 372252 398268 372304 398274
rect 372252 398210 372304 398216
rect 372356 393990 372384 399758
rect 372448 399758 372522 399786
rect 372448 397497 372476 399758
rect 372770 399752 372798 400044
rect 372724 399724 372798 399752
rect 372862 399752 372890 400044
rect 372954 399906 372982 400044
rect 372942 399900 372994 399906
rect 372942 399842 372994 399848
rect 373046 399752 373074 400044
rect 373138 399820 373166 400044
rect 373230 399945 373258 400044
rect 373216 399936 373272 399945
rect 373216 399871 373272 399880
rect 373322 399820 373350 400044
rect 373138 399792 373212 399820
rect 372862 399724 372936 399752
rect 373046 399724 373120 399752
rect 372528 399696 372580 399702
rect 372528 399638 372580 399644
rect 372620 399696 372672 399702
rect 372620 399638 372672 399644
rect 372540 398857 372568 399638
rect 372526 398848 372582 398857
rect 372526 398783 372582 398792
rect 372528 398064 372580 398070
rect 372528 398006 372580 398012
rect 372434 397488 372490 397497
rect 372434 397423 372490 397432
rect 372540 396074 372568 398006
rect 372632 397526 372660 399638
rect 372724 399401 372752 399724
rect 372804 399628 372856 399634
rect 372908 399616 372936 399724
rect 372908 399588 373028 399616
rect 372804 399570 372856 399576
rect 372710 399392 372766 399401
rect 372710 399327 372766 399336
rect 372712 399220 372764 399226
rect 372712 399162 372764 399168
rect 372724 398070 372752 399162
rect 372712 398064 372764 398070
rect 372712 398006 372764 398012
rect 372710 397896 372766 397905
rect 372710 397831 372766 397840
rect 372620 397520 372672 397526
rect 372620 397462 372672 397468
rect 372540 396046 372660 396074
rect 372344 393984 372396 393990
rect 372344 393926 372396 393932
rect 372632 391542 372660 396046
rect 372724 395865 372752 397831
rect 372710 395856 372766 395865
rect 372710 395791 372766 395800
rect 372712 393916 372764 393922
rect 372712 393858 372764 393864
rect 372620 391536 372672 391542
rect 372620 391478 372672 391484
rect 372724 391474 372752 393858
rect 372712 391468 372764 391474
rect 372712 391410 372764 391416
rect 372816 315858 372844 399570
rect 372894 399528 372950 399537
rect 372894 399463 372950 399472
rect 372908 315926 372936 399463
rect 373000 398177 373028 399588
rect 372986 398168 373042 398177
rect 372986 398103 373042 398112
rect 373092 398018 373120 399724
rect 373184 398154 373212 399792
rect 373276 399792 373350 399820
rect 373276 399650 373304 399792
rect 373414 399752 373442 400044
rect 373506 399906 373534 400044
rect 373494 399900 373546 399906
rect 373494 399842 373546 399848
rect 373598 399752 373626 400044
rect 373690 399820 373718 400044
rect 373782 399945 373810 400044
rect 373768 399936 373824 399945
rect 373768 399871 373824 399880
rect 373690 399792 373764 399820
rect 373414 399724 373488 399752
rect 373598 399724 373672 399752
rect 373276 399622 373396 399650
rect 373264 399560 373316 399566
rect 373264 399502 373316 399508
rect 373276 398410 373304 399502
rect 373264 398404 373316 398410
rect 373264 398346 373316 398352
rect 373368 398313 373396 399622
rect 373460 398546 373488 399724
rect 373540 399492 373592 399498
rect 373540 399434 373592 399440
rect 373448 398540 373500 398546
rect 373448 398482 373500 398488
rect 373354 398304 373410 398313
rect 373354 398239 373410 398248
rect 373184 398126 373488 398154
rect 373000 397990 373120 398018
rect 373356 398064 373408 398070
rect 373356 398006 373408 398012
rect 373000 393922 373028 397990
rect 373078 397624 373134 397633
rect 373078 397559 373134 397568
rect 372988 393916 373040 393922
rect 372988 393858 373040 393864
rect 372988 393780 373040 393786
rect 372988 393722 373040 393728
rect 373000 382974 373028 393722
rect 373092 389174 373120 397559
rect 373092 389146 373212 389174
rect 372988 382968 373040 382974
rect 372988 382910 373040 382916
rect 372896 315920 372948 315926
rect 372896 315862 372948 315868
rect 372804 315852 372856 315858
rect 372804 315794 372856 315800
rect 372160 305856 372212 305862
rect 372160 305798 372212 305804
rect 372068 301912 372120 301918
rect 372068 301854 372120 301860
rect 369952 300688 370004 300694
rect 369952 300630 370004 300636
rect 373184 297906 373212 389146
rect 373368 311642 373396 398006
rect 373356 311636 373408 311642
rect 373356 311578 373408 311584
rect 373460 304774 373488 398126
rect 373552 393786 373580 399434
rect 373644 399378 373672 399724
rect 373736 399498 373764 399792
rect 373874 399752 373902 400044
rect 373966 399906 373994 400044
rect 374058 399906 374086 400044
rect 373954 399900 374006 399906
rect 373954 399842 374006 399848
rect 374046 399900 374098 399906
rect 374046 399842 374098 399848
rect 374150 399786 374178 400044
rect 374104 399758 374178 399786
rect 374242 399786 374270 400044
rect 374334 399906 374362 400044
rect 374322 399900 374374 399906
rect 374322 399842 374374 399848
rect 374242 399758 374316 399786
rect 373874 399724 373948 399752
rect 373814 399664 373870 399673
rect 373814 399599 373870 399608
rect 373724 399492 373776 399498
rect 373724 399434 373776 399440
rect 373644 399350 373764 399378
rect 373630 399256 373686 399265
rect 373630 399191 373686 399200
rect 373540 393780 373592 393786
rect 373540 393722 373592 393728
rect 373644 310418 373672 399191
rect 373736 392970 373764 399350
rect 373828 398886 373856 399599
rect 373920 399226 373948 399724
rect 374000 399492 374052 399498
rect 374000 399434 374052 399440
rect 373908 399220 373960 399226
rect 373908 399162 373960 399168
rect 373908 399084 373960 399090
rect 373908 399026 373960 399032
rect 373816 398880 373868 398886
rect 373816 398822 373868 398828
rect 373920 398614 373948 399026
rect 373908 398608 373960 398614
rect 373908 398550 373960 398556
rect 374012 398070 374040 399434
rect 374000 398064 374052 398070
rect 374000 398006 374052 398012
rect 374104 393718 374132 399758
rect 374182 399664 374238 399673
rect 374182 399599 374238 399608
rect 374196 398970 374224 399599
rect 374288 399090 374316 399758
rect 374426 399650 374454 400044
rect 374518 399786 374546 400044
rect 374610 399906 374638 400044
rect 374598 399900 374650 399906
rect 374598 399842 374650 399848
rect 374518 399758 374592 399786
rect 374426 399622 374500 399650
rect 374368 399560 374420 399566
rect 374368 399502 374420 399508
rect 374276 399084 374328 399090
rect 374276 399026 374328 399032
rect 374196 398942 374316 398970
rect 374288 398041 374316 398942
rect 374274 398032 374330 398041
rect 374274 397967 374330 397976
rect 374276 394324 374328 394330
rect 374276 394266 374328 394272
rect 374092 393712 374144 393718
rect 374092 393654 374144 393660
rect 373724 392964 373776 392970
rect 373724 392906 373776 392912
rect 374184 392692 374236 392698
rect 374184 392634 374236 392640
rect 373998 392184 374054 392193
rect 373998 392119 374000 392128
rect 374052 392119 374054 392128
rect 374000 392090 374052 392096
rect 374196 315790 374224 392634
rect 374184 315784 374236 315790
rect 374184 315726 374236 315732
rect 374288 315518 374316 394266
rect 374380 394262 374408 399502
rect 374472 398857 374500 399622
rect 374458 398848 374514 398857
rect 374458 398783 374514 398792
rect 374564 398342 374592 399758
rect 374702 399650 374730 400044
rect 374794 399945 374822 400044
rect 374780 399936 374836 399945
rect 374886 399906 374914 400044
rect 374978 399906 375006 400044
rect 375070 399945 375098 400044
rect 375056 399936 375112 399945
rect 374780 399871 374836 399880
rect 374874 399900 374926 399906
rect 374874 399842 374926 399848
rect 374966 399900 375018 399906
rect 375056 399871 375112 399880
rect 374966 399842 375018 399848
rect 375162 399684 375190 400044
rect 375254 399752 375282 400044
rect 375346 399820 375374 400044
rect 375438 399945 375466 400044
rect 375424 399936 375480 399945
rect 375530 399906 375558 400044
rect 375622 399906 375650 400044
rect 375424 399871 375480 399880
rect 375518 399900 375570 399906
rect 375518 399842 375570 399848
rect 375610 399900 375662 399906
rect 375610 399842 375662 399848
rect 375714 399820 375742 400044
rect 375806 399945 375834 400044
rect 375792 399936 375848 399945
rect 375898 399906 375926 400044
rect 375792 399871 375848 399880
rect 375886 399900 375938 399906
rect 375886 399842 375938 399848
rect 375990 399838 376018 400044
rect 376082 399906 376110 400044
rect 376070 399900 376122 399906
rect 376070 399842 376122 399848
rect 375978 399832 376030 399838
rect 375346 399792 375420 399820
rect 375714 399792 375788 399820
rect 375254 399724 375328 399752
rect 375116 399656 375190 399684
rect 374702 399622 374868 399650
rect 374644 399560 374696 399566
rect 374642 399528 374644 399537
rect 374736 399560 374788 399566
rect 374696 399528 374698 399537
rect 374736 399502 374788 399508
rect 374642 399463 374698 399472
rect 374748 399378 374776 399502
rect 374656 399350 374776 399378
rect 374552 398336 374604 398342
rect 374552 398278 374604 398284
rect 374552 397452 374604 397458
rect 374552 397394 374604 397400
rect 374458 395312 374514 395321
rect 374458 395247 374514 395256
rect 374368 394256 374420 394262
rect 374368 394198 374420 394204
rect 374368 393916 374420 393922
rect 374368 393858 374420 393864
rect 374380 323610 374408 393858
rect 374472 341601 374500 395247
rect 374564 394210 374592 397394
rect 374656 394330 374684 399350
rect 374840 397497 374868 399622
rect 375012 399628 375064 399634
rect 375012 399570 375064 399576
rect 374918 399120 374974 399129
rect 374918 399055 374974 399064
rect 374826 397488 374882 397497
rect 374826 397423 374882 397432
rect 374736 395684 374788 395690
rect 374736 395626 374788 395632
rect 374644 394324 374696 394330
rect 374644 394266 374696 394272
rect 374564 394182 374684 394210
rect 374552 392556 374604 392562
rect 374552 392498 374604 392504
rect 374564 370569 374592 392498
rect 374550 370560 374606 370569
rect 374550 370495 374606 370504
rect 374458 341592 374514 341601
rect 374458 341527 374514 341536
rect 374368 323604 374420 323610
rect 374368 323546 374420 323552
rect 374276 315512 374328 315518
rect 374276 315454 374328 315460
rect 373632 310412 373684 310418
rect 373632 310354 373684 310360
rect 373448 304768 373500 304774
rect 373448 304710 373500 304716
rect 374656 299946 374684 394182
rect 374748 386170 374776 395626
rect 374828 393712 374880 393718
rect 374828 393654 374880 393660
rect 374736 386164 374788 386170
rect 374736 386106 374788 386112
rect 374840 377777 374868 393654
rect 374826 377768 374882 377777
rect 374826 377703 374882 377712
rect 374932 310486 374960 399055
rect 375024 393922 375052 399570
rect 375012 393916 375064 393922
rect 375012 393858 375064 393864
rect 375116 392698 375144 399656
rect 375300 399616 375328 399724
rect 375208 399588 375328 399616
rect 375104 392692 375156 392698
rect 375104 392634 375156 392640
rect 375208 392562 375236 399588
rect 375286 399528 375342 399537
rect 375286 399463 375342 399472
rect 375300 394466 375328 399463
rect 375392 398002 375420 399792
rect 375760 399786 375788 399792
rect 375838 399800 375894 399809
rect 375472 399764 375524 399770
rect 375760 399758 375838 399786
rect 375978 399774 376030 399780
rect 375838 399735 375894 399744
rect 375472 399706 375524 399712
rect 375380 397996 375432 398002
rect 375380 397938 375432 397944
rect 375288 394460 375340 394466
rect 375288 394402 375340 394408
rect 375288 394256 375340 394262
rect 375288 394198 375340 394204
rect 375196 392556 375248 392562
rect 375196 392498 375248 392504
rect 375300 311846 375328 394198
rect 375380 392828 375432 392834
rect 375380 392770 375432 392776
rect 375392 388618 375420 392770
rect 375484 391338 375512 399706
rect 375932 399696 375984 399702
rect 375562 399664 375618 399673
rect 375562 399599 375618 399608
rect 375852 399656 375932 399684
rect 375576 396778 375604 399599
rect 375656 399424 375708 399430
rect 375656 399366 375708 399372
rect 375564 396772 375616 396778
rect 375564 396714 375616 396720
rect 375668 395146 375696 399366
rect 375656 395140 375708 395146
rect 375656 395082 375708 395088
rect 375852 395026 375880 399656
rect 375932 399638 375984 399644
rect 376024 399628 376076 399634
rect 376024 399570 376076 399576
rect 375932 399560 375984 399566
rect 375932 399502 375984 399508
rect 375576 394998 375880 395026
rect 375472 391332 375524 391338
rect 375472 391274 375524 391280
rect 375380 388612 375432 388618
rect 375380 388554 375432 388560
rect 375576 317286 375604 394998
rect 375656 394936 375708 394942
rect 375656 394878 375708 394884
rect 375668 326398 375696 394878
rect 375944 392834 375972 399502
rect 375932 392828 375984 392834
rect 375932 392770 375984 392776
rect 376036 391377 376064 399570
rect 376174 399548 376202 400044
rect 376266 399945 376294 400044
rect 376252 399936 376308 399945
rect 376252 399871 376308 399880
rect 376358 399752 376386 400044
rect 376450 399906 376478 400044
rect 376542 399911 376570 400044
rect 376438 399900 376490 399906
rect 376438 399842 376490 399848
rect 376528 399902 376584 399911
rect 376634 399906 376662 400044
rect 376726 399945 376754 400044
rect 376712 399936 376768 399945
rect 376528 399837 376584 399846
rect 376622 399900 376674 399906
rect 376712 399871 376768 399880
rect 376622 399842 376674 399848
rect 376484 399764 376536 399770
rect 376358 399724 376432 399752
rect 376298 399664 376354 399673
rect 376298 399599 376354 399608
rect 376128 399520 376202 399548
rect 376128 391678 376156 399520
rect 376312 399378 376340 399599
rect 376220 399350 376340 399378
rect 376220 397866 376248 399350
rect 376300 399288 376352 399294
rect 376300 399230 376352 399236
rect 376312 398954 376340 399230
rect 376300 398948 376352 398954
rect 376300 398890 376352 398896
rect 376208 397860 376260 397866
rect 376208 397802 376260 397808
rect 376404 395486 376432 399724
rect 376484 399706 376536 399712
rect 376392 395480 376444 395486
rect 376392 395422 376444 395428
rect 376392 395276 376444 395282
rect 376392 395218 376444 395224
rect 376116 391672 376168 391678
rect 376116 391614 376168 391620
rect 376022 391368 376078 391377
rect 376022 391303 376078 391312
rect 376404 389174 376432 395218
rect 376312 389146 376432 389174
rect 375656 326392 375708 326398
rect 375656 326334 375708 326340
rect 375564 317280 375616 317286
rect 375564 317222 375616 317228
rect 375288 311840 375340 311846
rect 375288 311782 375340 311788
rect 374920 310480 374972 310486
rect 374920 310422 374972 310428
rect 375288 310480 375340 310486
rect 375288 310422 375340 310428
rect 375300 309806 375328 310422
rect 376312 310282 376340 389146
rect 376300 310276 376352 310282
rect 376300 310218 376352 310224
rect 375288 309800 375340 309806
rect 375288 309742 375340 309748
rect 374644 299940 374696 299946
rect 374644 299882 374696 299888
rect 376496 299334 376524 399706
rect 376818 399684 376846 400044
rect 376910 399906 376938 400044
rect 377002 399945 377030 400044
rect 376988 399936 377044 399945
rect 376898 399900 376950 399906
rect 377094 399906 377122 400044
rect 376988 399871 377044 399880
rect 377082 399900 377134 399906
rect 376898 399842 376950 399848
rect 377082 399842 377134 399848
rect 376944 399764 376996 399770
rect 377186 399752 377214 400044
rect 377278 399906 377306 400044
rect 377266 399900 377318 399906
rect 377266 399842 377318 399848
rect 377370 399786 377398 400044
rect 377324 399758 377398 399786
rect 377186 399724 377260 399752
rect 376944 399706 376996 399712
rect 376574 399664 376630 399673
rect 376574 399599 376630 399608
rect 376772 399656 376846 399684
rect 376588 397934 376616 399599
rect 376772 398274 376800 399656
rect 376852 399560 376904 399566
rect 376852 399502 376904 399508
rect 376760 398268 376812 398274
rect 376760 398210 376812 398216
rect 376760 398132 376812 398138
rect 376760 398074 376812 398080
rect 376576 397928 376628 397934
rect 376576 397870 376628 397876
rect 376772 397633 376800 398074
rect 376758 397624 376814 397633
rect 376758 397559 376814 397568
rect 376576 396772 376628 396778
rect 376576 396714 376628 396720
rect 376588 300626 376616 396714
rect 376668 395412 376720 395418
rect 376668 395354 376720 395360
rect 376680 390561 376708 395354
rect 376760 395344 376812 395350
rect 376760 395286 376812 395292
rect 376666 390552 376722 390561
rect 376666 390487 376722 390496
rect 376668 317280 376720 317286
rect 376668 317222 376720 317228
rect 376680 316742 376708 317222
rect 376668 316736 376720 316742
rect 376668 316678 376720 316684
rect 376576 300620 376628 300626
rect 376576 300562 376628 300568
rect 376484 299328 376536 299334
rect 376484 299270 376536 299276
rect 373172 297900 373224 297906
rect 373172 297842 373224 297848
rect 369308 297832 369360 297838
rect 369308 297774 369360 297780
rect 367468 297764 367520 297770
rect 367468 297706 367520 297712
rect 364984 297696 365036 297702
rect 364984 297638 365036 297644
rect 363420 297628 363472 297634
rect 363420 297570 363472 297576
rect 376772 292534 376800 395286
rect 376864 314362 376892 399502
rect 376956 395418 376984 399706
rect 377126 399664 377182 399673
rect 377048 399622 377126 399650
rect 376944 395412 376996 395418
rect 376944 395354 376996 395360
rect 377048 394398 377076 399622
rect 377126 399599 377182 399608
rect 377128 399492 377180 399498
rect 377128 399434 377180 399440
rect 377140 398206 377168 399434
rect 377128 398200 377180 398206
rect 377128 398142 377180 398148
rect 377036 394392 377088 394398
rect 377036 394334 377088 394340
rect 377232 394058 377260 399724
rect 377324 397458 377352 399758
rect 377462 399684 377490 400044
rect 377554 399752 377582 400044
rect 377646 399906 377674 400044
rect 377634 399900 377686 399906
rect 377634 399842 377686 399848
rect 377738 399786 377766 400044
rect 377830 399906 377858 400044
rect 377922 399906 377950 400044
rect 378014 399911 378042 400044
rect 377818 399900 377870 399906
rect 377818 399842 377870 399848
rect 377910 399900 377962 399906
rect 377910 399842 377962 399848
rect 378000 399902 378056 399911
rect 378106 399906 378134 400044
rect 378198 399945 378226 400044
rect 378184 399936 378240 399945
rect 378000 399837 378056 399846
rect 378094 399900 378146 399906
rect 378290 399906 378318 400044
rect 378184 399871 378240 399880
rect 378278 399900 378330 399906
rect 378094 399842 378146 399848
rect 378278 399842 378330 399848
rect 378138 399800 378194 399809
rect 377738 399758 378088 399786
rect 377554 399724 377628 399752
rect 377416 399656 377490 399684
rect 377312 397452 377364 397458
rect 377312 397394 377364 397400
rect 377312 396228 377364 396234
rect 377312 396170 377364 396176
rect 377220 394052 377272 394058
rect 377220 393994 377272 394000
rect 377036 393984 377088 393990
rect 377036 393926 377088 393932
rect 377048 334626 377076 393926
rect 377036 334620 377088 334626
rect 377036 334562 377088 334568
rect 377324 319025 377352 396170
rect 377416 396098 377444 399656
rect 377496 399560 377548 399566
rect 377494 399528 377496 399537
rect 377548 399528 377550 399537
rect 377494 399463 377550 399472
rect 377600 398478 377628 399724
rect 377680 399696 377732 399702
rect 377680 399638 377732 399644
rect 377772 399696 377824 399702
rect 377772 399638 377824 399644
rect 377588 398472 377640 398478
rect 377588 398414 377640 398420
rect 377588 398268 377640 398274
rect 377588 398210 377640 398216
rect 377404 396092 377456 396098
rect 377404 396034 377456 396040
rect 377600 389174 377628 398210
rect 377692 389706 377720 399638
rect 377784 393990 377812 399638
rect 377864 399628 377916 399634
rect 377864 399570 377916 399576
rect 377876 395962 377904 399570
rect 377956 399560 378008 399566
rect 377956 399502 378008 399508
rect 377968 398750 377996 399502
rect 377956 398744 378008 398750
rect 377956 398686 378008 398692
rect 377956 398472 378008 398478
rect 377956 398414 378008 398420
rect 377864 395956 377916 395962
rect 377864 395898 377916 395904
rect 377864 394052 377916 394058
rect 377864 393994 377916 394000
rect 377772 393984 377824 393990
rect 377772 393926 377824 393932
rect 377876 390153 377904 393994
rect 377862 390144 377918 390153
rect 377862 390079 377918 390088
rect 377968 389960 377996 398414
rect 378060 397089 378088 399758
rect 378382 399752 378410 400044
rect 378474 399809 378502 400044
rect 378138 399735 378194 399744
rect 378046 397080 378102 397089
rect 378046 397015 378102 397024
rect 378152 395282 378180 399735
rect 378336 399724 378410 399752
rect 378460 399800 378516 399809
rect 378460 399735 378516 399744
rect 378566 399752 378594 400044
rect 378658 399906 378686 400044
rect 378750 399945 378778 400044
rect 378736 399936 378792 399945
rect 378646 399900 378698 399906
rect 378736 399871 378792 399880
rect 378646 399842 378698 399848
rect 378692 399764 378744 399770
rect 378566 399724 378640 399752
rect 378230 399664 378286 399673
rect 378230 399599 378286 399608
rect 378244 396234 378272 399599
rect 378232 396228 378284 396234
rect 378232 396170 378284 396176
rect 378336 395418 378364 399724
rect 378416 399628 378468 399634
rect 378416 399570 378468 399576
rect 378324 395412 378376 395418
rect 378324 395354 378376 395360
rect 378322 395312 378378 395321
rect 378140 395276 378192 395282
rect 378322 395247 378378 395256
rect 378140 395218 378192 395224
rect 378140 395140 378192 395146
rect 378140 395082 378192 395088
rect 378152 390114 378180 395082
rect 378140 390108 378192 390114
rect 378140 390050 378192 390056
rect 377968 389932 378180 389960
rect 378152 389774 378180 389932
rect 377956 389768 378008 389774
rect 377956 389710 378008 389716
rect 378140 389768 378192 389774
rect 378140 389710 378192 389716
rect 377680 389700 377732 389706
rect 377680 389642 377732 389648
rect 377600 389146 377720 389174
rect 377310 319016 377366 319025
rect 377310 318951 377366 318960
rect 376852 314356 376904 314362
rect 376852 314298 376904 314304
rect 377692 313070 377720 389146
rect 377968 386102 377996 389710
rect 378048 389700 378100 389706
rect 378048 389642 378100 389648
rect 377956 386096 378008 386102
rect 377956 386038 378008 386044
rect 378060 316810 378088 389642
rect 378048 316804 378100 316810
rect 378048 316746 378100 316752
rect 378336 314294 378364 395247
rect 378428 323678 378456 399570
rect 378508 399492 378560 399498
rect 378508 399434 378560 399440
rect 378520 395350 378548 399434
rect 378612 399265 378640 399724
rect 378692 399706 378744 399712
rect 378598 399256 378654 399265
rect 378598 399191 378654 399200
rect 378704 395690 378732 399706
rect 378842 399684 378870 400044
rect 378934 399906 378962 400044
rect 379026 399906 379054 400044
rect 379118 399906 379146 400044
rect 378922 399900 378974 399906
rect 378922 399842 378974 399848
rect 379014 399900 379066 399906
rect 379014 399842 379066 399848
rect 379106 399900 379158 399906
rect 379106 399842 379158 399848
rect 379210 399786 379238 400044
rect 379164 399758 379238 399786
rect 378796 399656 378870 399684
rect 379060 399696 379112 399702
rect 378692 395684 378744 395690
rect 378692 395626 378744 395632
rect 378692 395480 378744 395486
rect 378692 395422 378744 395428
rect 378508 395344 378560 395350
rect 378508 395286 378560 395292
rect 378704 389174 378732 395422
rect 378796 395146 378824 399656
rect 379060 399638 379112 399644
rect 379072 397610 379100 399638
rect 378980 397582 379100 397610
rect 378784 395140 378836 395146
rect 378784 395082 378836 395088
rect 378980 390046 379008 397582
rect 379164 397497 379192 399758
rect 379302 399650 379330 400044
rect 379394 399906 379422 400044
rect 379486 399945 379514 400044
rect 379472 399936 379528 399945
rect 379382 399900 379434 399906
rect 379472 399871 379528 399880
rect 379382 399842 379434 399848
rect 379578 399838 379606 400044
rect 379566 399832 379618 399838
rect 379566 399774 379618 399780
rect 379428 399764 379480 399770
rect 379428 399706 379480 399712
rect 379256 399622 379330 399650
rect 379150 397488 379206 397497
rect 379150 397423 379206 397432
rect 379060 395480 379112 395486
rect 379060 395422 379112 395428
rect 378968 390040 379020 390046
rect 378968 389982 379020 389988
rect 378612 389146 378732 389174
rect 378416 323672 378468 323678
rect 378416 323614 378468 323620
rect 378324 314288 378376 314294
rect 378324 314230 378376 314236
rect 378336 313954 378364 314230
rect 378324 313948 378376 313954
rect 378324 313890 378376 313896
rect 377680 313064 377732 313070
rect 377680 313006 377732 313012
rect 378612 299470 378640 389146
rect 379072 318918 379100 395422
rect 379150 395312 379206 395321
rect 379150 395247 379206 395256
rect 379060 318912 379112 318918
rect 379060 318854 379112 318860
rect 379164 311545 379192 395247
rect 379256 314090 379284 399622
rect 379336 399560 379388 399566
rect 379336 399502 379388 399508
rect 379348 392834 379376 399502
rect 379440 399208 379468 399706
rect 379670 399684 379698 400044
rect 379762 399945 379790 400044
rect 379748 399936 379804 399945
rect 379854 399906 379882 400044
rect 379946 399945 379974 400044
rect 379932 399936 379988 399945
rect 379748 399871 379804 399880
rect 379842 399900 379894 399906
rect 379932 399871 379988 399880
rect 379842 399842 379894 399848
rect 379796 399764 379848 399770
rect 380038 399752 380066 400044
rect 379796 399706 379848 399712
rect 379992 399724 380066 399752
rect 379624 399656 379698 399684
rect 379440 399180 379560 399208
rect 379532 398041 379560 399180
rect 379624 399158 379652 399656
rect 379612 399152 379664 399158
rect 379612 399094 379664 399100
rect 379612 398948 379664 398954
rect 379808 398936 379836 399706
rect 379888 399492 379940 399498
rect 379888 399434 379940 399440
rect 379612 398890 379664 398896
rect 379716 398908 379836 398936
rect 379518 398032 379574 398041
rect 379518 397967 379574 397976
rect 379428 395344 379480 395350
rect 379428 395286 379480 395292
rect 379336 392828 379388 392834
rect 379336 392770 379388 392776
rect 379440 389978 379468 395286
rect 379428 389972 379480 389978
rect 379428 389914 379480 389920
rect 379624 315761 379652 398890
rect 379716 331294 379744 398908
rect 379900 398886 379928 399434
rect 379888 398880 379940 398886
rect 379888 398822 379940 398828
rect 379992 398818 380020 399724
rect 380130 399684 380158 400044
rect 380222 399707 380250 400044
rect 380314 399906 380342 400044
rect 380406 399911 380434 400044
rect 380302 399900 380354 399906
rect 380302 399842 380354 399848
rect 380392 399902 380448 399911
rect 380498 399906 380526 400044
rect 380590 399945 380618 400044
rect 380576 399936 380632 399945
rect 380392 399837 380448 399846
rect 380486 399900 380538 399906
rect 380576 399871 380632 399880
rect 380486 399842 380538 399848
rect 380682 399786 380710 400044
rect 380774 399906 380802 400044
rect 380866 399945 380894 400044
rect 380852 399936 380908 399945
rect 380762 399900 380814 399906
rect 380958 399906 380986 400044
rect 381050 399945 381078 400044
rect 381036 399936 381092 399945
rect 380852 399871 380908 399880
rect 380946 399900 380998 399906
rect 380762 399842 380814 399848
rect 381036 399871 381092 399880
rect 380946 399842 380998 399848
rect 381142 399809 381170 400044
rect 380806 399800 380862 399809
rect 380682 399758 380756 399786
rect 380084 399656 380158 399684
rect 380208 399698 380264 399707
rect 379796 398812 379848 398818
rect 379796 398754 379848 398760
rect 379980 398812 380032 398818
rect 379980 398754 380032 398760
rect 379808 395486 379836 398754
rect 379980 398676 380032 398682
rect 379980 398618 380032 398624
rect 379796 395480 379848 395486
rect 379796 395422 379848 395428
rect 379796 395344 379848 395350
rect 379796 395286 379848 395292
rect 379808 383382 379836 395286
rect 379888 391876 379940 391882
rect 379888 391818 379940 391824
rect 379900 387258 379928 391818
rect 379888 387252 379940 387258
rect 379888 387194 379940 387200
rect 379796 383376 379848 383382
rect 379796 383318 379848 383324
rect 379704 331288 379756 331294
rect 379704 331230 379756 331236
rect 379716 330585 379744 331230
rect 379702 330576 379758 330585
rect 379702 330511 379758 330520
rect 379610 315752 379666 315761
rect 379610 315687 379666 315696
rect 379992 315178 380020 398618
rect 380084 395298 380112 399656
rect 380532 399696 380584 399702
rect 380208 399633 380264 399642
rect 380346 399664 380402 399673
rect 380346 399599 380402 399608
rect 380452 399656 380532 399684
rect 380256 399560 380308 399566
rect 380256 399502 380308 399508
rect 380164 399288 380216 399294
rect 380164 399230 380216 399236
rect 380176 398818 380204 399230
rect 380268 399226 380296 399502
rect 380256 399220 380308 399226
rect 380256 399162 380308 399168
rect 380164 398812 380216 398818
rect 380164 398754 380216 398760
rect 380256 395412 380308 395418
rect 380256 395354 380308 395360
rect 380084 395270 380204 395298
rect 380072 392828 380124 392834
rect 380072 392770 380124 392776
rect 379980 315172 380032 315178
rect 379980 315114 380032 315120
rect 380084 314430 380112 392770
rect 380176 386753 380204 395270
rect 380268 387326 380296 395354
rect 380360 395350 380388 399599
rect 380348 395344 380400 395350
rect 380348 395286 380400 395292
rect 380256 387320 380308 387326
rect 380256 387262 380308 387268
rect 380162 386744 380218 386753
rect 380162 386679 380218 386688
rect 380072 314424 380124 314430
rect 380072 314366 380124 314372
rect 379244 314084 379296 314090
rect 379244 314026 379296 314032
rect 379150 311536 379206 311545
rect 379150 311471 379206 311480
rect 380452 307737 380480 399656
rect 380532 399638 380584 399644
rect 380622 399664 380678 399673
rect 380622 399599 380678 399608
rect 380532 399152 380584 399158
rect 380532 399094 380584 399100
rect 380544 390425 380572 399094
rect 380636 399022 380664 399599
rect 380624 399016 380676 399022
rect 380624 398958 380676 398964
rect 380728 391882 380756 399758
rect 381128 399800 381184 399809
rect 380862 399758 380940 399786
rect 380806 399735 380862 399744
rect 380808 399696 380860 399702
rect 380808 399638 380860 399644
rect 380820 398954 380848 399638
rect 380808 398948 380860 398954
rect 380808 398890 380860 398896
rect 380912 398546 380940 399758
rect 381234 399786 381262 400044
rect 381326 399906 381354 400044
rect 381418 399906 381446 400044
rect 381510 399906 381538 400044
rect 381314 399900 381366 399906
rect 381314 399842 381366 399848
rect 381406 399900 381458 399906
rect 381406 399842 381458 399848
rect 381498 399900 381550 399906
rect 381498 399842 381550 399848
rect 381602 399786 381630 400044
rect 381694 399906 381722 400044
rect 381682 399900 381734 399906
rect 381682 399842 381734 399848
rect 381786 399786 381814 400044
rect 381234 399758 381400 399786
rect 381602 399758 381676 399786
rect 381128 399735 381184 399744
rect 381266 399664 381322 399673
rect 381084 399628 381136 399634
rect 381266 399599 381268 399608
rect 381084 399570 381136 399576
rect 381320 399599 381322 399608
rect 381268 399570 381320 399576
rect 380900 398540 380952 398546
rect 380900 398482 380952 398488
rect 380806 398440 380862 398449
rect 380862 398398 381032 398426
rect 380806 398375 380862 398384
rect 380898 393544 380954 393553
rect 380898 393479 380954 393488
rect 380912 393446 380940 393479
rect 380900 393440 380952 393446
rect 380900 393382 380952 393388
rect 380716 391876 380768 391882
rect 380716 391818 380768 391824
rect 380530 390416 380586 390425
rect 380530 390351 380586 390360
rect 381004 389842 381032 398398
rect 381096 394194 381124 399570
rect 381176 399560 381228 399566
rect 381228 399508 381308 399514
rect 381176 399502 381308 399508
rect 381188 399486 381308 399502
rect 381176 399424 381228 399430
rect 381176 399366 381228 399372
rect 381084 394188 381136 394194
rect 381084 394130 381136 394136
rect 381084 393984 381136 393990
rect 381084 393926 381136 393932
rect 380992 389836 381044 389842
rect 380992 389778 381044 389784
rect 380900 327140 380952 327146
rect 380900 327082 380952 327088
rect 380912 326369 380940 327082
rect 380898 326360 380954 326369
rect 380898 326295 380954 326304
rect 380900 323060 380952 323066
rect 380900 323002 380952 323008
rect 380912 322250 380940 323002
rect 380900 322244 380952 322250
rect 380900 322186 380952 322192
rect 381096 308961 381124 393926
rect 381188 313041 381216 399366
rect 381280 394694 381308 399486
rect 381372 398834 381400 399758
rect 381452 399696 381504 399702
rect 381452 399638 381504 399644
rect 381544 399696 381596 399702
rect 381544 399638 381596 399644
rect 381464 399430 381492 399638
rect 381452 399424 381504 399430
rect 381452 399366 381504 399372
rect 381372 398806 381492 398834
rect 381464 398546 381492 398806
rect 381452 398540 381504 398546
rect 381452 398482 381504 398488
rect 381452 397928 381504 397934
rect 381452 397870 381504 397876
rect 381280 394666 381400 394694
rect 381268 392896 381320 392902
rect 381268 392838 381320 392844
rect 381280 323066 381308 392838
rect 381372 327146 381400 394666
rect 381360 327140 381412 327146
rect 381360 327082 381412 327088
rect 381268 323060 381320 323066
rect 381268 323002 381320 323008
rect 381174 313032 381230 313041
rect 381174 312967 381230 312976
rect 381464 311817 381492 397870
rect 381556 396982 381584 399638
rect 381648 399430 381676 399758
rect 381740 399758 381814 399786
rect 381878 399786 381906 400044
rect 381970 399906 381998 400044
rect 381958 399900 382010 399906
rect 381958 399842 382010 399848
rect 381878 399758 381952 399786
rect 381636 399424 381688 399430
rect 381636 399366 381688 399372
rect 381634 399256 381690 399265
rect 381634 399191 381690 399200
rect 381544 396976 381596 396982
rect 381544 396918 381596 396924
rect 381544 394732 381596 394738
rect 381544 394674 381596 394680
rect 381556 385937 381584 394674
rect 381648 389174 381676 399191
rect 381740 392902 381768 399758
rect 381820 399696 381872 399702
rect 381820 399638 381872 399644
rect 381728 392896 381780 392902
rect 381728 392838 381780 392844
rect 381648 389146 381768 389174
rect 381542 385928 381598 385937
rect 381542 385863 381598 385872
rect 381544 322992 381596 322998
rect 381544 322934 381596 322940
rect 381450 311808 381506 311817
rect 381450 311743 381506 311752
rect 381082 308952 381138 308961
rect 381082 308887 381138 308896
rect 380438 307728 380494 307737
rect 380438 307663 380494 307672
rect 381556 301510 381584 322934
rect 381740 307562 381768 389146
rect 381728 307556 381780 307562
rect 381728 307498 381780 307504
rect 381832 304842 381860 399638
rect 381924 399090 381952 399758
rect 382062 399752 382090 400044
rect 382154 399906 382182 400044
rect 382142 399900 382194 399906
rect 382142 399842 382194 399848
rect 382246 399820 382274 400044
rect 382338 399945 382366 400044
rect 382324 399936 382380 399945
rect 382430 399906 382458 400044
rect 382324 399871 382380 399880
rect 382418 399900 382470 399906
rect 382418 399842 382470 399848
rect 382246 399792 382320 399820
rect 382016 399724 382090 399752
rect 381912 399084 381964 399090
rect 381912 399026 381964 399032
rect 382016 393990 382044 399724
rect 382188 399696 382240 399702
rect 382188 399638 382240 399644
rect 382096 399424 382148 399430
rect 382096 399366 382148 399372
rect 382108 399158 382136 399366
rect 382096 399152 382148 399158
rect 382096 399094 382148 399100
rect 382094 398168 382150 398177
rect 382094 398103 382150 398112
rect 382108 397633 382136 398103
rect 382094 397624 382150 397633
rect 382094 397559 382150 397568
rect 382200 397497 382228 399638
rect 382292 399430 382320 399792
rect 382522 399786 382550 400044
rect 382384 399758 382550 399786
rect 382280 399424 382332 399430
rect 382280 399366 382332 399372
rect 382384 398478 382412 399758
rect 382614 399650 382642 400044
rect 382706 399752 382734 400044
rect 382798 399945 382826 400044
rect 382784 399936 382840 399945
rect 382784 399871 382840 399880
rect 382890 399820 382918 400044
rect 382982 399911 383010 400044
rect 382968 399902 383024 399911
rect 383074 399906 383102 400044
rect 383166 399945 383194 400044
rect 383152 399936 383208 399945
rect 382968 399837 383024 399846
rect 383062 399900 383114 399906
rect 383258 399906 383286 400044
rect 383152 399871 383208 399880
rect 383246 399900 383298 399906
rect 383062 399842 383114 399848
rect 383246 399842 383298 399848
rect 382844 399792 382918 399820
rect 383198 399800 383254 399809
rect 382706 399724 382780 399752
rect 382614 399622 382688 399650
rect 382556 399560 382608 399566
rect 382476 399520 382556 399548
rect 382372 398472 382424 398478
rect 382372 398414 382424 398420
rect 382186 397488 382242 397497
rect 382186 397423 382242 397432
rect 382280 397316 382332 397322
rect 382280 397258 382332 397264
rect 382004 393984 382056 393990
rect 382004 393926 382056 393932
rect 382292 387190 382320 397258
rect 382280 387184 382332 387190
rect 382280 387126 382332 387132
rect 382476 342961 382504 399520
rect 382556 399502 382608 399508
rect 382556 399424 382608 399430
rect 382556 399366 382608 399372
rect 382568 398070 382596 399366
rect 382660 398750 382688 399622
rect 382648 398744 382700 398750
rect 382648 398686 382700 398692
rect 382556 398064 382608 398070
rect 382556 398006 382608 398012
rect 382646 398032 382702 398041
rect 382646 397967 382702 397976
rect 382556 394052 382608 394058
rect 382556 393994 382608 394000
rect 382568 383314 382596 393994
rect 382556 383308 382608 383314
rect 382556 383250 382608 383256
rect 382462 342952 382518 342961
rect 382462 342887 382518 342896
rect 381820 304836 381872 304842
rect 381820 304778 381872 304784
rect 381544 301504 381596 301510
rect 381544 301446 381596 301452
rect 378600 299464 378652 299470
rect 378600 299406 378652 299412
rect 376760 292528 376812 292534
rect 376760 292470 376812 292476
rect 378140 292528 378192 292534
rect 378140 292470 378192 292476
rect 374092 260976 374144 260982
rect 374092 260918 374144 260924
rect 371240 255400 371292 255406
rect 371240 255342 371292 255348
rect 363604 140140 363656 140146
rect 363604 140082 363656 140088
rect 361578 62792 361634 62801
rect 361578 62727 361634 62736
rect 361592 16574 361620 62727
rect 360212 16546 361160 16574
rect 361592 16546 361896 16574
rect 359924 4072 359976 4078
rect 359924 4014 359976 4020
rect 359464 3392 359516 3398
rect 359464 3334 359516 3340
rect 359936 480 359964 4014
rect 361132 480 361160 16546
rect 345726 354 345838 480
rect 345308 326 345838 354
rect 345726 -960 345838 326
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 361868 354 361896 16546
rect 363616 4146 363644 140082
rect 369860 134632 369912 134638
rect 369860 134574 369912 134580
rect 365810 102912 365866 102921
rect 365810 102847 365866 102856
rect 363604 4140 363656 4146
rect 363604 4082 363656 4088
rect 364616 3732 364668 3738
rect 364616 3674 364668 3680
rect 363512 3392 363564 3398
rect 363512 3334 363564 3340
rect 363524 480 363552 3334
rect 364628 480 364656 3674
rect 365824 480 365852 102847
rect 368478 61432 368534 61441
rect 368478 61367 368534 61376
rect 368492 16574 368520 61367
rect 369872 16574 369900 134574
rect 368492 16546 369440 16574
rect 369872 16546 370176 16574
rect 367008 4140 367060 4146
rect 367008 4082 367060 4088
rect 367020 480 367048 4082
rect 368204 3868 368256 3874
rect 368204 3810 368256 3816
rect 368216 480 368244 3810
rect 369412 480 369440 16546
rect 362286 354 362398 480
rect 361868 326 362398 354
rect 362286 -960 362398 326
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370148 354 370176 16546
rect 370566 354 370678 480
rect 370148 326 370678 354
rect 371252 354 371280 255342
rect 372618 58576 372674 58585
rect 372618 58511 372674 58520
rect 372632 16574 372660 58511
rect 372632 16546 372936 16574
rect 372908 480 372936 16546
rect 374000 3664 374052 3670
rect 374000 3606 374052 3612
rect 374012 1850 374040 3606
rect 374104 3398 374132 260918
rect 376024 142860 376076 142866
rect 376024 142802 376076 142808
rect 376036 16574 376064 142802
rect 376760 133272 376812 133278
rect 376760 133214 376812 133220
rect 376772 16574 376800 133214
rect 378152 16574 378180 292470
rect 376036 16546 376156 16574
rect 376772 16546 377720 16574
rect 378152 16546 378456 16574
rect 376024 10328 376076 10334
rect 376024 10270 376076 10276
rect 374092 3392 374144 3398
rect 374092 3334 374144 3340
rect 375288 3392 375340 3398
rect 375288 3334 375340 3340
rect 374012 1822 374132 1850
rect 374104 480 374132 1822
rect 375300 480 375328 3334
rect 371670 354 371782 480
rect 371252 326 371782 354
rect 370566 -960 370678 326
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 354 376064 10270
rect 376128 3398 376156 16546
rect 376116 3392 376168 3398
rect 376116 3334 376168 3340
rect 377692 480 377720 16546
rect 376454 354 376566 480
rect 376036 326 376566 354
rect 376454 -960 376566 326
rect 377650 -960 377762 480
rect 378428 354 378456 16546
rect 379978 6488 380034 6497
rect 379978 6423 380034 6432
rect 379992 480 380020 6423
rect 381556 3738 381584 301446
rect 382660 297974 382688 397967
rect 382752 393854 382780 399724
rect 382844 398682 382872 399792
rect 383108 399764 383160 399770
rect 383350 399786 383378 400044
rect 383198 399735 383254 399744
rect 383304 399758 383378 399786
rect 383108 399706 383160 399712
rect 382832 398676 382884 398682
rect 382832 398618 382884 398624
rect 383016 398676 383068 398682
rect 383016 398618 383068 398624
rect 382832 398404 382884 398410
rect 382832 398346 382884 398352
rect 382740 393848 382792 393854
rect 382740 393790 382792 393796
rect 382844 315314 382872 398346
rect 383028 393938 383056 398618
rect 383120 394126 383148 399706
rect 383212 397322 383240 399735
rect 383304 398313 383332 399758
rect 383442 399650 383470 400044
rect 383396 399622 383470 399650
rect 383290 398304 383346 398313
rect 383290 398239 383346 398248
rect 383292 397928 383344 397934
rect 383292 397870 383344 397876
rect 383200 397316 383252 397322
rect 383200 397258 383252 397264
rect 383304 395350 383332 397870
rect 383292 395344 383344 395350
rect 383292 395286 383344 395292
rect 383108 394120 383160 394126
rect 383108 394062 383160 394068
rect 383396 394058 383424 399622
rect 383534 399514 383562 400044
rect 383626 399752 383654 400044
rect 383718 399906 383746 400044
rect 383810 399945 383838 400044
rect 383796 399936 383852 399945
rect 383706 399900 383758 399906
rect 383902 399906 383930 400044
rect 383796 399871 383852 399880
rect 383890 399900 383942 399906
rect 383706 399842 383758 399848
rect 383890 399842 383942 399848
rect 383750 399800 383806 399809
rect 383626 399724 383700 399752
rect 383994 399786 384022 400044
rect 384086 399911 384114 400044
rect 384072 399902 384128 399911
rect 384072 399837 384128 399846
rect 383750 399735 383806 399744
rect 383856 399758 384022 399786
rect 384178 399786 384206 400044
rect 384270 399906 384298 400044
rect 384258 399900 384310 399906
rect 384258 399842 384310 399848
rect 384362 399786 384390 400044
rect 384454 399911 384482 400044
rect 384440 399902 384496 399911
rect 384440 399837 384496 399846
rect 384546 399786 384574 400044
rect 384638 399906 384666 400044
rect 384626 399900 384678 399906
rect 384626 399842 384678 399848
rect 384730 399786 384758 400044
rect 384822 399906 384850 400044
rect 384810 399900 384862 399906
rect 384810 399842 384862 399848
rect 384914 399786 384942 400044
rect 385006 399911 385034 400044
rect 384992 399902 385048 399911
rect 384992 399837 385048 399846
rect 385098 399786 385126 400044
rect 384178 399758 384252 399786
rect 383488 399486 383562 399514
rect 383488 397633 383516 399486
rect 383568 399424 383620 399430
rect 383568 399366 383620 399372
rect 383580 397934 383608 399366
rect 383672 398410 383700 399724
rect 383660 398404 383712 398410
rect 383660 398346 383712 398352
rect 383660 398268 383712 398274
rect 383660 398210 383712 398216
rect 383568 397928 383620 397934
rect 383568 397870 383620 397876
rect 383568 397792 383620 397798
rect 383568 397734 383620 397740
rect 383474 397624 383530 397633
rect 383474 397559 383530 397568
rect 383384 394052 383436 394058
rect 383384 393994 383436 394000
rect 383028 393910 383424 393938
rect 383292 393848 383344 393854
rect 383292 393790 383344 393796
rect 382832 315308 382884 315314
rect 382832 315250 382884 315256
rect 383304 302734 383332 393790
rect 383396 322998 383424 393910
rect 383580 389174 383608 397734
rect 383672 397526 383700 398210
rect 383660 397520 383712 397526
rect 383660 397462 383712 397468
rect 383764 394074 383792 399735
rect 383856 394194 383884 399758
rect 383936 399696 383988 399702
rect 383936 399638 383988 399644
rect 384120 399696 384172 399702
rect 384120 399638 384172 399644
rect 383948 397934 383976 399638
rect 384132 399242 384160 399638
rect 384040 399214 384160 399242
rect 384040 398041 384068 399214
rect 384118 399120 384174 399129
rect 384118 399055 384174 399064
rect 384026 398032 384082 398041
rect 384026 397967 384082 397976
rect 383936 397928 383988 397934
rect 383936 397870 383988 397876
rect 383844 394188 383896 394194
rect 383844 394130 383896 394136
rect 383764 394046 383976 394074
rect 383844 393916 383896 393922
rect 383844 393858 383896 393864
rect 383752 393848 383804 393854
rect 383752 393790 383804 393796
rect 383488 389146 383608 389174
rect 383384 322992 383436 322998
rect 383384 322934 383436 322940
rect 383488 315450 383516 389146
rect 383764 340105 383792 393790
rect 383856 349110 383884 393858
rect 383948 356697 383976 394046
rect 384132 389174 384160 399055
rect 384224 397798 384252 399758
rect 384316 399758 384390 399786
rect 384500 399758 384574 399786
rect 384684 399758 384758 399786
rect 384868 399758 384942 399786
rect 385052 399758 385126 399786
rect 384212 397792 384264 397798
rect 384212 397734 384264 397740
rect 384212 395956 384264 395962
rect 384212 395898 384264 395904
rect 384224 393582 384252 395898
rect 384316 394738 384344 399758
rect 384500 399378 384528 399758
rect 384580 399696 384632 399702
rect 384580 399638 384632 399644
rect 384408 399350 384528 399378
rect 384408 397746 384436 399350
rect 384488 399220 384540 399226
rect 384488 399162 384540 399168
rect 384500 397866 384528 399162
rect 384592 398449 384620 399638
rect 384578 398440 384634 398449
rect 384578 398375 384634 398384
rect 384684 398177 384712 399758
rect 384868 399378 384896 399758
rect 384948 399696 385000 399702
rect 384948 399638 385000 399644
rect 384776 399350 384896 399378
rect 384670 398168 384726 398177
rect 384670 398103 384726 398112
rect 384488 397860 384540 397866
rect 384488 397802 384540 397808
rect 384408 397730 384712 397746
rect 384408 397724 384724 397730
rect 384408 397718 384672 397724
rect 384672 397666 384724 397672
rect 384396 397520 384448 397526
rect 384396 397462 384448 397468
rect 384304 394732 384356 394738
rect 384304 394674 384356 394680
rect 384212 393576 384264 393582
rect 384212 393518 384264 393524
rect 384040 389146 384160 389174
rect 384408 389174 384436 397462
rect 384672 396092 384724 396098
rect 384672 396034 384724 396040
rect 384684 393666 384712 396034
rect 384776 393854 384804 399350
rect 384854 399256 384910 399265
rect 384960 399226 384988 399638
rect 384854 399191 384910 399200
rect 384948 399220 385000 399226
rect 384764 393848 384816 393854
rect 384764 393790 384816 393796
rect 384684 393638 384804 393666
rect 384672 393576 384724 393582
rect 384672 393518 384724 393524
rect 384408 389146 384620 389174
rect 384040 366382 384068 389146
rect 384028 366376 384080 366382
rect 384028 366318 384080 366324
rect 383934 356688 383990 356697
rect 383934 356623 383990 356632
rect 383844 349104 383896 349110
rect 383844 349046 383896 349052
rect 384396 349104 384448 349110
rect 384396 349046 384448 349052
rect 384408 347818 384436 349046
rect 384396 347812 384448 347818
rect 384396 347754 384448 347760
rect 383750 340096 383806 340105
rect 383750 340031 383806 340040
rect 383476 315444 383528 315450
rect 383476 315386 383528 315392
rect 384408 313177 384436 347754
rect 384592 315382 384620 389146
rect 384580 315376 384632 315382
rect 384580 315318 384632 315324
rect 384684 314498 384712 393518
rect 384672 314492 384724 314498
rect 384672 314434 384724 314440
rect 384394 313168 384450 313177
rect 384394 313103 384450 313112
rect 383292 302728 383344 302734
rect 383292 302670 383344 302676
rect 384776 300801 384804 393638
rect 384868 388822 384896 399191
rect 384948 399162 385000 399168
rect 384946 398984 385002 398993
rect 384946 398919 385002 398928
rect 384856 388816 384908 388822
rect 384856 388758 384908 388764
rect 384960 323649 384988 398919
rect 385052 393854 385080 399758
rect 385190 399650 385218 400044
rect 385282 399786 385310 400044
rect 385374 399945 385402 400044
rect 385360 399936 385416 399945
rect 385466 399906 385494 400044
rect 385360 399871 385416 399880
rect 385454 399900 385506 399906
rect 385454 399842 385506 399848
rect 385282 399758 385356 399786
rect 385144 399622 385218 399650
rect 385144 393990 385172 399622
rect 385222 399528 385278 399537
rect 385222 399463 385278 399472
rect 385132 393984 385184 393990
rect 385132 393926 385184 393932
rect 385040 393848 385092 393854
rect 385040 393790 385092 393796
rect 385236 334014 385264 399463
rect 385328 395622 385356 399758
rect 385558 399650 385586 400044
rect 385650 399752 385678 400044
rect 385742 399906 385770 400044
rect 385834 399945 385862 400044
rect 385820 399936 385876 399945
rect 385730 399900 385782 399906
rect 385926 399906 385954 400044
rect 386018 399906 386046 400044
rect 385820 399871 385876 399880
rect 385914 399900 385966 399906
rect 385730 399842 385782 399848
rect 385914 399842 385966 399848
rect 386006 399900 386058 399906
rect 386006 399842 386058 399848
rect 386110 399786 386138 400044
rect 386202 399906 386230 400044
rect 386294 399945 386322 400044
rect 386280 399936 386336 399945
rect 386190 399900 386242 399906
rect 386386 399906 386414 400044
rect 386280 399871 386336 399880
rect 386374 399900 386426 399906
rect 386190 399842 386242 399848
rect 386374 399842 386426 399848
rect 386478 399838 386506 400044
rect 386466 399832 386518 399838
rect 386110 399758 386184 399786
rect 386466 399774 386518 399780
rect 386570 399786 386598 400044
rect 386662 399945 386690 400044
rect 386648 399936 386704 399945
rect 386648 399871 386704 399880
rect 386754 399786 386782 400044
rect 386846 399945 386874 400044
rect 386832 399936 386888 399945
rect 386938 399906 386966 400044
rect 387030 399906 387058 400044
rect 387122 399945 387150 400044
rect 387108 399936 387164 399945
rect 386832 399871 386888 399880
rect 386926 399900 386978 399906
rect 386926 399842 386978 399848
rect 387018 399900 387070 399906
rect 387108 399871 387164 399880
rect 387018 399842 387070 399848
rect 387214 399820 387242 400044
rect 387306 399922 387334 400044
rect 387412 400030 387472 400058
rect 387306 399894 387380 399922
rect 385650 399724 385724 399752
rect 385420 399622 385586 399650
rect 385420 396846 385448 399622
rect 385696 399566 385724 399724
rect 385868 399696 385920 399702
rect 385868 399638 385920 399644
rect 386052 399696 386104 399702
rect 386156 399673 386184 399758
rect 386328 399764 386380 399770
rect 386570 399758 386644 399786
rect 386328 399706 386380 399712
rect 386052 399638 386104 399644
rect 386142 399664 386198 399673
rect 385592 399560 385644 399566
rect 385498 399528 385554 399537
rect 385592 399502 385644 399508
rect 385684 399560 385736 399566
rect 385684 399502 385736 399508
rect 385498 399463 385554 399472
rect 385408 396840 385460 396846
rect 385408 396782 385460 396788
rect 385316 395616 385368 395622
rect 385316 395558 385368 395564
rect 385316 393984 385368 393990
rect 385316 393926 385368 393932
rect 385328 341465 385356 393926
rect 385512 389174 385540 399463
rect 385604 396137 385632 399502
rect 385684 399424 385736 399430
rect 385684 399366 385736 399372
rect 385590 396128 385646 396137
rect 385590 396063 385646 396072
rect 385696 393938 385724 399366
rect 385880 399242 385908 399638
rect 385776 399220 385828 399226
rect 385880 399214 386000 399242
rect 385776 399162 385828 399168
rect 385788 398818 385816 399162
rect 385868 399152 385920 399158
rect 385868 399094 385920 399100
rect 385880 399022 385908 399094
rect 385868 399016 385920 399022
rect 385868 398958 385920 398964
rect 385866 398848 385922 398857
rect 385776 398812 385828 398818
rect 385866 398783 385922 398792
rect 385776 398754 385828 398760
rect 385880 397526 385908 398783
rect 385868 397520 385920 397526
rect 385868 397462 385920 397468
rect 385696 393910 385908 393938
rect 385776 393848 385828 393854
rect 385776 393790 385828 393796
rect 385420 389146 385540 389174
rect 385420 359514 385448 389146
rect 385408 359508 385460 359514
rect 385408 359450 385460 359456
rect 385314 341456 385370 341465
rect 385314 341391 385370 341400
rect 385224 334008 385276 334014
rect 385224 333950 385276 333956
rect 385684 334008 385736 334014
rect 385684 333950 385736 333956
rect 384946 323640 385002 323649
rect 384946 323575 385002 323584
rect 385696 317257 385724 333950
rect 385788 324358 385816 393790
rect 385776 324352 385828 324358
rect 385776 324294 385828 324300
rect 385788 323785 385816 324294
rect 385774 323776 385830 323785
rect 385774 323711 385830 323720
rect 385880 322153 385908 393910
rect 385972 386034 386000 399214
rect 386064 397905 386092 399638
rect 386142 399599 386198 399608
rect 386050 397896 386106 397905
rect 386050 397831 386106 397840
rect 386052 397452 386104 397458
rect 386052 397394 386104 397400
rect 385960 386028 386012 386034
rect 385960 385970 386012 385976
rect 385866 322144 385922 322153
rect 385866 322079 385922 322088
rect 385682 317248 385738 317257
rect 385682 317183 385738 317192
rect 386064 313818 386092 397394
rect 386340 394942 386368 399706
rect 386510 399664 386566 399673
rect 386420 399628 386472 399634
rect 386510 399599 386566 399608
rect 386420 399570 386472 399576
rect 386328 394936 386380 394942
rect 386328 394878 386380 394884
rect 386432 392970 386460 399570
rect 386420 392964 386472 392970
rect 386420 392906 386472 392912
rect 386524 317121 386552 399599
rect 386616 393990 386644 399758
rect 386708 399758 386782 399786
rect 387168 399792 387242 399820
rect 386708 397662 386736 399758
rect 386788 399696 386840 399702
rect 386788 399638 386840 399644
rect 386972 399696 387024 399702
rect 386972 399638 387024 399644
rect 386696 397656 386748 397662
rect 386696 397598 386748 397604
rect 386800 397594 386828 399638
rect 386878 399528 386934 399537
rect 386878 399463 386934 399472
rect 386788 397588 386840 397594
rect 386788 397530 386840 397536
rect 386696 397384 386748 397390
rect 386892 397338 386920 399463
rect 386696 397326 386748 397332
rect 386604 393984 386656 393990
rect 386604 393926 386656 393932
rect 386604 390788 386656 390794
rect 386604 390730 386656 390736
rect 386616 321609 386644 390730
rect 386708 327729 386736 397326
rect 386800 397310 386920 397338
rect 386800 330449 386828 397310
rect 386984 394694 387012 399638
rect 386892 394666 387012 394694
rect 386892 390794 386920 394666
rect 386880 390788 386932 390794
rect 386880 390730 386932 390736
rect 386880 390652 386932 390658
rect 386880 390594 386932 390600
rect 386892 333305 386920 390594
rect 387168 389174 387196 399792
rect 387352 397390 387380 399894
rect 387340 397384 387392 397390
rect 387340 397326 387392 397332
rect 387340 393984 387392 393990
rect 387340 393926 387392 393932
rect 386984 389146 387196 389174
rect 386984 338774 387012 389146
rect 386972 338768 387024 338774
rect 386972 338710 387024 338716
rect 386878 333296 386934 333305
rect 386878 333231 386934 333240
rect 386786 330440 386842 330449
rect 386786 330375 386842 330384
rect 386694 327720 386750 327729
rect 386694 327655 386750 327664
rect 386602 321600 386658 321609
rect 386602 321535 386658 321544
rect 387062 321600 387118 321609
rect 387062 321535 387118 321544
rect 386510 317112 386566 317121
rect 386510 317047 386566 317056
rect 386052 313812 386104 313818
rect 386052 313754 386104 313760
rect 384762 300792 384818 300801
rect 384762 300727 384818 300736
rect 382648 297968 382700 297974
rect 382648 297910 382700 297916
rect 385040 253224 385092 253230
rect 385040 253166 385092 253172
rect 382280 251320 382332 251326
rect 382280 251262 382332 251268
rect 381636 151088 381688 151094
rect 381636 151030 381688 151036
rect 381648 3942 381676 151030
rect 382292 16574 382320 251262
rect 384302 155272 384358 155281
rect 384302 155207 384358 155216
rect 382292 16546 382412 16574
rect 381636 3936 381688 3942
rect 381636 3878 381688 3884
rect 381544 3732 381596 3738
rect 381544 3674 381596 3680
rect 381176 3392 381228 3398
rect 381176 3334 381228 3340
rect 381188 480 381216 3334
rect 382384 480 382412 16546
rect 383568 6316 383620 6322
rect 383568 6258 383620 6264
rect 383580 480 383608 6258
rect 384316 3874 384344 155207
rect 385052 16574 385080 253166
rect 385052 16546 386000 16574
rect 384764 3936 384816 3942
rect 384764 3878 384816 3884
rect 384304 3868 384356 3874
rect 384304 3810 384356 3816
rect 384776 480 384804 3878
rect 385972 480 386000 16546
rect 387076 3670 387104 321535
rect 387352 314265 387380 393926
rect 387444 390658 387472 400030
rect 387536 398954 387564 400318
rect 389546 400208 389602 400217
rect 389546 400143 389602 400152
rect 387984 399492 388036 399498
rect 387984 399434 388036 399440
rect 387524 398948 387576 398954
rect 387524 398890 387576 398896
rect 387800 398200 387852 398206
rect 387800 398142 387852 398148
rect 387432 390652 387484 390658
rect 387432 390594 387484 390600
rect 387338 314256 387394 314265
rect 387338 314191 387394 314200
rect 387812 304230 387840 398142
rect 387892 397792 387944 397798
rect 387892 397734 387944 397740
rect 387904 310185 387932 397734
rect 387996 311137 388024 399434
rect 389272 398744 389324 398750
rect 389272 398686 389324 398692
rect 389180 398608 389232 398614
rect 389180 398550 389232 398556
rect 388168 398404 388220 398410
rect 388168 398346 388220 398352
rect 388076 398064 388128 398070
rect 388076 398006 388128 398012
rect 388088 312322 388116 398006
rect 388180 314401 388208 398346
rect 388258 398304 388314 398313
rect 388258 398239 388314 398248
rect 388272 318102 388300 398239
rect 388260 318096 388312 318102
rect 388260 318038 388312 318044
rect 388166 314392 388222 314401
rect 388166 314327 388222 314336
rect 388076 312316 388128 312322
rect 388076 312258 388128 312264
rect 387982 311128 388038 311137
rect 387982 311063 388038 311072
rect 387890 310176 387946 310185
rect 387890 310111 387946 310120
rect 389192 306377 389220 398550
rect 389178 306368 389234 306377
rect 389178 306303 389234 306312
rect 389284 306241 389312 398686
rect 389364 398200 389416 398206
rect 389364 398142 389416 398148
rect 389376 308242 389404 398142
rect 389456 397928 389508 397934
rect 389456 397870 389508 397876
rect 389468 312594 389496 397870
rect 389560 313750 389588 400143
rect 390650 400072 390706 400081
rect 390650 400007 390706 400016
rect 392032 400036 392084 400042
rect 390560 399968 390612 399974
rect 390560 399910 390612 399916
rect 389640 398472 389692 398478
rect 389640 398414 389692 398420
rect 389652 317218 389680 398414
rect 389640 317212 389692 317218
rect 389640 317154 389692 317160
rect 389548 313744 389600 313750
rect 389548 313686 389600 313692
rect 389456 312588 389508 312594
rect 389456 312530 389508 312536
rect 390572 310049 390600 399910
rect 390664 312662 390692 400007
rect 392032 399978 392084 399984
rect 390928 397860 390980 397866
rect 390928 397802 390980 397808
rect 390744 397520 390796 397526
rect 390744 397462 390796 397468
rect 390756 314537 390784 397462
rect 390834 396944 390890 396953
rect 390834 396879 390890 396888
rect 390848 315217 390876 396879
rect 390940 317393 390968 397802
rect 391940 397588 391992 397594
rect 391940 397530 391992 397536
rect 390926 317384 390982 317393
rect 390926 317319 390982 317328
rect 390834 315208 390890 315217
rect 390834 315143 390890 315152
rect 390742 314528 390798 314537
rect 390742 314463 390798 314472
rect 390652 312656 390704 312662
rect 390652 312598 390704 312604
rect 390558 310040 390614 310049
rect 390558 309975 390614 309984
rect 389364 308236 389416 308242
rect 389364 308178 389416 308184
rect 389270 306232 389326 306241
rect 389270 306167 389326 306176
rect 391952 306105 391980 397530
rect 392044 309097 392072 399978
rect 580264 399492 580316 399498
rect 580264 399434 580316 399440
rect 393320 399084 393372 399090
rect 393320 399026 393372 399032
rect 392216 398540 392268 398546
rect 392216 398482 392268 398488
rect 392122 398032 392178 398041
rect 392122 397967 392178 397976
rect 392136 310321 392164 397967
rect 392228 312390 392256 398482
rect 392308 397724 392360 397730
rect 392308 397666 392360 397672
rect 392320 316470 392348 397666
rect 393136 397656 393188 397662
rect 393136 397598 393188 397604
rect 393148 394806 393176 397598
rect 393136 394800 393188 394806
rect 393136 394742 393188 394748
rect 392308 316464 392360 316470
rect 392308 316406 392360 316412
rect 392216 312384 392268 312390
rect 392216 312326 392268 312332
rect 393332 310457 393360 399026
rect 393504 399016 393556 399022
rect 393504 398958 393556 398964
rect 393412 398880 393464 398886
rect 393412 398822 393464 398828
rect 393424 313993 393452 398822
rect 393516 316674 393544 398958
rect 394976 398948 395028 398954
rect 394976 398890 395028 398896
rect 394792 395344 394844 395350
rect 394792 395286 394844 395292
rect 394700 394800 394752 394806
rect 394700 394742 394752 394748
rect 393504 316668 393556 316674
rect 393504 316610 393556 316616
rect 393410 313984 393466 313993
rect 393410 313919 393466 313928
rect 393318 310448 393374 310457
rect 393318 310383 393374 310392
rect 392122 310312 392178 310321
rect 392122 310247 392178 310256
rect 392030 309088 392086 309097
rect 392030 309023 392086 309032
rect 391938 306096 391994 306105
rect 391938 306031 391994 306040
rect 387800 304224 387852 304230
rect 387800 304166 387852 304172
rect 394712 290494 394740 394742
rect 394804 302190 394832 395286
rect 394884 394936 394936 394942
rect 394884 394878 394936 394884
rect 394896 303521 394924 394878
rect 394988 307766 395016 398890
rect 577502 387016 577558 387025
rect 577502 386951 577558 386960
rect 534724 369980 534776 369986
rect 534724 369922 534776 369928
rect 534080 347812 534132 347818
rect 534080 347754 534132 347760
rect 427818 338192 427874 338201
rect 427818 338127 427874 338136
rect 398932 315308 398984 315314
rect 398932 315250 398984 315256
rect 394976 307760 395028 307766
rect 394976 307702 395028 307708
rect 395988 307760 396040 307766
rect 395988 307702 396040 307708
rect 396000 307086 396028 307702
rect 395988 307080 396040 307086
rect 395988 307022 396040 307028
rect 394882 303512 394938 303521
rect 394882 303447 394938 303456
rect 395986 303512 396042 303521
rect 395986 303447 396042 303456
rect 396000 302938 396028 303447
rect 395988 302932 396040 302938
rect 395988 302874 396040 302880
rect 394792 302184 394844 302190
rect 394792 302126 394844 302132
rect 394700 290488 394752 290494
rect 394700 290430 394752 290436
rect 396080 259480 396132 259486
rect 396080 259422 396132 259428
rect 389180 256828 389232 256834
rect 389180 256770 389232 256776
rect 387800 131844 387852 131850
rect 387800 131786 387852 131792
rect 387156 6248 387208 6254
rect 387156 6190 387208 6196
rect 387064 3664 387116 3670
rect 387064 3606 387116 3612
rect 387168 480 387196 6190
rect 378846 354 378958 480
rect 378428 326 378958 354
rect 378846 -960 378958 326
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 387812 354 387840 131786
rect 389192 16574 389220 256770
rect 391940 253972 391992 253978
rect 391940 253914 391992 253920
rect 390560 126336 390612 126342
rect 390560 126278 390612 126284
rect 389192 16546 389496 16574
rect 389468 480 389496 16546
rect 390572 3398 390600 126278
rect 391952 16574 391980 253914
rect 394700 123548 394752 123554
rect 394700 123490 394752 123496
rect 394712 16574 394740 123490
rect 391952 16546 392624 16574
rect 394712 16546 395384 16574
rect 390650 6352 390706 6361
rect 390650 6287 390706 6296
rect 390560 3392 390612 3398
rect 390560 3334 390612 3340
rect 390664 480 390692 6287
rect 391848 3392 391900 3398
rect 391848 3334 391900 3340
rect 391860 480 391888 3334
rect 388230 354 388342 480
rect 387812 326 388342 354
rect 388230 -960 388342 326
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 354 392624 16546
rect 394238 6216 394294 6225
rect 394238 6151 394294 6160
rect 394252 480 394280 6151
rect 395356 480 395384 16546
rect 393014 354 393126 480
rect 392596 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 259422
rect 397458 21312 397514 21321
rect 397458 21247 397514 21256
rect 397472 16574 397500 21247
rect 397472 16546 397776 16574
rect 397748 480 397776 16546
rect 398840 3868 398892 3874
rect 398840 3810 398892 3816
rect 398852 1986 398880 3810
rect 398944 3398 398972 315250
rect 414020 309800 414072 309806
rect 414020 309742 414072 309748
rect 409880 307080 409932 307086
rect 409880 307022 409932 307028
rect 407120 248600 407172 248606
rect 407120 248542 407172 248548
rect 405740 147008 405792 147014
rect 405740 146950 405792 146956
rect 399484 138780 399536 138786
rect 399484 138722 399536 138728
rect 398932 3392 398984 3398
rect 398932 3334 398984 3340
rect 399496 3058 399524 138722
rect 404360 116612 404412 116618
rect 404360 116554 404412 116560
rect 400218 82104 400274 82113
rect 400218 82039 400274 82048
rect 400232 16574 400260 82039
rect 400232 16546 400904 16574
rect 400128 3392 400180 3398
rect 400128 3334 400180 3340
rect 399484 3052 399536 3058
rect 399484 2994 399536 3000
rect 398852 1958 398972 1986
rect 398944 480 398972 1958
rect 400140 480 400168 3334
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 400876 354 400904 16546
rect 403624 3800 403676 3806
rect 403624 3742 403676 3748
rect 402520 3052 402572 3058
rect 402520 2994 402572 3000
rect 402532 480 402560 2994
rect 403636 480 403664 3742
rect 401294 354 401406 480
rect 400876 326 401406 354
rect 401294 -960 401406 326
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404372 354 404400 116554
rect 405752 16574 405780 146950
rect 405752 16546 406056 16574
rect 406028 480 406056 16546
rect 407132 3210 407160 248542
rect 408500 130416 408552 130422
rect 408500 130358 408552 130364
rect 407210 54496 407266 54505
rect 407210 54431 407266 54440
rect 407224 3398 407252 54431
rect 408512 16574 408540 130358
rect 409892 16574 409920 307022
rect 412640 122120 412692 122126
rect 412640 122062 412692 122068
rect 411258 53136 411314 53145
rect 411258 53071 411314 53080
rect 411272 16574 411300 53071
rect 408512 16546 409184 16574
rect 409892 16546 410840 16574
rect 411272 16546 411944 16574
rect 407212 3392 407264 3398
rect 407212 3334 407264 3340
rect 408408 3392 408460 3398
rect 408408 3334 408460 3340
rect 407132 3182 407252 3210
rect 407224 480 407252 3182
rect 408420 480 408448 3334
rect 404790 354 404902 480
rect 404372 326 404902 354
rect 404790 -960 404902 326
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 354 409184 16546
rect 410812 480 410840 16546
rect 411916 480 411944 16546
rect 409574 354 409686 480
rect 409156 326 409686 354
rect 409574 -960 409686 326
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 354 412680 122062
rect 414032 16574 414060 309742
rect 416780 272536 416832 272542
rect 416780 272478 416832 272484
rect 415400 141500 415452 141506
rect 415400 141442 415452 141448
rect 414032 16546 414336 16574
rect 414308 480 414336 16546
rect 415412 2106 415440 141442
rect 416792 16574 416820 272478
rect 423772 247104 423824 247110
rect 423772 247046 423824 247052
rect 420920 243092 420972 243098
rect 420920 243034 420972 243040
rect 419540 137284 419592 137290
rect 419540 137226 419592 137232
rect 419552 16574 419580 137226
rect 416792 16546 417464 16574
rect 419552 16546 420224 16574
rect 415490 9344 415546 9353
rect 415490 9279 415546 9288
rect 415400 2100 415452 2106
rect 415400 2042 415452 2048
rect 415504 480 415532 9279
rect 416688 2100 416740 2106
rect 416688 2042 416740 2048
rect 416700 480 416728 2042
rect 413070 354 413182 480
rect 412652 326 413182 354
rect 413070 -960 413182 326
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 16546
rect 418986 9208 419042 9217
rect 418986 9143 419042 9152
rect 419000 480 419028 9143
rect 420196 480 420224 16546
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 417854 -960 417966 326
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 420932 354 420960 243034
rect 422944 129124 422996 129130
rect 422944 129066 422996 129072
rect 422576 9104 422628 9110
rect 422576 9046 422628 9052
rect 422588 480 422616 9046
rect 422956 3058 422984 129066
rect 423784 3398 423812 247046
rect 425060 183592 425112 183598
rect 425060 183534 425112 183540
rect 425072 16574 425100 183534
rect 426438 120864 426494 120873
rect 426438 120799 426494 120808
rect 426452 16574 426480 120799
rect 427832 16574 427860 338127
rect 513378 335472 513434 335481
rect 513378 335407 513434 335416
rect 481640 331288 481692 331294
rect 481640 331230 481692 331236
rect 429844 316736 429896 316742
rect 429844 316678 429896 316684
rect 425072 16546 425744 16574
rect 426452 16546 426848 16574
rect 427832 16546 428504 16574
rect 423772 3392 423824 3398
rect 423772 3334 423824 3340
rect 424968 3392 425020 3398
rect 424968 3334 425020 3340
rect 422944 3052 422996 3058
rect 422944 2994 422996 3000
rect 423772 3052 423824 3058
rect 423772 2994 423824 3000
rect 423784 480 423812 2994
rect 424980 480 425008 3334
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 425716 354 425744 16546
rect 426134 354 426246 480
rect 425716 326 426246 354
rect 426820 354 426848 16546
rect 428476 480 428504 16546
rect 429198 14512 429254 14521
rect 429198 14447 429254 14456
rect 427238 354 427350 480
rect 426820 326 427350 354
rect 426134 -960 426246 326
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429212 354 429240 14447
rect 429856 4146 429884 316678
rect 477498 313984 477554 313993
rect 466460 313948 466512 313954
rect 477498 313919 477554 313928
rect 466460 313890 466512 313896
rect 463700 260908 463752 260914
rect 463700 260850 463752 260856
rect 459560 257372 459612 257378
rect 459560 257314 459612 257320
rect 456800 256760 456852 256766
rect 456800 256702 456852 256708
rect 445760 255332 445812 255338
rect 445760 255274 445812 255280
rect 434720 251864 434772 251870
rect 434720 251806 434772 251812
rect 430580 156664 430632 156670
rect 430580 156606 430632 156612
rect 430592 16574 430620 156606
rect 433340 17264 433392 17270
rect 433340 17206 433392 17212
rect 433352 16574 433380 17206
rect 434732 16574 434760 251806
rect 441620 248532 441672 248538
rect 441620 248474 441672 248480
rect 438860 245676 438912 245682
rect 438860 245618 438912 245624
rect 436744 144288 436796 144294
rect 436744 144230 436796 144236
rect 430592 16546 430896 16574
rect 433352 16546 434024 16574
rect 434732 16546 435128 16574
rect 429844 4140 429896 4146
rect 429844 4082 429896 4088
rect 430868 480 430896 16546
rect 433248 9036 433300 9042
rect 433248 8978 433300 8984
rect 432052 4140 432104 4146
rect 432052 4082 432104 4088
rect 432064 480 432092 4082
rect 433260 480 433288 8978
rect 429630 354 429742 480
rect 429212 326 429742 354
rect 429630 -960 429742 326
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 433996 354 434024 16546
rect 434414 354 434526 480
rect 433996 326 434526 354
rect 435100 354 435128 16546
rect 436756 3058 436784 144230
rect 438872 16574 438900 245618
rect 440240 135992 440292 135998
rect 440240 135934 440292 135940
rect 438872 16546 439176 16574
rect 436834 9072 436890 9081
rect 436834 9007 436890 9016
rect 436744 3052 436796 3058
rect 436744 2994 436796 3000
rect 436848 2938 436876 9007
rect 437940 3052 437992 3058
rect 437940 2994 437992 3000
rect 436756 2910 436876 2938
rect 436756 480 436784 2910
rect 437952 480 437980 2994
rect 439148 480 439176 16546
rect 440252 2106 440280 135934
rect 441632 16574 441660 248474
rect 444380 127696 444432 127702
rect 444380 127638 444432 127644
rect 444392 16574 444420 127638
rect 441632 16546 442672 16574
rect 444392 16546 445064 16574
rect 440330 8936 440386 8945
rect 440330 8871 440386 8880
rect 440240 2100 440292 2106
rect 440240 2042 440292 2048
rect 440344 480 440372 8871
rect 441528 2100 441580 2106
rect 441528 2042 441580 2048
rect 441540 480 441568 2042
rect 442644 480 442672 16546
rect 443828 8968 443880 8974
rect 443828 8910 443880 8916
rect 443840 480 443868 8910
rect 445036 480 445064 16546
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 434414 -960 434526 326
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 445772 354 445800 255274
rect 452660 247716 452712 247722
rect 452660 247658 452712 247664
rect 448520 244520 448572 244526
rect 448520 244462 448572 244468
rect 447140 186380 447192 186386
rect 447140 186322 447192 186328
rect 447152 16574 447180 186322
rect 447152 16546 447456 16574
rect 447428 480 447456 16546
rect 448532 2514 448560 244462
rect 449900 187740 449952 187746
rect 449900 187682 449952 187688
rect 448610 118008 448666 118017
rect 448610 117943 448666 117952
rect 448520 2508 448572 2514
rect 448520 2450 448572 2456
rect 448624 480 448652 117943
rect 449912 16574 449940 187682
rect 451280 149728 451332 149734
rect 451280 149670 451332 149676
rect 451292 16574 451320 149670
rect 452672 16574 452700 247658
rect 455420 133204 455472 133210
rect 455420 133146 455472 133152
rect 454040 73840 454092 73846
rect 454040 73782 454092 73788
rect 449912 16546 450952 16574
rect 451292 16546 451688 16574
rect 452672 16546 453344 16574
rect 449808 2508 449860 2514
rect 449808 2450 449860 2456
rect 449820 480 449848 2450
rect 450924 480 450952 16546
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 451660 354 451688 16546
rect 453316 480 453344 16546
rect 452078 354 452190 480
rect 451660 326 452190 354
rect 452078 -960 452190 326
rect 453274 -960 453386 480
rect 454052 354 454080 73782
rect 455432 16574 455460 133146
rect 456812 16574 456840 256702
rect 458180 126268 458232 126274
rect 458180 126210 458232 126216
rect 458192 16574 458220 126210
rect 459572 16574 459600 257314
rect 462318 116512 462374 116521
rect 462318 116447 462374 116456
rect 460938 76528 460994 76537
rect 460938 76463 460994 76472
rect 460952 16574 460980 76463
rect 455432 16546 455736 16574
rect 456812 16546 456932 16574
rect 458192 16546 459232 16574
rect 459572 16546 459968 16574
rect 460952 16546 461624 16574
rect 455708 480 455736 16546
rect 456904 480 456932 16546
rect 458086 3632 458142 3641
rect 458086 3567 458142 3576
rect 458100 480 458128 3567
rect 459204 480 459232 16546
rect 454470 354 454582 480
rect 454052 326 454582 354
rect 454470 -960 454582 326
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 16546
rect 461596 480 461624 16546
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462332 354 462360 116447
rect 463712 16574 463740 260850
rect 465080 140072 465132 140078
rect 465080 140014 465132 140020
rect 465092 16574 465120 140014
rect 466472 16574 466500 313890
rect 471244 252680 471296 252686
rect 471244 252622 471296 252628
rect 470600 249824 470652 249830
rect 470600 249766 470652 249772
rect 468484 131776 468536 131782
rect 468484 131718 468536 131724
rect 463712 16546 464016 16574
rect 465092 16546 465856 16574
rect 466472 16546 467512 16574
rect 463988 480 464016 16546
rect 465170 3496 465226 3505
rect 465170 3431 465226 3440
rect 465184 480 465212 3431
rect 462750 354 462862 480
rect 462332 326 462862 354
rect 462750 -960 462862 326
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 465828 354 465856 16546
rect 467484 480 467512 16546
rect 468496 3534 468524 131718
rect 468300 3528 468352 3534
rect 468300 3470 468352 3476
rect 468484 3528 468536 3534
rect 468484 3470 468536 3476
rect 469864 3528 469916 3534
rect 469864 3470 469916 3476
rect 466246 354 466358 480
rect 465828 326 466358 354
rect 466246 -960 466358 326
rect 467442 -960 467554 480
rect 468312 354 468340 3470
rect 469876 480 469904 3470
rect 468638 354 468750 480
rect 468312 326 468750 354
rect 468638 -960 468750 326
rect 469834 -960 469946 480
rect 470612 354 470640 249766
rect 471256 3126 471284 252622
rect 476120 124908 476172 124914
rect 476120 124850 476172 124856
rect 472622 115152 472678 115161
rect 472622 115087 472678 115096
rect 472636 3534 472664 115087
rect 476132 16574 476160 124850
rect 477512 16574 477540 313919
rect 478880 173936 478932 173942
rect 478880 173878 478932 173884
rect 476132 16546 476528 16574
rect 477512 16546 478184 16574
rect 475752 6180 475804 6186
rect 475752 6122 475804 6128
rect 472624 3528 472676 3534
rect 472624 3470 472676 3476
rect 473452 3528 473504 3534
rect 473452 3470 473504 3476
rect 472256 3460 472308 3466
rect 472256 3402 472308 3408
rect 471244 3120 471296 3126
rect 471244 3062 471296 3068
rect 472268 480 472296 3402
rect 473464 480 473492 3470
rect 474556 3120 474608 3126
rect 474556 3062 474608 3068
rect 474568 480 474596 3062
rect 475764 480 475792 6122
rect 471030 354 471142 480
rect 470612 326 471142 354
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476500 354 476528 16546
rect 478156 480 478184 16546
rect 476918 354 477030 480
rect 476500 326 477030 354
rect 476918 -960 477030 326
rect 478114 -960 478226 480
rect 478892 354 478920 173878
rect 480260 129056 480312 129062
rect 480260 128998 480312 129004
rect 480272 16574 480300 128998
rect 481652 16574 481680 331230
rect 495440 327140 495492 327146
rect 495440 327082 495492 327088
rect 491300 252612 491352 252618
rect 491300 252554 491352 252560
rect 484400 248464 484452 248470
rect 484400 248406 484452 248412
rect 483020 153264 483072 153270
rect 483020 153206 483072 153212
rect 483032 16574 483060 153206
rect 484412 16574 484440 248406
rect 488540 238808 488592 238814
rect 488540 238750 488592 238756
rect 485778 111072 485834 111081
rect 485778 111007 485834 111016
rect 485792 16574 485820 111007
rect 487158 39264 487214 39273
rect 487158 39199 487214 39208
rect 480272 16546 480576 16574
rect 481652 16546 481772 16574
rect 483032 16546 484072 16574
rect 484412 16546 484808 16574
rect 485792 16546 486464 16574
rect 480548 480 480576 16546
rect 481744 480 481772 16546
rect 482834 3360 482890 3369
rect 482834 3295 482890 3304
rect 482848 480 482876 3295
rect 484044 480 484072 16546
rect 479310 354 479422 480
rect 478892 326 479422 354
rect 479310 -960 479422 326
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 484780 354 484808 16546
rect 486436 480 486464 16546
rect 485198 354 485310 480
rect 484780 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487172 354 487200 39199
rect 488552 16574 488580 238750
rect 490012 127628 490064 127634
rect 490012 127570 490064 127576
rect 489184 109744 489236 109750
rect 489184 109686 489236 109692
rect 488552 16546 488856 16574
rect 488828 480 488856 16546
rect 489196 4146 489224 109686
rect 490024 16574 490052 127570
rect 491312 16574 491340 252554
rect 494060 154624 494112 154630
rect 494060 154566 494112 154572
rect 492680 108316 492732 108322
rect 492680 108258 492732 108264
rect 492692 16574 492720 108258
rect 494072 16574 494100 154566
rect 490024 16546 490696 16574
rect 491312 16546 492352 16574
rect 492692 16546 493088 16574
rect 494072 16546 494744 16574
rect 489184 4140 489236 4146
rect 489184 4082 489236 4088
rect 489920 4140 489972 4146
rect 489920 4082 489972 4088
rect 489932 480 489960 4082
rect 487590 354 487702 480
rect 487172 326 487702 354
rect 487590 -960 487702 326
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490668 354 490696 16546
rect 492324 480 492352 16546
rect 491086 354 491198 480
rect 490668 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493060 354 493088 16546
rect 494716 480 494744 16546
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495452 354 495480 327082
rect 506480 322992 506532 322998
rect 506480 322934 506532 322940
rect 498200 312588 498252 312594
rect 498200 312530 498252 312536
rect 496818 106856 496874 106865
rect 496818 106791 496874 106800
rect 496832 16574 496860 106791
rect 496832 16546 497136 16574
rect 497108 480 497136 16546
rect 498212 3534 498240 312530
rect 502338 312488 502394 312497
rect 502338 312423 502394 312432
rect 498290 151192 498346 151201
rect 498290 151127 498346 151136
rect 498200 3528 498252 3534
rect 498200 3470 498252 3476
rect 498304 3346 498332 151127
rect 500960 148368 501012 148374
rect 500960 148310 501012 148316
rect 499580 35216 499632 35222
rect 499580 35158 499632 35164
rect 499592 16574 499620 35158
rect 500972 16574 501000 148310
rect 502352 16574 502380 312423
rect 503720 123480 503772 123486
rect 503720 123422 503772 123428
rect 499592 16546 500632 16574
rect 500972 16546 501368 16574
rect 502352 16546 503024 16574
rect 499028 3528 499080 3534
rect 499028 3470 499080 3476
rect 498212 3318 498332 3346
rect 498212 480 498240 3318
rect 495870 354 495982 480
rect 495452 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499040 354 499068 3470
rect 500604 480 500632 16546
rect 499366 354 499478 480
rect 499040 326 499478 354
rect 499366 -960 499478 326
rect 500562 -960 500674 480
rect 501340 354 501368 16546
rect 502996 480 503024 16546
rect 501758 354 501870 480
rect 501340 326 501870 354
rect 501758 -960 501870 326
rect 502954 -960 503066 480
rect 503732 354 503760 123422
rect 505376 15904 505428 15910
rect 505376 15846 505428 15852
rect 505388 480 505416 15846
rect 506492 480 506520 322934
rect 507860 153332 507912 153338
rect 507860 153274 507912 153280
rect 506570 105496 506626 105505
rect 506570 105431 506626 105440
rect 506584 16574 506612 105431
rect 507872 16574 507900 153274
rect 512000 152584 512052 152590
rect 512000 152526 512052 152532
rect 510618 104136 510674 104145
rect 510618 104071 510674 104080
rect 510632 16574 510660 104071
rect 506584 16546 507256 16574
rect 507872 16546 508912 16574
rect 510632 16546 511304 16574
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507228 354 507256 16546
rect 508884 480 508912 16546
rect 510068 3596 510120 3602
rect 510068 3538 510120 3544
rect 510080 480 510108 3538
rect 511276 480 511304 16546
rect 507646 354 507758 480
rect 507228 326 507758 354
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512012 354 512040 152526
rect 512430 354 512542 480
rect 512012 326 512542 354
rect 513392 354 513420 335407
rect 531320 273964 531372 273970
rect 531320 273906 531372 273912
rect 523132 267776 523184 267782
rect 523132 267718 523184 267724
rect 516140 244452 516192 244458
rect 516140 244394 516192 244400
rect 514024 145580 514076 145586
rect 514024 145522 514076 145528
rect 514036 3058 514064 145522
rect 514850 102776 514906 102785
rect 514850 102711 514906 102720
rect 514864 6914 514892 102711
rect 516152 16574 516180 244394
rect 518900 155984 518952 155990
rect 518900 155926 518952 155932
rect 517520 101448 517572 101454
rect 517520 101390 517572 101396
rect 517532 16574 517560 101390
rect 518912 16574 518940 155926
rect 522304 155236 522356 155242
rect 522304 155178 522356 155184
rect 520922 122088 520978 122097
rect 520922 122023 520978 122032
rect 516152 16546 517192 16574
rect 517532 16546 517928 16574
rect 518912 16546 519584 16574
rect 514772 6886 514892 6914
rect 514024 3052 514076 3058
rect 514024 2994 514076 3000
rect 514772 480 514800 6886
rect 515956 3052 516008 3058
rect 515956 2994 516008 3000
rect 515968 480 515996 2994
rect 517164 480 517192 16546
rect 513534 354 513646 480
rect 513392 326 513646 354
rect 512430 -960 512542 326
rect 513534 -960 513646 326
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 517900 354 517928 16546
rect 519556 480 519584 16546
rect 520740 3800 520792 3806
rect 520740 3742 520792 3748
rect 520752 480 520780 3742
rect 520936 3534 520964 122023
rect 522316 3534 522344 155178
rect 523144 16574 523172 267718
rect 527180 239420 527232 239426
rect 527180 239362 527232 239368
rect 525800 37936 525852 37942
rect 525800 37878 525852 37884
rect 524420 33788 524472 33794
rect 524420 33730 524472 33736
rect 524432 16574 524460 33730
rect 525812 16574 525840 37878
rect 527192 16574 527220 239362
rect 529938 149696 529994 149705
rect 529938 149631 529994 149640
rect 528558 98696 528614 98705
rect 528558 98631 528614 98640
rect 523144 16546 523816 16574
rect 524432 16546 525472 16574
rect 525812 16546 526208 16574
rect 527192 16546 527864 16574
rect 520924 3528 520976 3534
rect 520924 3470 520976 3476
rect 521844 3528 521896 3534
rect 521844 3470 521896 3476
rect 522304 3528 522356 3534
rect 522304 3470 522356 3476
rect 523040 3528 523092 3534
rect 523040 3470 523092 3476
rect 521856 480 521884 3470
rect 523052 480 523080 3470
rect 518318 354 518430 480
rect 517900 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 523788 354 523816 16546
rect 525444 480 525472 16546
rect 524206 354 524318 480
rect 523788 326 524318 354
rect 524206 -960 524318 326
rect 525402 -960 525514 480
rect 526180 354 526208 16546
rect 527836 480 527864 16546
rect 526598 354 526710 480
rect 526180 326 526710 354
rect 526598 -960 526710 326
rect 527794 -960 527906 480
rect 528572 354 528600 98631
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 529952 354 529980 149631
rect 531332 480 531360 273906
rect 532700 144220 532752 144226
rect 532700 144162 532752 144168
rect 531410 97200 531466 97209
rect 531410 97135 531466 97144
rect 531424 16574 531452 97135
rect 532712 16574 532740 144162
rect 534092 16574 534120 347754
rect 534736 313274 534764 369922
rect 552020 334008 552072 334014
rect 552020 333950 552072 333956
rect 547972 324352 548024 324358
rect 547972 324294 548024 324300
rect 534724 313268 534776 313274
rect 534724 313210 534776 313216
rect 538220 251252 538272 251258
rect 538220 251194 538272 251200
rect 536838 151056 536894 151065
rect 536838 150991 536894 151000
rect 535460 94512 535512 94518
rect 535460 94454 535512 94460
rect 535472 16574 535500 94454
rect 536852 16574 536880 150991
rect 531424 16546 532096 16574
rect 532712 16546 533752 16574
rect 534092 16546 534488 16574
rect 535472 16546 536144 16574
rect 536852 16546 537248 16574
rect 530094 354 530206 480
rect 529952 326 530206 354
rect 528990 -960 529102 326
rect 530094 -960 530206 326
rect 531290 -960 531402 480
rect 532068 354 532096 16546
rect 533724 480 533752 16546
rect 532486 354 532598 480
rect 532068 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534460 354 534488 16546
rect 536116 480 536144 16546
rect 537220 480 537248 16546
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538232 354 538260 251194
rect 540980 244384 541032 244390
rect 540980 244326 541032 244332
rect 539598 120728 539654 120737
rect 539598 120663 539654 120672
rect 539612 480 539640 120663
rect 539692 18624 539744 18630
rect 539692 18566 539744 18572
rect 539704 16574 539732 18566
rect 540992 16574 541020 244326
rect 543004 243024 543056 243030
rect 543004 242966 543056 242972
rect 542358 95840 542414 95849
rect 542358 95775 542414 95784
rect 542372 16574 542400 95775
rect 539704 16546 540376 16574
rect 540992 16546 542032 16574
rect 542372 16546 542768 16574
rect 538374 354 538486 480
rect 538232 326 538486 354
rect 538374 -960 538486 326
rect 539570 -960 539682 480
rect 540348 354 540376 16546
rect 542004 480 542032 16546
rect 540766 354 540878 480
rect 540348 326 540878 354
rect 540766 -960 540878 326
rect 541962 -960 542074 480
rect 542740 354 542768 16546
rect 543016 3194 543044 242966
rect 543738 148336 543794 148345
rect 543738 148271 543794 148280
rect 543752 16574 543780 148271
rect 547144 141432 547196 141438
rect 547144 141374 547196 141380
rect 543752 16546 544424 16574
rect 543004 3188 543056 3194
rect 543004 3130 543056 3136
rect 544396 480 544424 16546
rect 546684 7608 546736 7614
rect 546684 7550 546736 7556
rect 545488 3188 545540 3194
rect 545488 3130 545540 3136
rect 545500 480 545528 3130
rect 546696 480 546724 7550
rect 547156 4146 547184 141374
rect 547984 16574 548012 324294
rect 550640 152516 550692 152522
rect 550640 152458 550692 152464
rect 549258 93120 549314 93129
rect 549258 93055 549314 93064
rect 549272 16574 549300 93055
rect 550652 16574 550680 152458
rect 547984 16546 548656 16574
rect 549272 16546 550312 16574
rect 550652 16546 551048 16574
rect 547144 4140 547196 4146
rect 547144 4082 547196 4088
rect 547880 4140 547932 4146
rect 547880 4082 547932 4088
rect 547892 480 547920 4082
rect 543158 354 543270 480
rect 542740 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 548628 354 548656 16546
rect 550284 480 550312 16546
rect 549046 354 549158 480
rect 548628 326 549158 354
rect 549046 -960 549158 326
rect 550242 -960 550354 480
rect 551020 354 551048 16546
rect 552032 6914 552060 333950
rect 552662 311128 552718 311137
rect 552662 311063 552718 311072
rect 552676 16574 552704 311063
rect 570602 305008 570658 305017
rect 570602 304943 570658 304952
rect 565820 302932 565872 302938
rect 565820 302874 565872 302880
rect 558920 244316 558972 244322
rect 558920 244258 558972 244264
rect 557540 153876 557592 153882
rect 557540 153818 557592 153824
rect 554780 138712 554832 138718
rect 554780 138654 554832 138660
rect 553400 91792 553452 91798
rect 553400 91734 553452 91740
rect 553412 16574 553440 91734
rect 552676 16546 552796 16574
rect 553412 16546 553808 16574
rect 552032 6886 552704 6914
rect 552676 480 552704 6886
rect 552768 3194 552796 16546
rect 552756 3188 552808 3194
rect 552756 3130 552808 3136
rect 553780 480 553808 16546
rect 551438 354 551550 480
rect 551020 326 551550 354
rect 551438 -960 551550 326
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554792 354 554820 138654
rect 556252 90364 556304 90370
rect 556252 90306 556304 90312
rect 556264 16574 556292 90306
rect 557552 16574 557580 153818
rect 558932 16574 558960 244258
rect 563060 242956 563112 242962
rect 563060 242898 563112 242904
rect 561680 146940 561732 146946
rect 561680 146882 561732 146888
rect 560300 89004 560352 89010
rect 560300 88946 560352 88952
rect 560312 16574 560340 88946
rect 561692 16574 561720 146882
rect 556264 16546 556936 16574
rect 557552 16546 558592 16574
rect 558932 16546 559328 16574
rect 560312 16546 560432 16574
rect 561692 16546 562088 16574
rect 556160 3188 556212 3194
rect 556160 3130 556212 3136
rect 556172 480 556200 3130
rect 554934 354 555046 480
rect 554792 326 555046 354
rect 554934 -960 555046 326
rect 556130 -960 556242 480
rect 556908 354 556936 16546
rect 558564 480 558592 16546
rect 557326 354 557438 480
rect 556908 326 557438 354
rect 557326 -960 557438 326
rect 558522 -960 558634 480
rect 559300 354 559328 16546
rect 559718 354 559830 480
rect 559300 326 559830 354
rect 560404 354 560432 16546
rect 562060 480 562088 16546
rect 560822 354 560934 480
rect 560404 326 560934 354
rect 559718 -960 559830 326
rect 560822 -960 560934 326
rect 562018 -960 562130 480
rect 563072 354 563100 242898
rect 564440 136672 564492 136678
rect 564440 136614 564492 136620
rect 564452 3534 564480 136614
rect 564532 87644 564584 87650
rect 564532 87586 564584 87592
rect 564440 3528 564492 3534
rect 564440 3470 564492 3476
rect 564544 3346 564572 87586
rect 565832 16574 565860 302874
rect 569960 290488 570012 290494
rect 569960 290430 570012 290436
rect 567200 86284 567252 86290
rect 567200 86226 567252 86232
rect 567212 16574 567240 86226
rect 569224 84856 569276 84862
rect 569224 84798 569276 84804
rect 568580 36576 568632 36582
rect 568580 36518 568632 36524
rect 568592 16574 568620 36518
rect 565832 16546 566872 16574
rect 567212 16546 567608 16574
rect 568592 16546 568712 16574
rect 565268 3528 565320 3534
rect 565268 3470 565320 3476
rect 564452 3318 564572 3346
rect 564452 480 564480 3318
rect 563214 354 563326 480
rect 563072 326 563326 354
rect 563214 -960 563326 326
rect 564410 -960 564522 480
rect 565280 354 565308 3470
rect 566844 480 566872 16546
rect 565606 354 565718 480
rect 565280 326 565718 354
rect 565606 -960 565718 326
rect 566802 -960 566914 480
rect 567580 354 567608 16546
rect 567998 354 568110 480
rect 567580 326 568110 354
rect 568684 354 568712 16546
rect 569236 3194 569264 84798
rect 569972 16574 570000 290430
rect 569972 16546 570368 16574
rect 569224 3188 569276 3194
rect 569224 3130 569276 3136
rect 570340 480 570368 16546
rect 570616 3398 570644 304943
rect 577516 193186 577544 386951
rect 580276 378457 580304 399434
rect 580262 378448 580318 378457
rect 580262 378383 580318 378392
rect 577596 369912 577648 369918
rect 577596 369854 577648 369860
rect 577608 325514 577636 369854
rect 580632 369232 580684 369238
rect 580632 369174 580684 369180
rect 580356 369164 580408 369170
rect 580356 369106 580408 369112
rect 580262 366480 580318 366489
rect 580262 366415 580318 366424
rect 580172 365696 580224 365702
rect 580172 365638 580224 365644
rect 580184 365129 580212 365638
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 577596 325508 577648 325514
rect 577596 325450 577648 325456
rect 579620 313268 579672 313274
rect 579620 313210 579672 313216
rect 579632 312089 579660 313210
rect 579618 312080 579674 312089
rect 579618 312015 579674 312024
rect 580172 298784 580224 298790
rect 580170 298752 580172 298761
rect 580224 298752 580226 298761
rect 580170 298687 580226 298696
rect 577596 295384 577648 295390
rect 577596 295326 577648 295332
rect 577608 245614 577636 295326
rect 577596 245608 577648 245614
rect 579620 245608 579672 245614
rect 577596 245550 577648 245556
rect 579618 245576 579620 245585
rect 579672 245576 579674 245585
rect 579618 245511 579674 245520
rect 579620 233232 579672 233238
rect 579620 233174 579672 233180
rect 579632 232393 579660 233174
rect 579618 232384 579674 232393
rect 579618 232319 579674 232328
rect 579618 209128 579674 209137
rect 579618 209063 579674 209072
rect 579632 205737 579660 209063
rect 579618 205728 579674 205737
rect 579618 205663 579674 205672
rect 577504 193180 577556 193186
rect 577504 193122 577556 193128
rect 579620 193180 579672 193186
rect 579620 193122 579672 193128
rect 579632 192545 579660 193122
rect 579618 192536 579674 192545
rect 579618 192471 579674 192480
rect 579896 153196 579948 153202
rect 579896 153138 579948 153144
rect 579908 152697 579936 153138
rect 579894 152688 579950 152697
rect 579894 152623 579950 152632
rect 580276 139369 580304 366415
rect 580368 258913 580396 369106
rect 580538 366344 580594 366353
rect 580538 366279 580594 366288
rect 580446 364984 580502 364993
rect 580446 364919 580502 364928
rect 580354 258904 580410 258913
rect 580354 258839 580410 258848
rect 580354 200696 580410 200705
rect 580354 200631 580410 200640
rect 580262 139360 580318 139369
rect 580262 139295 580318 139304
rect 571984 135924 572036 135930
rect 571984 135866 572036 135872
rect 570604 3392 570656 3398
rect 570604 3334 570656 3340
rect 571996 3330 572024 135866
rect 575480 134564 575532 134570
rect 575480 134506 575532 134512
rect 574100 83496 574152 83502
rect 574100 83438 574152 83444
rect 574112 16574 574140 83438
rect 575492 16574 575520 134506
rect 580172 113144 580224 113150
rect 580172 113086 580224 113092
rect 580184 112849 580212 113086
rect 580170 112840 580226 112849
rect 580170 112775 580226 112784
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580262 100056 580318 100065
rect 580262 99991 580318 100000
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580276 86193 580304 99991
rect 580262 86184 580318 86193
rect 580262 86119 580318 86128
rect 578240 80708 578292 80714
rect 578240 80650 578292 80656
rect 578252 16574 578280 80650
rect 580262 71088 580318 71097
rect 580262 71023 580318 71032
rect 580276 46345 580304 71023
rect 580262 46336 580318 46345
rect 580262 46271 580318 46280
rect 580080 20664 580132 20670
rect 580080 20606 580132 20612
rect 580092 19825 580120 20606
rect 580078 19816 580134 19825
rect 580078 19751 580134 19760
rect 574112 16546 575152 16574
rect 575492 16546 575888 16574
rect 578252 16546 578648 16574
rect 573916 3664 573968 3670
rect 573916 3606 573968 3612
rect 571984 3324 572036 3330
rect 571984 3266 572036 3272
rect 572720 3324 572772 3330
rect 572720 3266 572772 3272
rect 571524 3188 571576 3194
rect 571524 3130 571576 3136
rect 571536 480 571564 3130
rect 572732 480 572760 3266
rect 573928 480 573956 3606
rect 575124 480 575152 16546
rect 569102 354 569214 480
rect 568684 326 569214 354
rect 567998 -960 568110 326
rect 569102 -960 569214 326
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 575860 354 575888 16546
rect 577412 3392 577464 3398
rect 577412 3334 577464 3340
rect 577424 480 577452 3334
rect 578620 480 578648 16546
rect 580368 6633 580396 200631
rect 580460 179217 580488 364919
rect 580552 219065 580580 366279
rect 580644 272241 580672 369174
rect 580736 351937 580764 400823
rect 580722 351928 580778 351937
rect 580722 351863 580778 351872
rect 580724 325508 580776 325514
rect 580724 325450 580776 325456
rect 580736 325281 580764 325450
rect 580722 325272 580778 325281
rect 580722 325207 580778 325216
rect 580630 272232 580686 272241
rect 580630 272167 580686 272176
rect 580538 219056 580594 219065
rect 580538 218991 580594 219000
rect 580538 209264 580594 209273
rect 580538 209199 580594 209208
rect 580446 179208 580502 179217
rect 580446 179143 580502 179152
rect 580552 126041 580580 209199
rect 580722 208992 580778 209001
rect 580722 208927 580778 208936
rect 580736 165889 580764 208927
rect 580722 165880 580778 165889
rect 580722 165815 580778 165824
rect 580538 126032 580594 126041
rect 580538 125967 580594 125976
rect 580354 6624 580410 6633
rect 580354 6559 580410 6568
rect 576278 354 576390 480
rect 575860 326 576390 354
rect 576278 -960 576390 326
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3422 671200 3478 671256
rect 2778 658144 2834 658200
rect 3422 632068 3424 632088
rect 3424 632068 3476 632088
rect 3476 632068 3478 632088
rect 3422 632032 3478 632068
rect 3422 619112 3478 619168
rect 3330 579944 3386 580000
rect 3238 566888 3294 566944
rect 3330 553832 3386 553888
rect 2962 527856 3018 527912
rect 3054 501744 3110 501800
rect 3054 475632 3110 475688
rect 3054 449520 3110 449576
rect 3514 606056 3570 606112
rect 3514 514820 3570 514856
rect 3514 514800 3516 514820
rect 3516 514800 3568 514820
rect 3568 514800 3570 514820
rect 3514 462596 3570 462632
rect 3514 462576 3516 462596
rect 3516 462576 3568 462596
rect 3568 462576 3570 462596
rect 3514 423544 3570 423600
rect 3422 410488 3478 410544
rect 3422 397468 3424 397488
rect 3424 397468 3476 397488
rect 3476 397468 3478 397488
rect 3422 397432 3478 397468
rect 3422 371320 3478 371376
rect 3146 358400 3202 358456
rect 3330 345344 3386 345400
rect 3422 319232 3478 319288
rect 4066 306176 4122 306232
rect 3422 293120 3478 293176
rect 3054 267144 3110 267200
rect 3422 254088 3478 254144
rect 3330 241032 3386 241088
rect 153014 241848 153070 241904
rect 151726 241712 151782 241768
rect 151634 241576 151690 241632
rect 150346 229744 150402 229800
rect 3422 214920 3478 214976
rect 3330 201864 3386 201920
rect 3146 188808 3202 188864
rect 3330 162832 3386 162888
rect 3146 110608 3202 110664
rect 3054 58520 3110 58576
rect 2870 32408 2926 32464
rect 3698 149776 3754 149832
rect 3606 136720 3662 136776
rect 3514 97552 3570 97608
rect 3514 84632 3570 84688
rect 3514 71576 3570 71632
rect 3514 45500 3516 45520
rect 3516 45500 3568 45520
rect 3568 45500 3570 45520
rect 3514 45464 3570 45500
rect 3422 19352 3478 19408
rect 3422 6432 3478 6488
rect 18602 145560 18658 145616
rect 20718 122032 20774 122088
rect 28998 153720 29054 153776
rect 34518 151000 34574 151056
rect 36542 130328 36598 130384
rect 44270 113736 44326 113792
rect 51078 151136 51134 151192
rect 53838 149640 53894 149696
rect 55218 131688 55274 131744
rect 59358 137264 59414 137320
rect 71042 153856 71098 153912
rect 64878 151272 64934 151328
rect 75918 148280 75974 148336
rect 80702 135904 80758 135960
rect 80058 126248 80114 126304
rect 84198 130464 84254 130520
rect 89718 152360 89774 152416
rect 100758 155216 100814 155272
rect 103518 146920 103574 146976
rect 110418 149776 110474 149832
rect 120722 147056 120778 147112
rect 117962 144064 118018 144120
rect 112442 122168 112498 122224
rect 126978 153992 127034 154048
rect 129002 136040 129058 136096
rect 129738 126384 129794 126440
rect 135350 149912 135406 149968
rect 136638 148416 136694 148472
rect 140778 139984 140834 140040
rect 147678 141344 147734 141400
rect 149702 151000 149758 151056
rect 151266 158888 151322 158944
rect 151542 158888 151598 158944
rect 152922 240760 152978 240816
rect 152554 159568 152610 159624
rect 152922 159568 152978 159624
rect 152830 156712 152886 156768
rect 152554 152360 152610 152416
rect 154118 220088 154174 220144
rect 153106 147464 153162 147520
rect 154118 147600 154174 147656
rect 157246 240896 157302 240952
rect 157062 240624 157118 240680
rect 155498 239400 155554 239456
rect 154578 153040 154634 153096
rect 155314 160112 155370 160168
rect 155774 239672 155830 239728
rect 155682 159840 155738 159896
rect 155590 156984 155646 157040
rect 155498 153856 155554 153912
rect 155314 153720 155370 153776
rect 155866 239536 155922 239592
rect 156510 156576 156566 156632
rect 155774 149640 155830 149696
rect 156694 159976 156750 160032
rect 156970 160384 157026 160440
rect 156878 159296 156934 159352
rect 156786 158752 156842 158808
rect 156878 156576 156934 156632
rect 158350 235320 158406 235376
rect 158258 228248 158314 228304
rect 158166 221448 158222 221504
rect 157798 211112 157854 211168
rect 157890 158480 157946 158536
rect 157338 157800 157394 157856
rect 157798 157800 157854 157856
rect 157246 157256 157302 157312
rect 157430 157392 157486 157448
rect 157338 155216 157394 155272
rect 157430 153992 157486 154048
rect 157338 153720 157394 153776
rect 156970 151136 157026 151192
rect 158258 160248 158314 160304
rect 158166 157528 158222 157584
rect 158074 157256 158130 157312
rect 158166 153040 158222 153096
rect 159822 231648 159878 231704
rect 159546 225528 159602 225584
rect 159362 160520 159418 160576
rect 158718 159160 158774 159216
rect 158626 158072 158682 158128
rect 158350 157392 158406 157448
rect 158258 148280 158314 148336
rect 159454 158616 159510 158672
rect 159730 157936 159786 157992
rect 160558 159704 160614 159760
rect 160006 158616 160062 158672
rect 160006 157664 160062 157720
rect 159822 156848 159878 156904
rect 161110 161880 161166 161936
rect 159362 151272 159418 151328
rect 160098 144744 160154 144800
rect 161386 144744 161442 144800
rect 162122 159840 162178 159896
rect 162582 211112 162638 211168
rect 164330 211248 164386 211304
rect 164882 211112 164938 211168
rect 165802 275168 165858 275224
rect 165434 211112 165490 211168
rect 168470 278024 168526 278080
rect 171322 287680 171378 287736
rect 165342 209616 165398 209672
rect 166814 209616 166870 209672
rect 180890 212064 180946 212120
rect 184202 289720 184258 289776
rect 186502 289584 186558 289640
rect 186318 289176 186374 289232
rect 185030 289040 185086 289096
rect 186686 289448 186742 289504
rect 187330 210024 187386 210080
rect 187790 289312 187846 289368
rect 184846 209616 184902 209672
rect 188802 209616 188858 209672
rect 189170 290672 189226 290728
rect 192022 290536 192078 290592
rect 190550 289992 190606 290048
rect 191838 289856 191894 289912
rect 190642 276664 190698 276720
rect 190734 243480 190790 243536
rect 192114 286320 192170 286376
rect 192482 232736 192538 232792
rect 193770 233144 193826 233200
rect 196254 210024 196310 210080
rect 196990 209616 197046 209672
rect 198462 209616 198518 209672
rect 171966 209480 172022 209536
rect 184754 209480 184810 209536
rect 188894 209480 188950 209536
rect 191746 209480 191802 209536
rect 192942 209480 192998 209536
rect 194414 209480 194470 209536
rect 195886 209480 195942 209536
rect 196898 209480 196954 209536
rect 197266 209480 197322 209536
rect 199566 209616 199622 209672
rect 201314 226208 201370 226264
rect 202786 321544 202842 321600
rect 199842 209616 199898 209672
rect 199934 209480 199990 209536
rect 202510 231648 202566 231704
rect 202786 219272 202842 219328
rect 202786 218864 202842 218920
rect 203982 235728 204038 235784
rect 203982 235456 204038 235512
rect 204902 307536 204958 307592
rect 204902 238448 204958 238504
rect 205270 230016 205326 230072
rect 205454 231784 205510 231840
rect 205362 228928 205418 228984
rect 205362 228248 205418 228304
rect 206466 304272 206522 304328
rect 206374 240896 206430 240952
rect 206650 238176 206706 238232
rect 206650 237632 206706 237688
rect 217966 321000 218022 321056
rect 206926 320864 206982 320920
rect 206834 316648 206890 316704
rect 210974 320728 211030 320784
rect 207938 319504 207994 319560
rect 207846 239400 207902 239456
rect 208030 319368 208086 319424
rect 205638 223488 205694 223544
rect 206650 223488 206706 223544
rect 207570 170312 207626 170368
rect 163042 159840 163098 159896
rect 162950 159704 163006 159760
rect 162950 159024 163006 159080
rect 163042 158616 163098 158672
rect 163410 159840 163466 159896
rect 163594 159840 163650 159896
rect 163410 159568 163466 159624
rect 163502 157972 163504 157992
rect 163504 157972 163556 157992
rect 163556 157972 163558 157992
rect 163502 157936 163558 157972
rect 163502 157428 163504 157448
rect 163504 157428 163556 157448
rect 163556 157428 163558 157448
rect 163502 157392 163558 157428
rect 163502 156460 163558 156496
rect 163502 156440 163504 156460
rect 163504 156440 163556 156460
rect 163556 156440 163558 156460
rect 163686 157800 163742 157856
rect 163870 158480 163926 158536
rect 163962 158344 164018 158400
rect 164238 159840 164294 159896
rect 164330 158752 164386 158808
rect 164238 158344 164294 158400
rect 164330 158208 164386 158264
rect 164146 157412 164202 157448
rect 164330 157800 164386 157856
rect 164146 157392 164148 157412
rect 164148 157392 164200 157412
rect 164200 157392 164202 157412
rect 164054 157120 164110 157176
rect 164698 159874 164754 159930
rect 164698 158616 164754 158672
rect 164606 158480 164662 158536
rect 164606 157936 164662 157992
rect 164882 158480 164938 158536
rect 164882 158344 164938 158400
rect 164790 157256 164846 157312
rect 165158 159704 165214 159760
rect 165342 159840 165398 159896
rect 165618 159840 165674 159896
rect 165158 158888 165214 158944
rect 165158 158480 165214 158536
rect 165250 157800 165306 157856
rect 165526 159704 165582 159760
rect 165618 159568 165674 159624
rect 165618 158888 165674 158944
rect 165710 158616 165766 158672
rect 165894 159024 165950 159080
rect 166262 159840 166318 159896
rect 166170 159704 166226 159760
rect 166354 159568 166410 159624
rect 166446 159160 166502 159216
rect 166354 158888 166410 158944
rect 165986 156984 166042 157040
rect 166262 158616 166318 158672
rect 166262 158072 166318 158128
rect 166262 157528 166318 157584
rect 166722 159840 166778 159896
rect 166814 159704 166870 159760
rect 166814 158616 166870 158672
rect 166722 158480 166778 158536
rect 167182 159840 167238 159896
rect 167182 159296 167238 159352
rect 167090 158616 167146 158672
rect 166998 157664 167054 157720
rect 167458 159840 167514 159896
rect 167642 159840 167698 159896
rect 167458 158344 167514 158400
rect 167918 159568 167974 159624
rect 168010 156576 168066 156632
rect 168286 159840 168342 159896
rect 168194 159704 168250 159760
rect 168470 159704 168526 159760
rect 168378 158344 168434 158400
rect 168286 158228 168342 158264
rect 168286 158208 168288 158228
rect 168288 158208 168340 158228
rect 168340 158208 168342 158228
rect 168562 158888 168618 158944
rect 168470 158208 168526 158264
rect 168470 158072 168526 158128
rect 168470 157664 168526 157720
rect 168746 159840 168802 159896
rect 168654 158616 168710 158672
rect 169022 159704 169078 159760
rect 168930 158072 168986 158128
rect 168838 156712 168894 156768
rect 169206 159840 169262 159896
rect 169298 159568 169354 159624
rect 169482 159840 169538 159896
rect 169390 159432 169446 159488
rect 169390 158616 169446 158672
rect 169482 158344 169538 158400
rect 169850 159432 169906 159488
rect 170126 157256 170182 157312
rect 170402 159840 170458 159896
rect 170586 159704 170642 159760
rect 170770 159704 170826 159760
rect 170586 158888 170642 158944
rect 170494 158208 170550 158264
rect 170954 159840 171010 159896
rect 170954 159740 170956 159760
rect 170956 159740 171008 159760
rect 171008 159740 171010 159760
rect 170954 159704 171010 159740
rect 171138 159840 171194 159896
rect 170678 158072 170734 158128
rect 171046 158616 171102 158672
rect 170862 158208 170918 158264
rect 170770 157528 170826 157584
rect 170954 158072 171010 158128
rect 171230 159568 171286 159624
rect 171414 159704 171470 159760
rect 171322 158616 171378 158672
rect 171506 159568 171562 159624
rect 171782 159840 171838 159896
rect 171598 158344 171654 158400
rect 172150 158616 172206 158672
rect 171966 158072 172022 158128
rect 172610 159840 172666 159896
rect 172702 159704 172758 159760
rect 172518 159568 172574 159624
rect 172886 159840 172942 159896
rect 172702 158208 172758 158264
rect 172242 153040 172298 153096
rect 173254 159704 173310 159760
rect 173070 158616 173126 158672
rect 173438 159704 173494 159760
rect 173438 159568 173494 159624
rect 173438 158888 173494 158944
rect 173346 157256 173402 157312
rect 173162 149096 173218 149152
rect 173714 159840 173770 159896
rect 173990 159840 174046 159896
rect 173898 159568 173954 159624
rect 173990 158344 174046 158400
rect 173990 158208 174046 158264
rect 174266 159704 174322 159760
rect 174542 159840 174598 159896
rect 174450 157664 174506 157720
rect 174818 159704 174874 159760
rect 174726 159024 174782 159080
rect 174818 158752 174874 158808
rect 174634 158616 174690 158672
rect 175094 159568 175150 159624
rect 175278 158344 175334 158400
rect 175278 158208 175334 158264
rect 175646 158616 175702 158672
rect 175922 159840 175978 159896
rect 175922 158208 175978 158264
rect 176382 158752 176438 158808
rect 176382 158616 176438 158672
rect 176382 157800 176438 157856
rect 176198 153040 176254 153096
rect 177026 159704 177082 159760
rect 177302 159840 177358 159896
rect 177210 157800 177266 157856
rect 177578 158616 177634 158672
rect 177762 158072 177818 158128
rect 177854 157936 177910 157992
rect 178958 159840 179014 159896
rect 179234 159704 179290 159760
rect 179142 158616 179198 158672
rect 179050 156576 179106 156632
rect 179786 159704 179842 159760
rect 180062 159840 180118 159896
rect 180338 159840 180394 159896
rect 180338 159704 180394 159760
rect 180614 159840 180670 159896
rect 179418 98640 179474 98696
rect 180890 159704 180946 159760
rect 181166 159840 181222 159896
rect 181442 158616 181498 158672
rect 181718 159704 181774 159760
rect 181902 159840 181958 159896
rect 181902 158888 181958 158944
rect 181994 158072 182050 158128
rect 182270 159840 182326 159896
rect 182546 158616 182602 158672
rect 182822 159840 182878 159896
rect 182822 158072 182878 158128
rect 183098 158616 183154 158672
rect 183282 159840 183338 159896
rect 183374 159704 183430 159760
rect 183466 158072 183522 158128
rect 183926 159840 183982 159896
rect 184202 159840 184258 159896
rect 184478 159704 184534 159760
rect 184754 159432 184810 159488
rect 185030 158616 185086 158672
rect 185858 158616 185914 158672
rect 186318 158752 186374 158808
rect 186134 141208 186190 141264
rect 186134 140800 186190 140856
rect 186686 158616 186742 158672
rect 186962 158072 187018 158128
rect 187238 158616 187294 158672
rect 187514 158616 187570 158672
rect 188066 158616 188122 158672
rect 188342 159840 188398 159896
rect 188434 159024 188490 159080
rect 188434 158752 188490 158808
rect 188618 158616 188674 158672
rect 188986 157256 189042 157312
rect 189170 158616 189226 158672
rect 189722 159840 189778 159896
rect 189630 159704 189686 159760
rect 189998 158616 190054 158672
rect 190274 158616 190330 158672
rect 190550 158888 190606 158944
rect 190458 158072 190514 158128
rect 189722 141480 189778 141536
rect 190826 159840 190882 159896
rect 190826 155760 190882 155816
rect 191102 159704 191158 159760
rect 191378 159840 191434 159896
rect 191654 159432 191710 159488
rect 191654 158072 191710 158128
rect 191930 158616 191986 158672
rect 192206 159704 192262 159760
rect 192022 152632 192078 152688
rect 192482 159840 192538 159896
rect 192390 157528 192446 157584
rect 192390 157256 192446 157312
rect 192482 156032 192538 156088
rect 192758 159840 192814 159896
rect 193034 158616 193090 158672
rect 193310 158072 193366 158128
rect 193126 156032 193182 156088
rect 193586 159840 193642 159896
rect 193402 155216 193458 155272
rect 193310 152088 193366 152144
rect 193586 152088 193642 152144
rect 194138 158616 194194 158672
rect 194414 159840 194470 159896
rect 194506 156712 194562 156768
rect 194690 158072 194746 158128
rect 194966 159840 195022 159896
rect 195242 159704 195298 159760
rect 194966 149912 195022 149968
rect 195610 158616 195666 158672
rect 195794 159840 195850 159896
rect 195886 158616 195942 158672
rect 193862 28192 193918 28248
rect 196070 158616 196126 158672
rect 196070 158072 196126 158128
rect 196346 159840 196402 159896
rect 196622 159704 196678 159760
rect 196622 151408 196678 151464
rect 196898 159840 196954 159896
rect 196806 155896 196862 155952
rect 197174 159840 197230 159896
rect 197082 153584 197138 153640
rect 197266 158616 197322 158672
rect 196346 147056 196402 147112
rect 197082 144336 197138 144392
rect 196622 17176 196678 17232
rect 197910 159840 197966 159896
rect 198002 159704 198058 159760
rect 197910 159432 197966 159488
rect 197910 158344 197966 158400
rect 197910 158072 197966 158128
rect 197910 155352 197966 155408
rect 197910 154944 197966 155000
rect 197910 150048 197966 150104
rect 198278 158616 198334 158672
rect 198370 158344 198426 158400
rect 198554 159840 198610 159896
rect 198462 156440 198518 156496
rect 198830 159840 198886 159896
rect 198830 157800 198886 157856
rect 197542 139304 197598 139360
rect 198646 139304 198702 139360
rect 197358 116456 197414 116512
rect 199106 159840 199162 159896
rect 199198 158616 199254 158672
rect 199106 157936 199162 157992
rect 199382 159840 199438 159896
rect 199382 159740 199384 159760
rect 199384 159740 199436 159760
rect 199436 159740 199438 159760
rect 199382 159704 199438 159740
rect 199014 148824 199070 148880
rect 199658 154672 199714 154728
rect 199566 151136 199622 151192
rect 199474 148688 199530 148744
rect 199842 158616 199898 158672
rect 200118 159296 200174 159352
rect 200210 158616 200266 158672
rect 199934 158344 199990 158400
rect 200394 158888 200450 158944
rect 200026 157936 200082 157992
rect 200302 157936 200358 157992
rect 199934 157800 199990 157856
rect 199842 154536 199898 154592
rect 200302 152496 200358 152552
rect 200670 157256 200726 157312
rect 200302 152224 200358 152280
rect 200946 158616 201002 158672
rect 201038 158344 201094 158400
rect 200854 156848 200910 156904
rect 201038 156848 201094 156904
rect 201314 159840 201370 159896
rect 201406 159024 201462 159080
rect 201498 158752 201554 158808
rect 201406 158344 201462 158400
rect 201130 151544 201186 151600
rect 201314 157392 201370 157448
rect 201038 150184 201094 150240
rect 201222 144336 201278 144392
rect 200210 144064 200266 144120
rect 201130 144064 201186 144120
rect 201866 156032 201922 156088
rect 201682 154808 201738 154864
rect 202142 158344 202198 158400
rect 202326 159840 202382 159896
rect 202326 159432 202382 159488
rect 202418 158616 202474 158672
rect 202694 157936 202750 157992
rect 202694 154808 202750 154864
rect 202878 159432 202934 159488
rect 202970 158616 203026 158672
rect 202878 155488 202934 155544
rect 203154 154400 203210 154456
rect 203522 159840 203578 159896
rect 203430 159704 203486 159760
rect 203798 159840 203854 159896
rect 203614 154672 203670 154728
rect 202694 144336 202750 144392
rect 203798 151680 203854 151736
rect 204074 159704 204130 159760
rect 203982 158616 204038 158672
rect 204350 158616 204406 158672
rect 204258 158344 204314 158400
rect 203706 144336 203762 144392
rect 203706 143928 203762 143984
rect 204166 155488 204222 155544
rect 204074 150320 204130 150376
rect 204626 159840 204682 159896
rect 204534 155216 204590 155272
rect 204902 159024 204958 159080
rect 204718 148960 204774 149016
rect 205178 159840 205234 159896
rect 204718 139304 204774 139360
rect 205178 158344 205234 158400
rect 205454 159704 205510 159760
rect 205638 159704 205694 159760
rect 205454 155216 205510 155272
rect 205362 154264 205418 154320
rect 205178 151272 205234 151328
rect 204994 139168 205050 139224
rect 206282 159840 206338 159896
rect 206190 159024 206246 159080
rect 206558 159840 206614 159896
rect 206834 159840 206890 159896
rect 206558 147600 206614 147656
rect 207018 158616 207074 158672
rect 207294 159840 207350 159896
rect 207386 159704 207442 159760
rect 207110 158072 207166 158128
rect 208950 238176 209006 238232
rect 208766 234504 208822 234560
rect 208490 233688 208546 233744
rect 208766 233552 208822 233608
rect 208306 224304 208362 224360
rect 207754 202136 207810 202192
rect 207846 188264 207902 188320
rect 207754 166368 207810 166424
rect 207662 166096 207718 166152
rect 207386 157800 207442 157856
rect 207294 157664 207350 157720
rect 207662 158208 207718 158264
rect 207478 155760 207534 155816
rect 207938 184184 207994 184240
rect 208766 173576 208822 173632
rect 208030 173440 208086 173496
rect 208122 166368 208178 166424
rect 208214 161336 208270 161392
rect 208214 160248 208270 160304
rect 208214 158072 208270 158128
rect 208398 160656 208454 160712
rect 208398 160112 208454 160168
rect 208122 157664 208178 157720
rect 208306 157800 208362 157856
rect 208490 157936 208546 157992
rect 208398 155896 208454 155952
rect 209318 304680 209374 304736
rect 209594 240760 209650 240816
rect 210146 306992 210202 307048
rect 209686 235592 209742 235648
rect 209410 234504 209466 234560
rect 210330 239672 210386 239728
rect 210146 234368 210202 234424
rect 209226 173576 209282 173632
rect 209134 159568 209190 159624
rect 209410 158344 209466 158400
rect 208490 153584 208546 153640
rect 210330 157528 210386 157584
rect 210514 158072 210570 158128
rect 210790 239672 210846 239728
rect 210790 239264 210846 239320
rect 215022 319912 215078 319968
rect 213090 319640 213146 319696
rect 210974 236544 211030 236600
rect 210790 156440 210846 156496
rect 210422 155624 210478 155680
rect 210422 154808 210478 154864
rect 211618 297336 211674 297392
rect 212078 307400 212134 307456
rect 211710 239128 211766 239184
rect 211710 154944 211766 155000
rect 211158 149504 211214 149560
rect 212078 238312 212134 238368
rect 212354 315288 212410 315344
rect 212170 236408 212226 236464
rect 213090 239536 213146 239592
rect 213090 156712 213146 156768
rect 212170 153992 212226 154048
rect 212538 151000 212594 151056
rect 211894 144608 211950 144664
rect 213458 240352 213514 240408
rect 213458 152360 213514 152416
rect 213918 156576 213974 156632
rect 213366 147328 213422 147384
rect 214654 237088 214710 237144
rect 214838 235320 214894 235376
rect 215114 236816 215170 236872
rect 215022 153720 215078 153776
rect 216126 307264 216182 307320
rect 216126 236952 216182 237008
rect 215850 148552 215906 148608
rect 215298 147736 215354 147792
rect 215850 147736 215906 147792
rect 214746 147192 214802 147248
rect 217414 241168 217470 241224
rect 217782 315424 217838 315480
rect 217506 238720 217562 238776
rect 217414 237224 217470 237280
rect 217414 236816 217470 236872
rect 216678 139984 216734 140040
rect 218058 291760 218114 291816
rect 217782 237224 217838 237280
rect 217690 156984 217746 157040
rect 218978 307128 219034 307184
rect 218610 237224 218666 237280
rect 218702 232328 218758 232384
rect 218058 201320 218114 201376
rect 218518 201320 218574 201376
rect 218058 200640 218114 200696
rect 217598 152768 217654 152824
rect 217414 141344 217470 141400
rect 218886 239944 218942 240000
rect 219346 291760 219402 291816
rect 219990 291624 220046 291680
rect 219990 239536 220046 239592
rect 219898 238992 219954 239048
rect 220082 228248 220138 228304
rect 222106 372816 222162 372872
rect 222014 312432 222070 312488
rect 220726 290400 220782 290456
rect 221186 241848 221242 241904
rect 220634 238856 220690 238912
rect 220450 236136 220506 236192
rect 220450 232736 220506 232792
rect 220910 239264 220966 239320
rect 221462 240896 221518 240952
rect 221462 239400 221518 239456
rect 221462 233688 221518 233744
rect 220174 152496 220230 152552
rect 221830 246336 221886 246392
rect 224866 370096 224922 370152
rect 224222 369960 224278 370016
rect 222014 246336 222070 246392
rect 228362 369280 228418 369336
rect 225602 369144 225658 369200
rect 225694 321136 225750 321192
rect 224222 290128 224278 290184
rect 224222 289856 224278 289912
rect 225786 317464 225842 317520
rect 227166 318552 227222 318608
rect 227166 301552 227222 301608
rect 225786 295296 225842 295352
rect 226154 291216 226210 291272
rect 227718 291760 227774 291816
rect 227626 290400 227682 290456
rect 228362 291352 228418 291408
rect 229926 368600 229982 368656
rect 230018 323584 230074 323640
rect 233330 318416 233386 318472
rect 233330 315560 233386 315616
rect 231582 289856 231638 289912
rect 238574 315968 238630 316024
rect 238574 306448 238630 306504
rect 238758 314064 238814 314120
rect 234158 290128 234214 290184
rect 234158 289856 234214 289912
rect 238666 306176 238722 306232
rect 238666 296792 238722 296848
rect 238666 296656 238722 296712
rect 238666 290128 238722 290184
rect 240874 292576 240930 292632
rect 242254 371320 242310 371376
rect 243542 360848 243598 360904
rect 242530 316920 242586 316976
rect 241058 289720 241114 289776
rect 242714 292440 242770 292496
rect 244278 290128 244334 290184
rect 248418 368872 248474 368928
rect 244830 289756 244832 289776
rect 244832 289756 244884 289776
rect 244884 289756 244886 289776
rect 244830 289720 244886 289756
rect 246394 353912 246450 353968
rect 246946 290672 247002 290728
rect 245474 289448 245530 289504
rect 247774 357992 247830 358048
rect 247682 291624 247738 291680
rect 247682 291216 247738 291272
rect 248234 291216 248290 291272
rect 253202 370368 253258 370424
rect 251822 369008 251878 369064
rect 250442 368328 250498 368384
rect 250442 363568 250498 363624
rect 249798 312704 249854 312760
rect 249706 291896 249762 291952
rect 251178 292168 251234 292224
rect 250442 291488 250498 291544
rect 250810 291080 250866 291136
rect 250626 289992 250682 290048
rect 251546 292032 251602 292088
rect 251914 362208 251970 362264
rect 252650 292304 252706 292360
rect 251914 292032 251970 292088
rect 251822 290536 251878 290592
rect 252098 290536 252154 290592
rect 251914 289856 251970 289912
rect 253294 292304 253350 292360
rect 266174 402056 266230 402112
rect 260746 396752 260802 396808
rect 260654 389952 260710 390008
rect 259274 388320 259330 388376
rect 259182 318008 259238 318064
rect 262034 389816 262090 389872
rect 260746 306856 260802 306912
rect 261942 310392 261998 310448
rect 266082 391176 266138 391232
rect 263322 314200 263378 314256
rect 264886 310120 264942 310176
rect 269026 400560 269082 400616
rect 266266 396616 266322 396672
rect 266174 307536 266230 307592
rect 267002 395392 267058 395448
rect 266358 317328 266414 317384
rect 267554 317328 267610 317384
rect 267370 313520 267426 313576
rect 267554 302776 267610 302832
rect 267094 291080 267150 291136
rect 248970 289584 249026 289640
rect 247038 289448 247094 289504
rect 247498 289312 247554 289368
rect 268658 394032 268714 394088
rect 268842 314472 268898 314528
rect 270314 397976 270370 398032
rect 269670 387096 269726 387152
rect 269578 385600 269634 385656
rect 269026 304816 269082 304872
rect 269026 304272 269082 304328
rect 267646 260072 267702 260128
rect 267554 241848 267610 241904
rect 222198 240624 222254 240680
rect 222290 240372 222346 240408
rect 222290 240352 222292 240372
rect 222292 240352 222344 240372
rect 222344 240352 222346 240372
rect 222106 240216 222162 240272
rect 222014 238040 222070 238096
rect 222014 233008 222070 233064
rect 221922 232328 221978 232384
rect 222198 239808 222254 239864
rect 222888 239844 222890 239864
rect 222890 239844 222942 239864
rect 222942 239844 222944 239864
rect 222382 239672 222438 239728
rect 222198 218728 222254 218784
rect 222888 239808 222944 239844
rect 223532 239808 223588 239864
rect 223118 238856 223174 238912
rect 220082 141208 220138 141264
rect 223486 239400 223542 239456
rect 223026 224304 223082 224360
rect 223486 238176 223542 238232
rect 223992 239808 224048 239864
rect 224130 239828 224186 239864
rect 224130 239808 224132 239828
rect 224132 239808 224184 239828
rect 224184 239808 224186 239828
rect 224360 239808 224416 239864
rect 223854 239692 223910 239728
rect 223854 239672 223856 239692
rect 223856 239672 223908 239692
rect 223908 239672 223910 239692
rect 223762 238892 223764 238912
rect 223764 238892 223816 238912
rect 223816 238892 223818 238912
rect 223762 238856 223818 238892
rect 223670 238448 223726 238504
rect 223670 238176 223726 238232
rect 223578 232600 223634 232656
rect 223762 219272 223818 219328
rect 223670 162152 223726 162208
rect 224912 239808 224968 239864
rect 224590 237632 224646 237688
rect 224498 229472 224554 229528
rect 224498 229336 224554 229392
rect 224314 226208 224370 226264
rect 224222 224440 224278 224496
rect 224038 159160 224094 159216
rect 225096 239808 225152 239864
rect 224406 170312 224462 170368
rect 225050 224168 225106 224224
rect 225326 239400 225382 239456
rect 225510 239264 225566 239320
rect 225786 239808 225842 239864
rect 225694 239556 225750 239592
rect 225694 239536 225696 239556
rect 225696 239536 225748 239556
rect 225748 239536 225750 239556
rect 225418 225936 225474 225992
rect 224958 217912 225014 217968
rect 225694 237496 225750 237552
rect 225602 231240 225658 231296
rect 224222 142704 224278 142760
rect 223026 138488 223082 138544
rect 225878 236272 225934 236328
rect 226568 239808 226624 239864
rect 226522 239536 226578 239592
rect 226614 238992 226670 239048
rect 226614 238176 226670 238232
rect 225786 224168 225842 224224
rect 225786 142568 225842 142624
rect 225878 140528 225934 140584
rect 226522 235864 226578 235920
rect 227028 239672 227084 239728
rect 226982 239400 227038 239456
rect 226982 238992 227038 239048
rect 226890 230424 226946 230480
rect 226798 217776 226854 217832
rect 227258 237768 227314 237824
rect 227672 239808 227728 239864
rect 227442 239692 227498 239728
rect 227442 239672 227444 239692
rect 227444 239672 227496 239692
rect 227496 239672 227498 239692
rect 227442 239436 227444 239456
rect 227444 239436 227496 239456
rect 227496 239436 227498 239456
rect 227442 239400 227498 239436
rect 227166 231784 227222 231840
rect 228132 239808 228188 239864
rect 228454 239808 228510 239864
rect 227994 239672 228050 239728
rect 228178 239264 228234 239320
rect 227994 238720 228050 238776
rect 227902 217504 227958 217560
rect 227718 211928 227774 211984
rect 228362 239672 228418 239728
rect 229236 239808 229292 239864
rect 228454 235728 228510 235784
rect 228638 239536 228694 239592
rect 228362 232464 228418 232520
rect 228178 228928 228234 228984
rect 228086 161744 228142 161800
rect 226430 120944 226486 121000
rect 228822 239400 228878 239456
rect 229282 239692 229338 239728
rect 229282 239672 229284 239692
rect 229284 239672 229336 239692
rect 229336 239672 229338 239692
rect 229282 239556 229338 239592
rect 229282 239536 229284 239556
rect 229284 239536 229336 239556
rect 229336 239536 229338 239556
rect 229190 238720 229246 238776
rect 229466 239672 229522 239728
rect 229788 239808 229844 239864
rect 229558 239536 229614 239592
rect 229374 238312 229430 238368
rect 228454 142840 228510 142896
rect 229742 238312 229798 238368
rect 229742 237904 229798 237960
rect 229650 237224 229706 237280
rect 229650 236136 229706 236192
rect 229650 236000 229706 236056
rect 230340 239808 230396 239864
rect 230294 239672 230350 239728
rect 230018 239400 230074 239456
rect 230294 239436 230296 239456
rect 230296 239436 230348 239456
rect 230348 239436 230350 239456
rect 230294 239400 230350 239436
rect 229926 236544 229982 236600
rect 230478 235728 230534 235784
rect 229742 227296 229798 227352
rect 229650 217368 229706 217424
rect 230018 188264 230074 188320
rect 230800 239844 230802 239864
rect 230802 239844 230854 239864
rect 230854 239844 230856 239864
rect 230800 239808 230856 239844
rect 231168 239808 231224 239864
rect 230202 220768 230258 220824
rect 231122 239672 231178 239728
rect 231904 239808 231960 239864
rect 230846 231104 230902 231160
rect 230478 220360 230534 220416
rect 230478 217640 230534 217696
rect 230570 217232 230626 217288
rect 231122 238720 231178 238776
rect 231122 238176 231178 238232
rect 231490 239672 231546 239728
rect 231766 239572 231768 239592
rect 231768 239572 231820 239592
rect 231820 239572 231822 239592
rect 231766 239536 231822 239572
rect 231950 239536 232006 239592
rect 231122 231512 231178 231568
rect 231030 217096 231086 217152
rect 231306 221312 231362 221368
rect 231214 218728 231270 218784
rect 231398 173440 231454 173496
rect 231674 215872 231730 215928
rect 232042 238720 232098 238776
rect 232318 239672 232374 239728
rect 232226 237360 232282 237416
rect 233192 239808 233248 239864
rect 233422 239828 233478 239864
rect 233422 239808 233424 239828
rect 233424 239808 233476 239828
rect 233476 239808 233478 239828
rect 232870 239536 232926 239592
rect 232778 238584 232834 238640
rect 232870 235728 232926 235784
rect 233054 235320 233110 235376
rect 232410 215056 232466 215112
rect 231950 213560 232006 213616
rect 231582 184184 231638 184240
rect 231306 145696 231362 145752
rect 231214 138896 231270 138952
rect 229742 138760 229798 138816
rect 230478 124752 230534 124808
rect 232778 213288 232834 213344
rect 233422 239672 233478 239728
rect 233330 239536 233386 239592
rect 233238 239400 233294 239456
rect 233238 238720 233294 238776
rect 233238 229880 233294 229936
rect 232686 149776 232742 149832
rect 232594 138624 232650 138680
rect 233698 239672 233754 239728
rect 234296 239808 234352 239864
rect 233606 238584 233662 238640
rect 233790 239420 233846 239456
rect 233790 239400 233792 239420
rect 233792 239400 233844 239420
rect 233844 239400 233846 239420
rect 233974 239400 234030 239456
rect 233882 236000 233938 236056
rect 233790 231376 233846 231432
rect 233606 220224 233662 220280
rect 234158 238584 234214 238640
rect 234066 236000 234122 236056
rect 233974 232872 234030 232928
rect 234434 239672 234490 239728
rect 234848 239808 234904 239864
rect 234526 238176 234582 238232
rect 234434 238040 234490 238096
rect 234894 239400 234950 239456
rect 235078 239672 235134 239728
rect 234986 236272 235042 236328
rect 235170 236680 235226 236736
rect 235538 239672 235594 239728
rect 235446 238720 235502 238776
rect 234802 213152 234858 213208
rect 235354 229744 235410 229800
rect 236090 239672 236146 239728
rect 236320 239808 236376 239864
rect 236504 239808 236560 239864
rect 235906 239400 235962 239456
rect 236182 239400 236238 239456
rect 235538 153040 235594 153096
rect 234710 98776 234766 98832
rect 236550 239672 236606 239728
rect 236458 238720 236514 238776
rect 236458 238176 236514 238232
rect 236366 237496 236422 237552
rect 236182 236988 236184 237008
rect 236184 236988 236236 237008
rect 236236 236988 236238 237008
rect 236182 236952 236238 236988
rect 236182 236136 236238 236192
rect 236734 238720 236790 238776
rect 236642 235184 236698 235240
rect 236366 213696 236422 213752
rect 236182 213016 236238 213072
rect 237010 239400 237066 239456
rect 236918 238176 236974 238232
rect 237332 239842 237388 239898
rect 237654 239672 237710 239728
rect 237194 237768 237250 237824
rect 237286 237088 237342 237144
rect 236826 226752 236882 226808
rect 236734 218864 236790 218920
rect 236918 224712 236974 224768
rect 236826 153856 236882 153912
rect 237470 235728 237526 235784
rect 238528 239896 238584 239898
rect 238528 239844 238530 239896
rect 238530 239844 238582 239896
rect 238582 239844 238584 239896
rect 238528 239842 238584 239844
rect 238298 239400 238354 239456
rect 238896 239808 238952 239864
rect 239540 239808 239596 239864
rect 238666 239400 238722 239456
rect 237930 236952 237986 237008
rect 238114 236680 238170 236736
rect 236734 142976 236790 143032
rect 236642 141480 236698 141536
rect 238390 236952 238446 237008
rect 238942 239436 238944 239456
rect 238944 239436 238996 239456
rect 238996 239436 238998 239456
rect 238942 239400 238998 239436
rect 239310 239436 239312 239456
rect 239312 239436 239364 239456
rect 239364 239436 239366 239456
rect 239310 239400 239366 239436
rect 238850 238176 238906 238232
rect 238758 235592 238814 235648
rect 238666 235456 238722 235512
rect 238298 221448 238354 221504
rect 238114 144200 238170 144256
rect 238942 237496 238998 237552
rect 238850 213832 238906 213888
rect 238574 159432 238630 159488
rect 238482 154264 238538 154320
rect 238298 144064 238354 144120
rect 240138 238720 240194 238776
rect 240368 239808 240424 239864
rect 240828 239808 240884 239864
rect 240322 238584 240378 238640
rect 240690 238720 240746 238776
rect 240874 238176 240930 238232
rect 240874 234232 240930 234288
rect 240690 233824 240746 233880
rect 241196 239842 241252 239898
rect 241702 239808 241758 239864
rect 240690 233144 240746 233200
rect 241150 238584 241206 238640
rect 240690 224712 240746 224768
rect 239770 159296 239826 159352
rect 239678 157120 239734 157176
rect 239494 141616 239550 141672
rect 241242 236680 241298 236736
rect 241426 238584 241482 238640
rect 241426 238040 241482 238096
rect 242116 239808 242172 239864
rect 241242 226344 241298 226400
rect 241150 221584 241206 221640
rect 240874 154128 240930 154184
rect 241886 236680 241942 236736
rect 241794 234368 241850 234424
rect 241978 227024 242034 227080
rect 241978 226344 242034 226400
rect 243128 239842 243184 239898
rect 242898 239400 242954 239456
rect 243266 239672 243322 239728
rect 243082 235864 243138 235920
rect 243266 239400 243322 239456
rect 243266 236816 243322 236872
rect 243082 235320 243138 235376
rect 242806 234096 242862 234152
rect 242254 223216 242310 223272
rect 242806 224984 242862 225040
rect 242254 142024 242310 142080
rect 243450 239672 243506 239728
rect 243358 233552 243414 233608
rect 244738 239828 244794 239864
rect 244738 239808 244740 239828
rect 244740 239808 244792 239828
rect 244792 239808 244794 239828
rect 244462 239400 244518 239456
rect 243910 213424 243966 213480
rect 244738 238176 244794 238232
rect 245382 239808 245438 239864
rect 245290 239400 245346 239456
rect 245382 238584 245438 238640
rect 245658 239672 245714 239728
rect 245934 233144 245990 233200
rect 246348 239842 246404 239898
rect 246394 239708 246396 239728
rect 246396 239708 246448 239728
rect 246448 239708 246450 239728
rect 246394 239672 246450 239708
rect 246992 239808 247048 239864
rect 244278 122168 244334 122224
rect 246394 143248 246450 143304
rect 247544 239808 247600 239864
rect 247314 239400 247370 239456
rect 247866 239400 247922 239456
rect 247682 233824 247738 233880
rect 248142 239692 248198 239728
rect 248142 239672 248144 239692
rect 248144 239672 248196 239692
rect 248196 239672 248198 239692
rect 248648 239808 248704 239864
rect 248326 234232 248382 234288
rect 248878 239692 248934 239728
rect 248878 239672 248880 239692
rect 248880 239672 248932 239692
rect 248932 239672 248934 239692
rect 249752 239808 249808 239864
rect 249890 239708 249892 239728
rect 249892 239708 249944 239728
rect 249944 239708 249946 239728
rect 248786 236408 248842 236464
rect 248786 228520 248842 228576
rect 249522 239400 249578 239456
rect 248970 228520 249026 228576
rect 249338 228384 249394 228440
rect 249890 239672 249946 239708
rect 249890 236680 249946 236736
rect 249430 161064 249486 161120
rect 250304 239842 250360 239898
rect 250074 231920 250130 231976
rect 250534 222128 250590 222184
rect 247682 112376 247738 112432
rect 250994 239672 251050 239728
rect 250718 238584 250774 238640
rect 250810 237904 250866 237960
rect 251454 239672 251510 239728
rect 250994 238720 251050 238776
rect 250902 232736 250958 232792
rect 250902 231920 250958 231976
rect 250534 149912 250590 149968
rect 251822 239808 251878 239864
rect 251914 239672 251970 239728
rect 252098 236408 252154 236464
rect 252604 239842 252660 239898
rect 252742 239672 252798 239728
rect 252558 239400 252614 239456
rect 251178 214784 251234 214840
rect 251270 95920 251326 95976
rect 252558 231376 252614 231432
rect 252466 230016 252522 230072
rect 253018 239400 253074 239456
rect 252926 236544 252982 236600
rect 253294 238040 253350 238096
rect 253386 237224 253442 237280
rect 253110 236680 253166 236736
rect 253018 235184 253074 235240
rect 253662 235728 253718 235784
rect 253846 239400 253902 239456
rect 253110 218048 253166 218104
rect 253110 214512 253166 214568
rect 253294 151272 253350 151328
rect 253938 223080 253994 223136
rect 254720 239808 254776 239864
rect 254490 232328 254546 232384
rect 255134 239672 255190 239728
rect 256100 239842 256156 239898
rect 254858 237768 254914 237824
rect 254398 223080 254454 223136
rect 255134 238584 255190 238640
rect 255410 237904 255466 237960
rect 255226 233144 255282 233200
rect 255042 219136 255098 219192
rect 255042 214920 255098 214976
rect 254766 151408 254822 151464
rect 255686 239128 255742 239184
rect 255594 237768 255650 237824
rect 256054 239708 256056 239728
rect 256056 239708 256108 239728
rect 256108 239708 256110 239728
rect 256054 239672 256110 239708
rect 255962 239400 256018 239456
rect 255870 238720 255926 238776
rect 255778 236680 255834 236736
rect 255686 231376 255742 231432
rect 255778 230424 255834 230480
rect 256146 230424 256202 230480
rect 256054 221992 256110 222048
rect 256238 220224 256294 220280
rect 256238 214648 256294 214704
rect 256054 148688 256110 148744
rect 255318 142860 255374 142896
rect 255318 142840 255320 142860
rect 255320 142840 255372 142860
rect 255372 142840 255374 142860
rect 257158 239672 257214 239728
rect 257250 238720 257306 238776
rect 257250 235728 257306 235784
rect 257250 235320 257306 235376
rect 256974 231512 257030 231568
rect 257618 239400 257674 239456
rect 257526 235048 257582 235104
rect 258124 239808 258180 239864
rect 257526 202136 257582 202192
rect 258538 239692 258594 239728
rect 258538 239672 258540 239692
rect 258540 239672 258592 239692
rect 258592 239672 258594 239692
rect 258078 239400 258134 239456
rect 257434 161200 257490 161256
rect 257618 160928 257674 160984
rect 257526 150048 257582 150104
rect 258262 238312 258318 238368
rect 258354 238040 258410 238096
rect 258814 239400 258870 239456
rect 259090 238720 259146 238776
rect 258998 236680 259054 236736
rect 258814 231104 258870 231160
rect 259458 239708 259460 239728
rect 259460 239708 259512 239728
rect 259512 239708 259514 239728
rect 259458 239672 259514 239708
rect 259182 233280 259238 233336
rect 259274 232328 259330 232384
rect 259734 239400 259790 239456
rect 259642 238448 259698 238504
rect 259734 238332 259790 238368
rect 259734 238312 259736 238332
rect 259736 238312 259788 238332
rect 259788 238312 259790 238332
rect 259734 232192 259790 232248
rect 258814 148824 258870 148880
rect 260516 239808 260572 239864
rect 260792 239808 260848 239864
rect 260470 239400 260526 239456
rect 260378 238720 260434 238776
rect 260378 238584 260434 238640
rect 260654 239400 260710 239456
rect 260654 238584 260710 238640
rect 260562 238040 260618 238096
rect 260470 236408 260526 236464
rect 260746 238312 260802 238368
rect 259918 227296 259974 227352
rect 260102 223352 260158 223408
rect 261436 239808 261492 239864
rect 261390 239672 261446 239728
rect 261022 238584 261078 238640
rect 261022 238312 261078 238368
rect 261298 238584 261354 238640
rect 261390 236136 261446 236192
rect 261666 239672 261722 239728
rect 261942 239400 261998 239456
rect 260930 226208 260986 226264
rect 260286 162016 260342 162072
rect 260194 161336 260250 161392
rect 258538 140664 258594 140720
rect 259550 130328 259606 130384
rect 255318 127608 255374 127664
rect 260930 146104 260986 146160
rect 262632 239808 262688 239864
rect 262402 239400 262458 239456
rect 262126 238176 262182 238232
rect 261666 233008 261722 233064
rect 261850 235048 261906 235104
rect 262310 230832 262366 230888
rect 262586 238720 262642 238776
rect 263184 239808 263240 239864
rect 262494 234504 262550 234560
rect 262862 230152 262918 230208
rect 261850 161880 261906 161936
rect 263598 239692 263654 239728
rect 263598 239672 263600 239692
rect 263600 239672 263652 239692
rect 263652 239672 263654 239692
rect 263598 238176 263654 238232
rect 263506 237632 263562 237688
rect 263322 235184 263378 235240
rect 263046 223488 263102 223544
rect 263782 237632 263838 237688
rect 263782 233824 263838 233880
rect 264104 239808 264160 239864
rect 264150 238720 264206 238776
rect 264058 236544 264114 236600
rect 264656 239808 264712 239864
rect 264886 239672 264942 239728
rect 264702 239420 264758 239456
rect 264702 239400 264704 239420
rect 264704 239400 264756 239420
rect 264756 239400 264758 239420
rect 263690 166232 263746 166288
rect 263598 165008 263654 165064
rect 263046 163512 263102 163568
rect 264334 226208 264390 226264
rect 264886 239400 264942 239456
rect 265392 239808 265448 239864
rect 265162 238720 265218 238776
rect 264978 236680 265034 236736
rect 264610 226752 264666 226808
rect 265530 239708 265532 239728
rect 265532 239708 265584 239728
rect 265584 239708 265586 239728
rect 265530 239672 265586 239708
rect 265254 231784 265310 231840
rect 264978 190984 265034 191040
rect 264334 179968 264390 180024
rect 262954 154400 263010 154456
rect 262862 139304 262918 139360
rect 266036 239844 266038 239864
rect 266038 239844 266090 239864
rect 266090 239844 266092 239864
rect 266036 239808 266092 239844
rect 265714 237088 265770 237144
rect 265806 235320 265862 235376
rect 265714 231784 265770 231840
rect 265622 228928 265678 228984
rect 265622 228792 265678 228848
rect 266312 239672 266368 239728
rect 266174 238720 266230 238776
rect 266358 238176 266414 238232
rect 266082 233824 266138 233880
rect 265990 228792 266046 228848
rect 265714 177248 265770 177304
rect 265622 166368 265678 166424
rect 266818 239672 266874 239728
rect 267002 237768 267058 237824
rect 266910 237088 266966 237144
rect 266634 236680 266690 236736
rect 266910 235456 266966 235512
rect 267002 235048 267058 235104
rect 266818 233960 266874 234016
rect 266450 171672 266506 171728
rect 267186 229880 267242 229936
rect 267738 250416 267794 250472
rect 268014 247560 268070 247616
rect 267922 246336 267978 246392
rect 267738 241576 267794 241632
rect 267738 240216 267794 240272
rect 267370 228656 267426 228712
rect 267278 227432 267334 227488
rect 267462 182824 267518 182880
rect 267278 173304 267334 173360
rect 267094 173168 267150 173224
rect 267002 169088 267058 169144
rect 267922 240080 267978 240136
rect 268290 243616 268346 243672
rect 268106 242256 268162 242312
rect 268198 241576 268254 241632
rect 268014 239944 268070 240000
rect 267922 235456 267978 235512
rect 267830 235184 267886 235240
rect 267646 178608 267702 178664
rect 267554 164872 267610 164928
rect 266174 163376 266230 163432
rect 268474 265512 268530 265568
rect 268566 257352 268622 257408
rect 268474 243616 268530 243672
rect 268474 243480 268530 243536
rect 268750 247832 268806 247888
rect 269118 265512 269174 265568
rect 269118 257388 269120 257408
rect 269120 257388 269172 257408
rect 269172 257388 269174 257408
rect 269118 257352 269174 257388
rect 268842 246472 268898 246528
rect 268842 240624 268898 240680
rect 268658 238720 268714 238776
rect 268382 238312 268438 238368
rect 268106 235048 268162 235104
rect 269302 240488 269358 240544
rect 269670 313792 269726 313848
rect 269670 308760 269726 308816
rect 269486 250688 269542 250744
rect 269578 241440 269634 241496
rect 269486 240216 269542 240272
rect 268934 237224 268990 237280
rect 268014 229880 268070 229936
rect 269118 235728 269174 235784
rect 269578 235592 269634 235648
rect 270406 395256 270462 395312
rect 270130 320320 270186 320376
rect 269854 318144 269910 318200
rect 269762 246608 269818 246664
rect 269946 245112 270002 245168
rect 270130 241712 270186 241768
rect 270222 239264 270278 239320
rect 270130 237224 270186 237280
rect 267922 155624 267978 155680
rect 267830 155488 267886 155544
rect 267922 141752 267978 141808
rect 265622 97280 265678 97336
rect 270314 234368 270370 234424
rect 269762 151544 269818 151600
rect 269762 151136 269818 151192
rect 269118 32408 269174 32464
rect 270590 238584 270646 238640
rect 270590 157256 270646 157312
rect 271418 395664 271474 395720
rect 271418 320864 271474 320920
rect 270682 155216 270738 155272
rect 271050 238448 271106 238504
rect 271234 238040 271290 238096
rect 270958 235320 271014 235376
rect 271694 393896 271750 393952
rect 271786 392536 271842 392592
rect 272522 388456 272578 388512
rect 272246 316648 272302 316704
rect 271786 315968 271842 316024
rect 271786 315016 271842 315072
rect 271694 313656 271750 313712
rect 271694 313384 271750 313440
rect 271602 309576 271658 309632
rect 271786 237360 271842 237416
rect 271694 231376 271750 231432
rect 272798 383016 272854 383072
rect 272522 319776 272578 319832
rect 272798 321408 272854 321464
rect 272798 321000 272854 321056
rect 272982 321408 273038 321464
rect 272798 317056 272854 317112
rect 272614 231104 272670 231160
rect 272982 317192 273038 317248
rect 272982 316648 273038 316704
rect 272982 316240 273038 316296
rect 272798 230424 272854 230480
rect 273994 395800 274050 395856
rect 273718 321000 273774 321056
rect 273166 319232 273222 319288
rect 273166 151680 273222 151736
rect 273166 151000 273222 151056
rect 273442 238176 273498 238232
rect 273994 319640 274050 319696
rect 273810 316104 273866 316160
rect 275926 403008 275982 403064
rect 275558 391312 275614 391368
rect 275466 382880 275522 382936
rect 274546 319640 274602 319696
rect 274546 319096 274602 319152
rect 274178 288360 274234 288416
rect 274546 241304 274602 241360
rect 274546 236408 274602 236464
rect 274362 235864 274418 235920
rect 273626 160792 273682 160848
rect 273534 158888 273590 158944
rect 272246 137944 272302 138000
rect 275282 320184 275338 320240
rect 275558 320728 275614 320784
rect 275466 320592 275522 320648
rect 275558 320456 275614 320512
rect 275466 320184 275522 320240
rect 275374 235864 275430 235920
rect 275190 148960 275246 149016
rect 276018 369416 276074 369472
rect 276018 368600 276074 368656
rect 276386 368600 276442 368656
rect 275834 301280 275890 301336
rect 275650 150184 275706 150240
rect 275190 148280 275246 148336
rect 276202 158752 276258 158808
rect 277122 395528 277178 395584
rect 276938 316376 276994 316432
rect 277674 358828 277730 358864
rect 277674 358808 277676 358828
rect 277676 358808 277728 358828
rect 277728 358808 277730 358828
rect 277490 240216 277546 240272
rect 277030 155080 277086 155136
rect 278042 321408 278098 321464
rect 278042 320592 278098 320648
rect 278042 315152 278098 315208
rect 277766 314336 277822 314392
rect 277858 240216 277914 240272
rect 277950 236272 278006 236328
rect 278318 321000 278374 321056
rect 278042 222808 278098 222864
rect 277490 160656 277546 160712
rect 276110 109656 276166 109712
rect 279146 384240 279202 384296
rect 278870 228248 278926 228304
rect 278962 159024 279018 159080
rect 279606 320048 279662 320104
rect 279606 317872 279662 317928
rect 280710 451424 280766 451480
rect 280066 401784 280122 401840
rect 281078 449112 281134 449168
rect 280710 371628 280712 371648
rect 280712 371628 280764 371648
rect 280764 371628 280766 371648
rect 280710 371592 280766 371628
rect 280434 369688 280490 369744
rect 280434 369280 280490 369336
rect 279790 236952 279846 237008
rect 280158 221856 280214 221912
rect 280710 356768 280766 356824
rect 280710 345752 280766 345808
rect 280710 319776 280766 319832
rect 280710 317872 280766 317928
rect 281170 372136 281226 372192
rect 281262 356768 281318 356824
rect 281078 345752 281134 345808
rect 281446 372000 281502 372056
rect 281630 320456 281686 320512
rect 281722 320184 281778 320240
rect 281998 319776 282054 319832
rect 281814 319504 281870 319560
rect 281722 319368 281778 319424
rect 281906 319368 281962 319424
rect 281998 318960 282054 319016
rect 286322 448976 286378 449032
rect 284482 444896 284538 444952
rect 282274 371864 282330 371920
rect 285034 401920 285090 401976
rect 285126 392672 285182 392728
rect 284574 372816 284630 372872
rect 284482 369960 284538 370016
rect 286690 372952 286746 373008
rect 286046 372680 286102 372736
rect 284942 370096 284998 370152
rect 284850 369960 284906 370016
rect 286046 370096 286102 370152
rect 285080 369552 285136 369608
rect 290002 372136 290058 372192
rect 289634 371456 289690 371512
rect 289358 370640 289414 370696
rect 288024 369688 288080 369744
rect 287288 369552 287344 369608
rect 291934 439456 291990 439512
rect 293314 400832 293370 400888
rect 290646 372272 290702 372328
rect 291842 372272 291898 372328
rect 290646 371320 290702 371376
rect 290094 369416 290150 369472
rect 293314 372000 293370 372056
rect 295338 398112 295394 398168
rect 298742 399744 298798 399800
rect 297362 371864 297418 371920
rect 300122 451560 300178 451616
rect 298926 400968 298982 401024
rect 300214 449928 300270 449984
rect 300306 400016 300362 400072
rect 300122 370096 300178 370152
rect 300398 381792 300454 381848
rect 301594 446392 301650 446448
rect 302974 398248 303030 398304
rect 302974 385736 303030 385792
rect 302974 370776 303030 370832
rect 302744 369824 302800 369880
rect 304998 395936 305054 395992
rect 305090 395120 305146 395176
rect 308402 452784 308458 452840
rect 307942 390632 307998 390688
rect 312542 448840 312598 448896
rect 309782 447752 309838 447808
rect 309966 391856 310022 391912
rect 309782 375400 309838 375456
rect 310242 371728 310298 371784
rect 310702 371592 310758 371648
rect 310610 370232 310666 370288
rect 302146 369416 302202 369472
rect 303342 369416 303398 369472
rect 310702 369824 310758 369880
rect 311576 369824 311632 369880
rect 312818 399472 312874 399528
rect 312726 387640 312782 387696
rect 312082 369688 312138 369744
rect 311806 369552 311862 369608
rect 314014 450064 314070 450120
rect 313922 401240 313978 401296
rect 313554 370368 313610 370424
rect 315302 399608 315358 399664
rect 314382 369552 314438 369608
rect 315854 369824 315910 369880
rect 319718 401104 319774 401160
rect 319902 369552 319958 369608
rect 323766 399880 323822 399936
rect 324226 389952 324282 390008
rect 324318 385736 324374 385792
rect 321374 369552 321430 369608
rect 324870 370776 324926 370832
rect 311438 369416 311494 369472
rect 313186 369416 313242 369472
rect 314290 369416 314346 369472
rect 318706 369416 318762 369472
rect 319810 369416 319866 369472
rect 321282 369416 321338 369472
rect 285816 369280 285872 369336
rect 287288 369280 287344 369336
rect 309000 369280 309056 369336
rect 310104 369280 310160 369336
rect 282274 360848 282330 360904
rect 282182 353912 282238 353968
rect 327446 333240 327502 333296
rect 327538 330384 327594 330440
rect 327446 321544 327502 321600
rect 282274 321272 282330 321328
rect 282274 320728 282330 320784
rect 283240 320728 283296 320784
rect 284252 320728 284308 320784
rect 287472 320728 287528 320784
rect 288208 320728 288264 320784
rect 290600 320728 290656 320784
rect 291152 320728 291208 320784
rect 291888 320728 291944 320784
rect 292624 320728 292680 320784
rect 296488 320728 296544 320784
rect 297316 320728 297372 320784
rect 298144 320728 298200 320784
rect 299064 320728 299120 320784
rect 303388 320728 303444 320784
rect 306700 320728 306756 320784
rect 308816 320728 308872 320784
rect 323536 320728 323592 320784
rect 324088 320728 324144 320784
rect 324364 320728 324420 320784
rect 325192 320728 325248 320784
rect 325744 320728 325800 320784
rect 327032 320728 327088 320784
rect 283332 320592 283388 320648
rect 283608 320592 283664 320648
rect 286184 320592 286240 320648
rect 313048 320592 313104 320648
rect 315808 320592 315864 320648
rect 317096 320592 317152 320648
rect 317648 320592 317704 320648
rect 318016 320592 318072 320648
rect 318200 320592 318256 320648
rect 318936 320592 318992 320648
rect 319212 320592 319268 320648
rect 282274 320456 282330 320512
rect 282872 320456 282928 320512
rect 283976 320456 284032 320512
rect 286552 320456 286608 320512
rect 288668 320456 288724 320512
rect 292348 320456 292404 320512
rect 293728 320456 293784 320512
rect 294004 320456 294060 320512
rect 294832 320456 294888 320512
rect 297868 320456 297924 320512
rect 298604 320456 298660 320512
rect 305596 320456 305652 320512
rect 308356 320456 308412 320512
rect 310380 320456 310436 320512
rect 322064 320456 322120 320512
rect 322248 320456 322304 320512
rect 323352 320456 323408 320512
rect 323812 320456 323868 320512
rect 324640 320456 324696 320512
rect 326112 320456 326168 320512
rect 284344 320320 284400 320376
rect 285448 320320 285504 320376
rect 285724 320320 285780 320376
rect 287748 320320 287804 320376
rect 289496 320320 289552 320376
rect 290048 320320 290104 320376
rect 291704 320320 291760 320376
rect 307896 320320 307952 320376
rect 309552 320320 309608 320376
rect 310104 320320 310160 320376
rect 310288 320320 310344 320376
rect 310656 320320 310712 320376
rect 311392 320320 311448 320376
rect 316452 320320 316508 320376
rect 320132 320320 320188 320376
rect 320316 320320 320372 320376
rect 320776 320320 320832 320376
rect 321604 320320 321660 320376
rect 323260 320320 323316 320376
rect 324272 320320 324328 320376
rect 325468 320320 325524 320376
rect 326388 320320 326444 320376
rect 327400 320320 327456 320376
rect 282504 320184 282560 320240
rect 292808 320184 292864 320240
rect 293176 320184 293232 320240
rect 294188 320184 294244 320240
rect 294556 320184 294612 320240
rect 295936 320184 295992 320240
rect 297040 320184 297096 320240
rect 297408 320184 297464 320240
rect 298420 320184 298476 320240
rect 302008 320184 302064 320240
rect 307988 320184 308044 320240
rect 312036 320184 312092 320240
rect 312680 320184 312736 320240
rect 313600 320184 313656 320240
rect 314152 320184 314208 320240
rect 316636 320184 316692 320240
rect 317740 320184 317796 320240
rect 282550 319504 282606 319560
rect 283148 320048 283204 320104
rect 282090 306856 282146 306912
rect 282090 235048 282146 235104
rect 281078 231648 281134 231704
rect 280802 218592 280858 218648
rect 282826 318688 282882 318744
rect 283010 319096 283066 319152
rect 283102 318824 283158 318880
rect 282458 238992 282514 239048
rect 282458 233960 282514 234016
rect 283286 319368 283342 319424
rect 283286 317600 283342 317656
rect 283792 320048 283848 320104
rect 283746 319368 283802 319424
rect 283654 317464 283710 317520
rect 284298 319776 284354 319832
rect 284022 317736 284078 317792
rect 284712 320048 284768 320104
rect 284390 317736 284446 317792
rect 284206 317192 284262 317248
rect 283470 296112 283526 296168
rect 282918 238856 282974 238912
rect 282918 236000 282974 236056
rect 280158 108296 280214 108352
rect 283470 236816 283526 236872
rect 283470 236000 283526 236056
rect 284114 241168 284170 241224
rect 283930 225800 283986 225856
rect 284574 318688 284630 318744
rect 284390 241984 284446 242040
rect 285172 320048 285228 320104
rect 284666 295024 284722 295080
rect 284666 293936 284722 293992
rect 285586 319640 285642 319696
rect 285402 318552 285458 318608
rect 285402 317736 285458 317792
rect 286276 320048 286332 320104
rect 285862 319232 285918 319288
rect 286046 310256 286102 310312
rect 285310 302912 285366 302968
rect 285218 301960 285274 302016
rect 285126 293936 285182 293992
rect 284758 240896 284814 240952
rect 285126 239536 285182 239592
rect 284758 237360 284814 237416
rect 285126 233824 285182 233880
rect 284390 94424 284446 94480
rect 287104 320048 287160 320104
rect 287334 319640 287390 319696
rect 285310 227024 285366 227080
rect 285218 222944 285274 223000
rect 286506 309712 286562 309768
rect 286598 295160 286654 295216
rect 286874 295160 286930 295216
rect 287242 298968 287298 299024
rect 288300 320048 288356 320104
rect 287794 319640 287850 319696
rect 287702 319232 287758 319288
rect 287978 319640 288034 319696
rect 288254 319776 288310 319832
rect 288576 320048 288632 320104
rect 288944 320048 289000 320104
rect 287794 295976 287850 296032
rect 286690 231104 286746 231160
rect 287058 26832 287114 26888
rect 288162 315696 288218 315752
rect 288162 314880 288218 314936
rect 288622 319232 288678 319288
rect 288714 319096 288770 319152
rect 288438 310392 288494 310448
rect 287978 296248 288034 296304
rect 288254 298968 288310 299024
rect 289312 320048 289368 320104
rect 289680 320048 289736 320104
rect 289864 320048 289920 320104
rect 289174 317464 289230 317520
rect 289450 319640 289506 319696
rect 289358 317328 289414 317384
rect 288898 294888 288954 294944
rect 289174 310800 289230 310856
rect 289174 239400 289230 239456
rect 289726 319776 289782 319832
rect 289634 318280 289690 318336
rect 290416 320048 290472 320104
rect 290094 318280 290150 318336
rect 290278 319640 290334 319696
rect 290462 319776 290518 319832
rect 290094 317464 290150 317520
rect 290002 311480 290058 311536
rect 290876 320048 290932 320104
rect 291428 320048 291484 320104
rect 291106 319640 291162 319696
rect 290738 319096 290794 319152
rect 290830 318824 290886 318880
rect 290738 316784 290794 316840
rect 289634 294480 289690 294536
rect 291014 318824 291070 318880
rect 291198 315696 291254 315752
rect 291106 310392 291162 310448
rect 290646 247968 290702 248024
rect 291382 301824 291438 301880
rect 291842 319232 291898 319288
rect 291658 294344 291714 294400
rect 292164 320048 292220 320104
rect 292118 319640 292174 319696
rect 291842 317736 291898 317792
rect 292026 318144 292082 318200
rect 292486 319660 292542 319696
rect 292486 319640 292488 319660
rect 292488 319640 292540 319660
rect 292540 319640 292542 319660
rect 292670 319504 292726 319560
rect 293268 319878 293324 319934
rect 290554 220768 290610 220824
rect 292118 301824 292174 301880
rect 292394 300192 292450 300248
rect 292118 220496 292174 220552
rect 293038 319640 293094 319696
rect 293452 320048 293508 320104
rect 292670 314472 292726 314528
rect 294280 320048 294336 320104
rect 293590 319504 293646 319560
rect 292302 220632 292358 220688
rect 293682 317464 293738 317520
rect 293866 313656 293922 313712
rect 294464 320048 294520 320104
rect 294142 319776 294198 319832
rect 294142 319232 294198 319288
rect 294234 318416 294290 318472
rect 294740 320048 294796 320104
rect 294418 319776 294474 319832
rect 294510 319096 294566 319152
rect 294418 315968 294474 316024
rect 293958 298832 294014 298888
rect 294694 315696 294750 315752
rect 294694 315424 294750 315480
rect 294602 236544 294658 236600
rect 293314 218592 293370 218648
rect 295476 319878 295532 319934
rect 295154 299376 295210 299432
rect 294786 230016 294842 230072
rect 296120 320048 296176 320104
rect 296304 320048 296360 320104
rect 295614 319640 295670 319696
rect 296166 319776 296222 319832
rect 295338 304408 295394 304464
rect 295338 301416 295394 301472
rect 295338 235864 295394 235920
rect 296166 319640 296222 319696
rect 296258 313928 296314 313984
rect 295062 227160 295118 227216
rect 297224 320048 297280 320104
rect 296350 304544 296406 304600
rect 297086 319232 297142 319288
rect 297086 318552 297142 318608
rect 297592 320048 297648 320104
rect 298052 320048 298108 320104
rect 297270 319640 297326 319696
rect 297178 318280 297234 318336
rect 297178 317600 297234 317656
rect 297086 317464 297142 317520
rect 296902 316648 296958 316704
rect 297730 317464 297786 317520
rect 296626 235864 296682 235920
rect 298006 319776 298062 319832
rect 297822 304136 297878 304192
rect 298190 319640 298246 319696
rect 298190 317872 298246 317928
rect 298374 319232 298430 319288
rect 298098 314200 298154 314256
rect 298098 308488 298154 308544
rect 298880 319878 298936 319934
rect 299248 320048 299304 320104
rect 298742 319640 298798 319696
rect 297914 293120 297970 293176
rect 298190 236680 298246 236736
rect 298834 308624 298890 308680
rect 299294 319640 299350 319696
rect 299294 318008 299350 318064
rect 299018 302096 299074 302152
rect 299616 320048 299672 320104
rect 299570 319640 299626 319696
rect 300030 317464 300086 317520
rect 299846 314472 299902 314528
rect 299846 312568 299902 312624
rect 300720 320048 300776 320104
rect 300904 320048 300960 320104
rect 300306 317872 300362 317928
rect 299294 293392 299350 293448
rect 299018 236680 299074 236736
rect 298190 150320 298246 150376
rect 299386 150320 299442 150376
rect 299386 149640 299442 149696
rect 300582 302232 300638 302288
rect 301272 319878 301328 319934
rect 300858 313540 300914 313576
rect 300858 313520 300860 313540
rect 300860 313520 300912 313540
rect 300912 313520 300914 313540
rect 300674 301688 300730 301744
rect 300582 293256 300638 293312
rect 300306 230288 300362 230344
rect 300122 224848 300178 224904
rect 301732 320048 301788 320104
rect 301318 319640 301374 319696
rect 301226 314336 301282 314392
rect 302192 320048 302248 320104
rect 301502 315832 301558 315888
rect 301410 315560 301466 315616
rect 301226 313384 301282 313440
rect 301502 315152 301558 315208
rect 301870 319640 301926 319696
rect 301778 315696 301834 315752
rect 301686 314200 301742 314256
rect 301134 303456 301190 303512
rect 301134 302948 301136 302968
rect 301136 302948 301188 302968
rect 301188 302948 301190 302968
rect 301134 302912 301190 302948
rect 301962 317464 302018 317520
rect 302560 319878 302616 319934
rect 302836 320048 302892 320104
rect 302146 319096 302202 319152
rect 302698 319640 302754 319696
rect 302330 318144 302386 318200
rect 302698 318688 302754 318744
rect 302238 300192 302294 300248
rect 302698 307128 302754 307184
rect 303066 317872 303122 317928
rect 303066 316648 303122 316704
rect 303342 319660 303398 319696
rect 303342 319640 303344 319660
rect 303344 319640 303396 319660
rect 303396 319640 303398 319660
rect 303250 317464 303306 317520
rect 303250 316376 303306 316432
rect 303940 320048 303996 320104
rect 304216 320048 304272 320104
rect 304584 320048 304640 320104
rect 303434 303456 303490 303512
rect 303526 303184 303582 303240
rect 303526 297628 303582 297664
rect 303526 297608 303528 297628
rect 303528 297608 303580 297628
rect 303580 297608 303582 297628
rect 303158 239128 303214 239184
rect 304078 319504 304134 319560
rect 304262 319640 304318 319696
rect 304538 319640 304594 319696
rect 304262 317872 304318 317928
rect 304538 318008 304594 318064
rect 304446 317464 304502 317520
rect 304170 297880 304226 297936
rect 304170 290808 304226 290864
rect 305136 319878 305192 319934
rect 304998 319504 305054 319560
rect 304906 316240 304962 316296
rect 304998 309848 305054 309904
rect 305182 319232 305238 319288
rect 305872 320048 305928 320104
rect 306332 320048 306388 320104
rect 305458 289720 305514 289776
rect 306010 305632 306066 305688
rect 305826 301416 305882 301472
rect 301962 6024 302018 6080
rect 305826 221720 305882 221776
rect 306746 319776 306802 319832
rect 306976 320048 307032 320104
rect 306746 317464 306802 317520
rect 307528 320048 307584 320104
rect 307482 318280 307538 318336
rect 307206 317872 307262 317928
rect 307574 314608 307630 314664
rect 307758 313148 307760 313168
rect 307760 313148 307812 313168
rect 307812 313148 307814 313168
rect 307758 313112 307814 313148
rect 307758 301960 307814 302016
rect 307574 290400 307630 290456
rect 307114 228384 307170 228440
rect 308632 320048 308688 320104
rect 309736 320048 309792 320104
rect 307850 291760 307906 291816
rect 308954 307264 309010 307320
rect 309138 312160 309194 312216
rect 309598 319776 309654 319832
rect 309506 318552 309562 318608
rect 309920 320048 309976 320104
rect 309874 319776 309930 319832
rect 310150 319812 310152 319832
rect 310152 319812 310204 319832
rect 310204 319812 310206 319832
rect 310150 319776 310206 319812
rect 309782 308352 309838 308408
rect 310150 319504 310206 319560
rect 310242 319232 310298 319288
rect 310150 291760 310206 291816
rect 310058 289176 310114 289232
rect 310932 320048 310988 320104
rect 310702 319504 310758 319560
rect 311668 320048 311724 320104
rect 310702 304408 310758 304464
rect 310886 304272 310942 304328
rect 310702 303728 310758 303784
rect 310886 303592 310942 303648
rect 310150 234232 310206 234288
rect 311944 320048 312000 320104
rect 311898 319660 311954 319696
rect 311898 319640 311900 319660
rect 311900 319640 311952 319660
rect 311952 319640 311954 319660
rect 311898 312840 311954 312896
rect 311254 303728 311310 303784
rect 311438 303592 311494 303648
rect 311530 299240 311586 299296
rect 312772 320048 312828 320104
rect 312358 315424 312414 315480
rect 312542 317464 312598 317520
rect 312818 319776 312874 319832
rect 313094 319776 313150 319832
rect 312082 304544 312138 304600
rect 313416 320048 313472 320104
rect 313692 319776 313748 319832
rect 313278 319640 313334 319696
rect 313370 317872 313426 317928
rect 313278 317736 313334 317792
rect 313186 312568 313242 312624
rect 313646 319504 313702 319560
rect 313646 318960 313702 319016
rect 314106 319640 314162 319696
rect 313830 317872 313886 317928
rect 314014 317872 314070 317928
rect 313278 303320 313334 303376
rect 314428 320048 314484 320104
rect 314658 319776 314714 319832
rect 314888 320048 314944 320104
rect 314198 319232 314254 319288
rect 314106 315968 314162 316024
rect 314106 314472 314162 314528
rect 314382 304136 314438 304192
rect 315256 320048 315312 320104
rect 315578 319660 315634 319696
rect 315578 319640 315580 319660
rect 315580 319640 315632 319660
rect 315632 319640 315634 319660
rect 314842 303592 314898 303648
rect 315578 317872 315634 317928
rect 315762 317464 315818 317520
rect 316176 320048 316232 320104
rect 316038 319640 316094 319696
rect 315394 258712 315450 258768
rect 316130 317600 316186 317656
rect 316912 320048 316968 320104
rect 316866 318552 316922 318608
rect 316866 318416 316922 318472
rect 317050 319640 317106 319696
rect 317142 318688 317198 318744
rect 317142 318552 317198 318608
rect 317050 317056 317106 317112
rect 317234 317464 317290 317520
rect 318292 320048 318348 320104
rect 317510 319096 317566 319152
rect 317418 318960 317474 319016
rect 316590 311752 316646 311808
rect 316682 299240 316738 299296
rect 316866 267008 316922 267064
rect 316774 264152 316830 264208
rect 316682 251776 316738 251832
rect 315486 222128 315542 222184
rect 317234 311752 317290 311808
rect 317878 319676 317880 319696
rect 317880 319676 317932 319696
rect 317932 319676 317934 319696
rect 317878 319640 317934 319676
rect 317878 319504 317934 319560
rect 318154 319504 318210 319560
rect 318568 320048 318624 320104
rect 318246 319368 318302 319424
rect 318338 319096 318394 319152
rect 318430 317464 318486 317520
rect 319120 320048 319176 320104
rect 317878 311208 317934 311264
rect 317694 306312 317750 306368
rect 317694 304952 317750 305008
rect 317418 299240 317474 299296
rect 318062 299240 318118 299296
rect 318982 319368 319038 319424
rect 318890 318688 318946 318744
rect 318890 318008 318946 318064
rect 318522 311208 318578 311264
rect 318338 304952 318394 305008
rect 318246 300736 318302 300792
rect 318154 262792 318210 262848
rect 318062 244840 318118 244896
rect 318246 250416 318302 250472
rect 319258 319776 319314 319832
rect 319258 319096 319314 319152
rect 318982 309032 319038 309088
rect 319672 320048 319728 320104
rect 319442 315152 319498 315208
rect 319534 313792 319590 313848
rect 319810 318824 319866 318880
rect 319902 318552 319958 318608
rect 320178 319640 320234 319696
rect 320270 317464 320326 317520
rect 320684 320048 320740 320104
rect 320454 319368 320510 319424
rect 320178 316104 320234 316160
rect 321328 320048 321384 320104
rect 321236 319878 321292 319934
rect 320822 319368 320878 319424
rect 321006 318960 321062 319016
rect 320914 317872 320970 317928
rect 321006 317736 321062 317792
rect 320822 315696 320878 315752
rect 319994 315152 320050 315208
rect 319718 305904 319774 305960
rect 319534 250688 319590 250744
rect 319902 309032 319958 309088
rect 319902 308488 319958 308544
rect 319626 242120 319682 242176
rect 321006 315696 321062 315752
rect 320914 312976 320970 313032
rect 320730 304408 320786 304464
rect 321374 319640 321430 319696
rect 321742 319660 321798 319696
rect 321742 319640 321744 319660
rect 321744 319640 321796 319660
rect 321796 319640 321798 319660
rect 321558 318280 321614 318336
rect 321466 312976 321522 313032
rect 321098 307672 321154 307728
rect 321282 304292 321338 304328
rect 321282 304272 321284 304292
rect 321284 304272 321336 304292
rect 321336 304272 321338 304292
rect 321098 257216 321154 257272
rect 321742 319504 321798 319560
rect 321834 319368 321890 319424
rect 322524 320048 322580 320104
rect 322110 319776 322166 319832
rect 322294 319640 322350 319696
rect 322110 319096 322166 319152
rect 322110 318960 322166 319016
rect 322202 317464 322258 317520
rect 322478 319504 322534 319560
rect 322386 316784 322442 316840
rect 322662 319640 322718 319696
rect 322018 311072 322074 311128
rect 322202 311072 322258 311128
rect 322110 310936 322166 310992
rect 321926 310120 321982 310176
rect 321834 309032 321890 309088
rect 321742 306176 321798 306232
rect 321742 304952 321798 305008
rect 321650 301416 321706 301472
rect 321006 247560 321062 247616
rect 322294 309032 322350 309088
rect 322202 243480 322258 243536
rect 322938 319096 322994 319152
rect 323214 319640 323270 319696
rect 323214 317872 323270 317928
rect 322570 310120 322626 310176
rect 322938 309984 322994 310040
rect 322938 309712 322994 309768
rect 323214 312840 323270 312896
rect 323490 318960 323546 319016
rect 323490 318144 323546 318200
rect 323398 314608 323454 314664
rect 323306 310256 323362 310312
rect 323030 309032 323086 309088
rect 322846 304952 322902 305008
rect 322754 290536 322810 290592
rect 322570 253136 322626 253192
rect 322478 246336 322534 246392
rect 323582 314336 323638 314392
rect 323858 313112 323914 313168
rect 323490 300600 323546 300656
rect 324042 319640 324098 319696
rect 324042 318416 324098 318472
rect 324042 318008 324098 318064
rect 324226 318960 324282 319016
rect 324502 318688 324558 318744
rect 324134 312840 324190 312896
rect 324042 309032 324098 309088
rect 322938 273808 322994 273864
rect 323766 287680 323822 287736
rect 324916 320048 324972 320104
rect 324962 319640 325018 319696
rect 324870 317328 324926 317384
rect 324686 313656 324742 313712
rect 325054 318960 325110 319016
rect 325238 318960 325294 319016
rect 325422 318960 325478 319016
rect 325238 317192 325294 317248
rect 325146 314472 325202 314528
rect 324410 311208 324466 311264
rect 324962 311208 325018 311264
rect 324226 310256 324282 310312
rect 323582 247696 323638 247752
rect 311898 106936 311954 106992
rect 315302 100136 315358 100192
rect 318062 69536 318118 69592
rect 322386 229744 322442 229800
rect 325146 301960 325202 302016
rect 325330 314472 325386 314528
rect 325330 313928 325386 313984
rect 325422 301960 325478 302016
rect 325146 264288 325202 264344
rect 325054 244976 325110 245032
rect 326848 320048 326904 320104
rect 327216 320048 327272 320104
rect 326342 319524 326398 319560
rect 326342 319504 326344 319524
rect 326344 319504 326396 319524
rect 326396 319504 326398 319524
rect 326158 315560 326214 315616
rect 326066 312704 326122 312760
rect 327630 321544 327686 321600
rect 327630 320728 327686 320784
rect 327630 320492 327632 320512
rect 327632 320492 327684 320512
rect 327684 320492 327686 320512
rect 327630 320456 327686 320492
rect 327630 320320 327686 320376
rect 326802 319504 326858 319560
rect 326710 318960 326766 319016
rect 326618 317600 326674 317656
rect 326618 316240 326674 316296
rect 326526 314200 326582 314256
rect 325974 307536 326030 307592
rect 325882 306040 325938 306096
rect 325790 302776 325846 302832
rect 326434 307536 326490 307592
rect 326342 249056 326398 249112
rect 326802 317056 326858 317112
rect 327078 319504 327134 319560
rect 326986 317464 327042 317520
rect 326894 316648 326950 316704
rect 326802 316240 326858 316296
rect 327446 318960 327502 319016
rect 326986 312704 327042 312760
rect 326710 309712 326766 309768
rect 326802 306040 326858 306096
rect 326894 303456 326950 303512
rect 326894 302776 326950 302832
rect 326618 271088 326674 271144
rect 326526 260072 326582 260128
rect 326434 246200 326490 246256
rect 327262 317736 327318 317792
rect 327170 253272 327226 253328
rect 326342 228792 326398 228848
rect 327354 315288 327410 315344
rect 327354 313656 327410 313712
rect 327814 357992 327870 358048
rect 328366 366424 328422 366480
rect 327906 341536 327962 341592
rect 327998 327664 328054 327720
rect 327906 321136 327962 321192
rect 327814 321000 327870 321056
rect 327814 320456 327870 320512
rect 327906 320320 327962 320376
rect 328366 321408 328422 321464
rect 328366 321136 328422 321192
rect 327998 317736 328054 317792
rect 328918 320048 328974 320104
rect 328458 316648 328514 316704
rect 327630 247832 327686 247888
rect 328458 309576 328514 309632
rect 327538 229880 327594 229936
rect 322938 12960 322994 13016
rect 328918 317872 328974 317928
rect 330482 398384 330538 398440
rect 329194 319912 329250 319968
rect 329194 319368 329250 319424
rect 329194 318280 329250 318336
rect 329378 386008 329434 386064
rect 330298 323720 330354 323776
rect 329838 322904 329894 322960
rect 330298 322904 330354 322960
rect 329378 318008 329434 318064
rect 329194 316240 329250 316296
rect 329378 316104 329434 316160
rect 329746 318688 329802 318744
rect 329654 318552 329710 318608
rect 329746 317600 329802 317656
rect 329010 311344 329066 311400
rect 329010 311072 329066 311128
rect 330206 321272 330262 321328
rect 329930 318008 329986 318064
rect 330390 310392 330446 310448
rect 330390 310120 330446 310176
rect 331954 397296 332010 397352
rect 330758 397160 330814 397216
rect 330574 396480 330630 396536
rect 330942 321272 330998 321328
rect 331218 327120 331274 327176
rect 330850 311616 330906 311672
rect 330758 309984 330814 310040
rect 330758 309712 330814 309768
rect 331678 320048 331734 320104
rect 331310 318552 331366 318608
rect 331494 318144 331550 318200
rect 332322 318144 332378 318200
rect 332414 314608 332470 314664
rect 332690 317600 332746 317656
rect 332046 236544 332102 236600
rect 331494 235184 331550 235240
rect 331310 233960 331366 234016
rect 331218 231784 331274 231840
rect 329838 228928 329894 228984
rect 332874 319232 332930 319288
rect 332690 235320 332746 235376
rect 333610 315968 333666 316024
rect 334990 450200 335046 450256
rect 333978 371864 334034 371920
rect 334622 368736 334678 368792
rect 333978 319912 334034 319968
rect 333886 319640 333942 319696
rect 333886 319232 333942 319288
rect 333702 312704 333758 312760
rect 333518 237224 333574 237280
rect 332874 233144 332930 233200
rect 334070 315424 334126 315480
rect 333978 233008 334034 233064
rect 334530 320592 334586 320648
rect 334530 320320 334586 320376
rect 334254 312604 334256 312624
rect 334256 312604 334308 312624
rect 334308 312604 334310 312624
rect 334254 312568 334310 312604
rect 334254 237904 334310 237960
rect 334898 395120 334954 395176
rect 335910 400424 335966 400480
rect 335818 395800 335874 395856
rect 334990 368328 335046 368384
rect 334990 317464 335046 317520
rect 335174 315424 335230 315480
rect 337474 454144 337530 454200
rect 337658 454008 337714 454064
rect 336554 400288 336610 400344
rect 336738 321544 336794 321600
rect 335542 233824 335598 233880
rect 336830 320320 336886 320376
rect 336922 320184 336978 320240
rect 337934 325080 337990 325136
rect 338210 321000 338266 321056
rect 338118 320592 338174 320648
rect 337934 320320 337990 320376
rect 338118 320184 338174 320240
rect 336830 227568 336886 227624
rect 336738 227432 336794 227488
rect 338210 319096 338266 319152
rect 338210 316512 338266 316568
rect 339222 397840 339278 397896
rect 339406 449656 339462 449712
rect 340234 448568 340290 448624
rect 339406 368600 339462 368656
rect 339498 321816 339554 321872
rect 339958 321816 340014 321872
rect 339314 320184 339370 320240
rect 339222 315288 339278 315344
rect 340050 321136 340106 321192
rect 339590 316648 339646 316704
rect 340510 334600 340566 334656
rect 340510 316648 340566 316704
rect 340878 451696 340934 451752
rect 340970 438232 341026 438288
rect 340970 436756 341026 436792
rect 340970 436736 340972 436756
rect 340972 436736 341024 436756
rect 341024 436736 341026 436756
rect 340970 428460 341026 428496
rect 340970 428440 340972 428460
rect 340972 428440 341024 428460
rect 341024 428440 341026 428460
rect 347778 452648 347834 452704
rect 345570 451832 345626 451888
rect 340970 405728 341026 405784
rect 340878 399200 340934 399256
rect 340878 398792 340934 398848
rect 341062 398792 341118 398848
rect 345202 451424 345258 451480
rect 341890 438232 341946 438288
rect 341798 436736 341854 436792
rect 341706 428440 341762 428496
rect 341614 405728 341670 405784
rect 342074 403008 342130 403064
rect 341982 402056 342038 402112
rect 341706 400696 341762 400752
rect 341614 400016 341670 400072
rect 341062 398248 341118 398304
rect 341430 398248 341486 398304
rect 340878 324944 340934 325000
rect 341522 368600 341578 368656
rect 340878 223488 340934 223544
rect 330390 6840 330446 6896
rect 333886 6704 333942 6760
rect 337474 6568 337530 6624
rect 342074 399336 342130 399392
rect 345938 451560 345994 451616
rect 352930 451288 352986 451344
rect 347272 449656 347328 449712
rect 346536 449520 346592 449576
rect 344466 449384 344522 449440
rect 345202 449384 345258 449440
rect 349342 449384 349398 449440
rect 353390 449384 353446 449440
rect 358082 449384 358138 449440
rect 358634 451560 358690 451616
rect 359554 451288 359610 451344
rect 360152 449928 360208 449984
rect 361670 452512 361726 452568
rect 361670 452104 361726 452160
rect 362222 452512 362278 452568
rect 368018 452784 368074 452840
rect 368570 452512 368626 452568
rect 368570 451424 368626 451480
rect 369490 452512 369546 452568
rect 371330 454144 371386 454200
rect 370088 450200 370144 450256
rect 371422 451696 371478 451752
rect 372802 454008 372858 454064
rect 372618 452512 372674 452568
rect 373400 450064 373456 450120
rect 374090 452512 374146 452568
rect 373998 451424 374054 451480
rect 378690 451288 378746 451344
rect 580170 697176 580226 697232
rect 580262 683848 580318 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 579986 630808 580042 630864
rect 580170 617480 580226 617536
rect 580170 590960 580226 591016
rect 580170 577632 580226 577688
rect 580170 564304 580226 564360
rect 579894 537784 579950 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580354 511264 580410 511320
rect 580170 484608 580226 484664
rect 580078 471416 580134 471472
rect 580170 458088 580226 458144
rect 371928 449520 371984 449576
rect 370594 449420 370596 449440
rect 370596 449420 370648 449440
rect 370648 449420 370650 449440
rect 370594 449384 370650 449420
rect 372066 449384 372122 449440
rect 372802 449384 372858 449440
rect 375010 449384 375066 449440
rect 383106 449384 383162 449440
rect 383842 449384 383898 449440
rect 384302 449384 384358 449440
rect 385682 449384 385738 449440
rect 343960 449248 344016 449304
rect 346904 449248 346960 449304
rect 368984 449248 369040 449304
rect 374872 449248 374928 449304
rect 385544 449248 385600 449304
rect 342442 439456 342498 439512
rect 580170 431568 580226 431624
rect 580262 418240 580318 418296
rect 580170 404912 580226 404968
rect 580722 400832 580778 400888
rect 342258 395392 342314 395448
rect 342258 389136 342314 389192
rect 342810 398112 342866 398168
rect 342350 325216 342406 325272
rect 343362 396752 343418 396808
rect 344006 399200 344062 399256
rect 343638 394304 343694 394360
rect 343270 383424 343326 383480
rect 343730 391176 343786 391232
rect 343454 387368 343510 387424
rect 344190 395800 344246 395856
rect 344190 386960 344246 387016
rect 344098 312840 344154 312896
rect 344466 398928 344522 398984
rect 344650 398928 344706 398984
rect 344650 388184 344706 388240
rect 345018 396072 345074 396128
rect 345110 391040 345166 391096
rect 345386 388864 345442 388920
rect 345662 399200 345718 399256
rect 345846 397976 345902 398032
rect 346214 398948 346270 398984
rect 346214 398928 346216 398948
rect 346216 398928 346268 398948
rect 346268 398928 346270 398948
rect 346122 395392 346178 395448
rect 345478 320728 345534 320784
rect 345846 381656 345902 381712
rect 346720 399880 346776 399936
rect 346766 399744 346822 399800
rect 347088 399880 347144 399936
rect 347824 399880 347880 399936
rect 346674 398948 346730 398984
rect 346674 398928 346676 398948
rect 346676 398928 346728 398948
rect 346728 398928 346730 398948
rect 346858 399336 346914 399392
rect 346398 394984 346454 395040
rect 346214 388456 346270 388512
rect 346122 320864 346178 320920
rect 347226 399492 347282 399528
rect 347226 399472 347228 399492
rect 347228 399472 347280 399492
rect 347280 399472 347282 399492
rect 347226 397704 347282 397760
rect 347410 398656 347466 398712
rect 347502 395664 347558 395720
rect 348468 399880 348524 399936
rect 347870 398112 347926 398168
rect 347778 396616 347834 396672
rect 347318 394984 347374 395040
rect 347870 394848 347926 394904
rect 347502 383288 347558 383344
rect 348330 397296 348386 397352
rect 348146 395392 348202 395448
rect 348928 399880 348984 399936
rect 348606 397568 348662 397624
rect 348422 388728 348478 388784
rect 348422 387504 348478 387560
rect 349296 399880 349352 399936
rect 349158 398792 349214 398848
rect 349250 396752 349306 396808
rect 348514 379344 348570 379400
rect 349526 388592 349582 388648
rect 349434 378800 349490 378856
rect 350860 399880 350916 399936
rect 349802 397840 349858 397896
rect 349986 398384 350042 398440
rect 349986 398248 350042 398304
rect 349986 397568 350042 397624
rect 349986 395392 350042 395448
rect 349618 321952 349674 322008
rect 349986 378664 350042 378720
rect 349986 377576 350042 377632
rect 350722 396752 350778 396808
rect 350630 393508 350686 393544
rect 350630 393488 350632 393508
rect 350632 393488 350684 393508
rect 350684 393488 350686 393508
rect 351596 399880 351652 399936
rect 351274 399472 351330 399528
rect 351090 397840 351146 397896
rect 350998 379072 351054 379128
rect 350906 373360 350962 373416
rect 351458 379208 351514 379264
rect 351826 397976 351882 398032
rect 352010 394168 352066 394224
rect 352286 398384 352342 398440
rect 352286 384376 352342 384432
rect 352194 377304 352250 377360
rect 352562 396480 352618 396536
rect 342350 219272 342406 219328
rect 340970 72392 341026 72448
rect 343638 113736 343694 113792
rect 352930 399472 352986 399528
rect 353252 399880 353308 399936
rect 353022 397432 353078 397488
rect 353206 399472 353262 399528
rect 353804 399880 353860 399936
rect 353390 398928 353446 398984
rect 353298 397432 353354 397488
rect 353574 399200 353630 399256
rect 353114 392264 353170 392320
rect 353298 390224 353354 390280
rect 354356 399880 354412 399936
rect 353850 391720 353906 391776
rect 353758 391448 353814 391504
rect 354310 395528 354366 395584
rect 354218 395256 354274 395312
rect 354034 391584 354090 391640
rect 354816 399880 354872 399936
rect 355276 399880 355332 399936
rect 354034 390224 354090 390280
rect 354310 389680 354366 389736
rect 354954 396616 355010 396672
rect 355322 399200 355378 399256
rect 355690 398792 355746 398848
rect 355598 380160 355654 380216
rect 356656 399880 356712 399936
rect 355966 397160 356022 397216
rect 355966 393624 356022 393680
rect 357116 399880 357172 399936
rect 357852 399880 357908 399936
rect 356702 398112 356758 398168
rect 356426 394440 356482 394496
rect 355322 305768 355378 305824
rect 356886 393760 356942 393816
rect 357530 392400 357586 392456
rect 358404 399880 358460 399936
rect 357990 397432 358046 397488
rect 358358 396616 358414 396672
rect 357806 387232 357862 387288
rect 357622 381520 357678 381576
rect 358542 395256 358598 395312
rect 358818 397568 358874 397624
rect 359508 399880 359564 399936
rect 359002 399200 359058 399256
rect 359186 399508 359188 399528
rect 359188 399508 359240 399528
rect 359240 399508 359242 399528
rect 359186 399472 359242 399508
rect 360060 399880 360116 399936
rect 359784 399744 359840 399800
rect 359278 396480 359334 396536
rect 359002 394984 359058 395040
rect 360888 399744 360944 399800
rect 361532 399880 361588 399936
rect 354678 64096 354734 64152
rect 351642 3712 351698 3768
rect 354034 3712 354090 3768
rect 358726 9424 358782 9480
rect 361992 399880 362048 399936
rect 361486 398792 361542 398848
rect 361486 397704 361542 397760
rect 363280 399880 363336 399936
rect 363648 399880 363704 399936
rect 364200 399880 364256 399936
rect 362866 397976 362922 398032
rect 362774 393080 362830 393136
rect 363234 394440 363290 394496
rect 364154 399472 364210 399528
rect 364062 395528 364118 395584
rect 364752 399880 364808 399936
rect 364522 395256 364578 395312
rect 364522 394984 364578 395040
rect 364338 392672 364394 392728
rect 364706 395120 364762 395176
rect 364614 373496 364670 373552
rect 365304 399880 365360 399936
rect 365120 399744 365176 399800
rect 366040 399744 366096 399800
rect 365074 399472 365130 399528
rect 365166 395936 365222 395992
rect 367236 399880 367292 399936
rect 367604 399880 367660 399936
rect 366546 398676 366602 398712
rect 366546 398656 366548 398676
rect 366548 398656 366600 398676
rect 366600 398656 366602 398676
rect 366362 397296 366418 397352
rect 366270 383152 366326 383208
rect 366638 397296 366694 397352
rect 367190 397296 367246 397352
rect 367190 395936 367246 395992
rect 367466 398112 367522 398168
rect 368708 399880 368764 399936
rect 367834 397976 367890 398032
rect 368294 397976 368350 398032
rect 368662 398520 368718 398576
rect 369168 399880 369224 399936
rect 368754 397840 368810 397896
rect 368478 392672 368534 392728
rect 368846 377440 368902 377496
rect 369536 399880 369592 399936
rect 369720 399880 369776 399936
rect 370364 399880 370420 399936
rect 370272 399744 370328 399800
rect 370640 399880 370696 399936
rect 369030 395664 369086 395720
rect 369398 391856 369454 391912
rect 369858 399200 369914 399256
rect 370042 398656 370098 398712
rect 370226 398384 370282 398440
rect 370502 399472 370558 399528
rect 370686 399200 370742 399256
rect 370594 398520 370650 398576
rect 370594 398384 370650 398440
rect 371008 399846 371064 399902
rect 370778 397704 370834 397760
rect 370686 393896 370742 393952
rect 371468 399880 371524 399936
rect 371146 399472 371202 399528
rect 371054 397840 371110 397896
rect 371652 399880 371708 399936
rect 371330 399200 371386 399256
rect 372020 399846 372076 399902
rect 371698 399200 371754 399256
rect 370686 308760 370742 308816
rect 372664 399846 372720 399902
rect 372250 398656 372306 398712
rect 373216 399880 373272 399936
rect 372526 398792 372582 398848
rect 372434 397432 372490 397488
rect 372710 399336 372766 399392
rect 372710 397840 372766 397896
rect 372710 395800 372766 395856
rect 372894 399472 372950 399528
rect 372986 398112 373042 398168
rect 373768 399880 373824 399936
rect 373354 398248 373410 398304
rect 373078 397568 373134 397624
rect 373814 399608 373870 399664
rect 373630 399200 373686 399256
rect 374182 399608 374238 399664
rect 374274 397976 374330 398032
rect 373998 392148 374054 392184
rect 373998 392128 374000 392148
rect 374000 392128 374052 392148
rect 374052 392128 374054 392148
rect 374458 398792 374514 398848
rect 374780 399880 374836 399936
rect 375056 399880 375112 399936
rect 375424 399880 375480 399936
rect 375792 399880 375848 399936
rect 374642 399508 374644 399528
rect 374644 399508 374696 399528
rect 374696 399508 374698 399528
rect 374642 399472 374698 399508
rect 374458 395256 374514 395312
rect 374918 399064 374974 399120
rect 374826 397432 374882 397488
rect 374550 370504 374606 370560
rect 374458 341536 374514 341592
rect 374826 377712 374882 377768
rect 375286 399472 375342 399528
rect 375838 399744 375894 399800
rect 375562 399608 375618 399664
rect 376252 399880 376308 399936
rect 376528 399846 376584 399902
rect 376712 399880 376768 399936
rect 376298 399608 376354 399664
rect 376022 391312 376078 391368
rect 376988 399880 377044 399936
rect 376574 399608 376630 399664
rect 376758 397568 376814 397624
rect 376666 390496 376722 390552
rect 377126 399608 377182 399664
rect 378000 399846 378056 399902
rect 378184 399880 378240 399936
rect 377494 399508 377496 399528
rect 377496 399508 377548 399528
rect 377548 399508 377550 399528
rect 377494 399472 377550 399508
rect 377862 390088 377918 390144
rect 378138 399744 378194 399800
rect 378046 397024 378102 397080
rect 378460 399744 378516 399800
rect 378736 399880 378792 399936
rect 378230 399608 378286 399664
rect 378322 395256 378378 395312
rect 377310 318960 377366 319016
rect 378598 399200 378654 399256
rect 379472 399880 379528 399936
rect 379150 397432 379206 397488
rect 379150 395256 379206 395312
rect 379748 399880 379804 399936
rect 379932 399880 379988 399936
rect 379518 397976 379574 398032
rect 380392 399846 380448 399902
rect 380576 399880 380632 399936
rect 380852 399880 380908 399936
rect 381036 399880 381092 399936
rect 379702 330520 379758 330576
rect 379610 315696 379666 315752
rect 380208 399642 380264 399698
rect 380346 399608 380402 399664
rect 380162 386688 380218 386744
rect 379150 311480 379206 311536
rect 380622 399608 380678 399664
rect 380806 399744 380862 399800
rect 381128 399744 381184 399800
rect 381266 399628 381322 399664
rect 381266 399608 381268 399628
rect 381268 399608 381320 399628
rect 381320 399608 381322 399628
rect 380806 398384 380862 398440
rect 380898 393488 380954 393544
rect 380530 390360 380586 390416
rect 380898 326304 380954 326360
rect 381174 312976 381230 313032
rect 381634 399200 381690 399256
rect 381542 385872 381598 385928
rect 381450 311752 381506 311808
rect 381082 308896 381138 308952
rect 380438 307672 380494 307728
rect 382324 399880 382380 399936
rect 382094 398112 382150 398168
rect 382094 397568 382150 397624
rect 382784 399880 382840 399936
rect 382968 399846 383024 399902
rect 383152 399880 383208 399936
rect 382186 397432 382242 397488
rect 382646 397976 382702 398032
rect 382462 342896 382518 342952
rect 361578 62736 361634 62792
rect 365810 102856 365866 102912
rect 368478 61376 368534 61432
rect 372618 58520 372674 58576
rect 379978 6432 380034 6488
rect 383198 399744 383254 399800
rect 383290 398248 383346 398304
rect 383796 399880 383852 399936
rect 383750 399744 383806 399800
rect 384072 399846 384128 399902
rect 384440 399846 384496 399902
rect 384992 399846 385048 399902
rect 383474 397568 383530 397624
rect 384118 399064 384174 399120
rect 384026 397976 384082 398032
rect 384578 398384 384634 398440
rect 384670 398112 384726 398168
rect 384854 399200 384910 399256
rect 383934 356632 383990 356688
rect 383750 340040 383806 340096
rect 384394 313112 384450 313168
rect 384946 398928 385002 398984
rect 385360 399880 385416 399936
rect 385222 399472 385278 399528
rect 385820 399880 385876 399936
rect 386280 399880 386336 399936
rect 386648 399880 386704 399936
rect 386832 399880 386888 399936
rect 387108 399880 387164 399936
rect 385498 399472 385554 399528
rect 385590 396072 385646 396128
rect 385866 398792 385922 398848
rect 385314 341400 385370 341456
rect 384946 323584 385002 323640
rect 385774 323720 385830 323776
rect 386142 399608 386198 399664
rect 386050 397840 386106 397896
rect 385866 322088 385922 322144
rect 385682 317192 385738 317248
rect 386510 399608 386566 399664
rect 386878 399472 386934 399528
rect 386878 333240 386934 333296
rect 386786 330384 386842 330440
rect 386694 327664 386750 327720
rect 386602 321544 386658 321600
rect 387062 321544 387118 321600
rect 386510 317056 386566 317112
rect 384762 300736 384818 300792
rect 384302 155216 384358 155272
rect 389546 400152 389602 400208
rect 387338 314200 387394 314256
rect 388258 398248 388314 398304
rect 388166 314336 388222 314392
rect 387982 311072 388038 311128
rect 387890 310120 387946 310176
rect 389178 306312 389234 306368
rect 390650 400016 390706 400072
rect 390834 396888 390890 396944
rect 390926 317328 390982 317384
rect 390834 315152 390890 315208
rect 390742 314472 390798 314528
rect 390558 309984 390614 310040
rect 389270 306176 389326 306232
rect 392122 397976 392178 398032
rect 393410 313928 393466 313984
rect 393318 310392 393374 310448
rect 392122 310256 392178 310312
rect 392030 309032 392086 309088
rect 391938 306040 391994 306096
rect 577502 386960 577558 387016
rect 427818 338136 427874 338192
rect 394882 303456 394938 303512
rect 395986 303456 396042 303512
rect 390650 6296 390706 6352
rect 394238 6160 394294 6216
rect 397458 21256 397514 21312
rect 400218 82048 400274 82104
rect 407210 54440 407266 54496
rect 411258 53080 411314 53136
rect 415490 9288 415546 9344
rect 418986 9152 419042 9208
rect 426438 120808 426494 120864
rect 513378 335416 513434 335472
rect 429198 14456 429254 14512
rect 477498 313928 477554 313984
rect 436834 9016 436890 9072
rect 440330 8880 440386 8936
rect 448610 117952 448666 118008
rect 462318 116456 462374 116512
rect 460938 76472 460994 76528
rect 458086 3576 458142 3632
rect 465170 3440 465226 3496
rect 472622 115096 472678 115152
rect 485778 111016 485834 111072
rect 487158 39208 487214 39264
rect 482834 3304 482890 3360
rect 496818 106800 496874 106856
rect 502338 312432 502394 312488
rect 498290 151136 498346 151192
rect 506570 105440 506626 105496
rect 510618 104080 510674 104136
rect 514850 102720 514906 102776
rect 520922 122032 520978 122088
rect 529938 149640 529994 149696
rect 528558 98640 528614 98696
rect 531410 97144 531466 97200
rect 536838 151000 536894 151056
rect 539598 120672 539654 120728
rect 542358 95784 542414 95840
rect 543738 148280 543794 148336
rect 549258 93064 549314 93120
rect 552662 311072 552718 311128
rect 570602 304952 570658 305008
rect 580262 378392 580318 378448
rect 580262 366424 580318 366480
rect 580170 365064 580226 365120
rect 579618 312024 579674 312080
rect 580170 298732 580172 298752
rect 580172 298732 580224 298752
rect 580224 298732 580226 298752
rect 580170 298696 580226 298732
rect 579618 245556 579620 245576
rect 579620 245556 579672 245576
rect 579672 245556 579674 245576
rect 579618 245520 579674 245556
rect 579618 232328 579674 232384
rect 579618 209072 579674 209128
rect 579618 205672 579674 205728
rect 579618 192480 579674 192536
rect 579894 152632 579950 152688
rect 580538 366288 580594 366344
rect 580446 364928 580502 364984
rect 580354 258848 580410 258904
rect 580354 200640 580410 200696
rect 580262 139304 580318 139360
rect 580170 112784 580226 112840
rect 580262 100000 580318 100056
rect 580170 99456 580226 99512
rect 580262 86128 580318 86184
rect 580262 71032 580318 71088
rect 580262 46280 580318 46336
rect 580078 19760 580134 19816
rect 580722 351872 580778 351928
rect 580722 325216 580778 325272
rect 580630 272176 580686 272232
rect 580538 219000 580594 219056
rect 580538 209208 580594 209264
rect 580446 179152 580502 179208
rect 580722 208936 580778 208992
rect 580722 165824 580778 165880
rect 580538 125976 580594 126032
rect 580354 6568 580410 6624
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580257 683906 580323 683909
rect 583520 683906 584960 683996
rect 580257 683904 584960 683906
rect 580257 683848 580262 683904
rect 580318 683848 584960 683904
rect 580257 683846 584960 683848
rect 580257 683843 580323 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3417 671258 3483 671261
rect -960 671256 3483 671258
rect -960 671200 3422 671256
rect 3478 671200 3483 671256
rect -960 671198 3483 671200
rect -960 671108 480 671198
rect 3417 671195 3483 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 2773 658202 2839 658205
rect -960 658200 2839 658202
rect -960 658144 2778 658200
rect 2834 658144 2839 658200
rect -960 658142 2839 658144
rect -960 658052 480 658142
rect 2773 658139 2839 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 579981 630866 580047 630869
rect 583520 630866 584960 630956
rect 579981 630864 584960 630866
rect 579981 630808 579986 630864
rect 580042 630808 584960 630864
rect 579981 630806 584960 630808
rect 579981 630803 580047 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3417 619170 3483 619173
rect -960 619168 3483 619170
rect -960 619112 3422 619168
rect 3478 619112 3483 619168
rect -960 619110 3483 619112
rect -960 619020 480 619110
rect 3417 619107 3483 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3509 606114 3575 606117
rect -960 606112 3575 606114
rect -960 606056 3514 606112
rect 3570 606056 3575 606112
rect -960 606054 3575 606056
rect -960 605964 480 606054
rect 3509 606051 3575 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580165 591018 580231 591021
rect 583520 591018 584960 591108
rect 580165 591016 584960 591018
rect 580165 590960 580170 591016
rect 580226 590960 584960 591016
rect 580165 590958 584960 590960
rect 580165 590955 580231 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3233 566946 3299 566949
rect -960 566944 3299 566946
rect -960 566888 3238 566944
rect 3294 566888 3299 566944
rect -960 566886 3299 566888
rect -960 566796 480 566886
rect 3233 566883 3299 566886
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3325 553890 3391 553893
rect -960 553888 3391 553890
rect -960 553832 3330 553888
rect 3386 553832 3391 553888
rect -960 553830 3391 553832
rect -960 553740 480 553830
rect 3325 553827 3391 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 579889 537842 579955 537845
rect 583520 537842 584960 537932
rect 579889 537840 584960 537842
rect 579889 537784 579894 537840
rect 579950 537784 584960 537840
rect 579889 537782 584960 537784
rect 579889 537779 579955 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 2957 527914 3023 527917
rect -960 527912 3023 527914
rect -960 527856 2962 527912
rect 3018 527856 3023 527912
rect -960 527854 3023 527856
rect -960 527764 480 527854
rect 2957 527851 3023 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3509 514858 3575 514861
rect -960 514856 3575 514858
rect -960 514800 3514 514856
rect 3570 514800 3575 514856
rect -960 514798 3575 514800
rect -960 514708 480 514798
rect 3509 514795 3575 514798
rect 580349 511322 580415 511325
rect 583520 511322 584960 511412
rect 580349 511320 584960 511322
rect 580349 511264 580354 511320
rect 580410 511264 584960 511320
rect 580349 511262 584960 511264
rect 580349 511259 580415 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3049 501802 3115 501805
rect -960 501800 3115 501802
rect -960 501744 3054 501800
rect 3110 501744 3115 501800
rect -960 501742 3115 501744
rect -960 501652 480 501742
rect 3049 501739 3115 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3049 475690 3115 475693
rect -960 475688 3115 475690
rect -960 475632 3054 475688
rect 3110 475632 3115 475688
rect -960 475630 3115 475632
rect -960 475540 480 475630
rect 3049 475627 3115 475630
rect 580073 471474 580139 471477
rect 583520 471474 584960 471564
rect 580073 471472 584960 471474
rect 580073 471416 580078 471472
rect 580134 471416 584960 471472
rect 580073 471414 584960 471416
rect 580073 471411 580139 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3509 462634 3575 462637
rect -960 462632 3575 462634
rect -960 462576 3514 462632
rect 3570 462576 3575 462632
rect -960 462574 3575 462576
rect -960 462484 480 462574
rect 3509 462571 3575 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect 337469 454202 337535 454205
rect 371325 454202 371391 454205
rect 337469 454200 371391 454202
rect 337469 454144 337474 454200
rect 337530 454144 371330 454200
rect 371386 454144 371391 454200
rect 337469 454142 371391 454144
rect 337469 454139 337535 454142
rect 371325 454139 371391 454142
rect 337653 454066 337719 454069
rect 372797 454066 372863 454069
rect 337653 454064 372863 454066
rect 337653 454008 337658 454064
rect 337714 454008 372802 454064
rect 372858 454008 372863 454064
rect 337653 454006 372863 454008
rect 337653 454003 337719 454006
rect 372797 454003 372863 454006
rect 308397 452842 308463 452845
rect 368013 452842 368079 452845
rect 308397 452840 368079 452842
rect 308397 452784 308402 452840
rect 308458 452784 368018 452840
rect 368074 452784 368079 452840
rect 308397 452782 368079 452784
rect 308397 452779 308463 452782
rect 368013 452779 368079 452782
rect 279918 452644 279924 452708
rect 279988 452706 279994 452708
rect 347773 452706 347839 452709
rect 279988 452704 347839 452706
rect 279988 452648 347778 452704
rect 347834 452648 347839 452704
rect 279988 452646 347839 452648
rect 279988 452644 279994 452646
rect 347773 452643 347839 452646
rect 361665 452570 361731 452573
rect 362217 452570 362283 452573
rect 361665 452568 362283 452570
rect 361665 452512 361670 452568
rect 361726 452512 362222 452568
rect 362278 452512 362283 452568
rect 361665 452510 362283 452512
rect 361665 452507 361731 452510
rect 362217 452507 362283 452510
rect 368565 452570 368631 452573
rect 369485 452570 369551 452573
rect 372613 452572 372679 452573
rect 374085 452572 374151 452573
rect 372613 452570 372660 452572
rect 368565 452568 369551 452570
rect 368565 452512 368570 452568
rect 368626 452512 369490 452568
rect 369546 452512 369551 452568
rect 368565 452510 369551 452512
rect 372568 452568 372660 452570
rect 372568 452512 372618 452568
rect 372568 452510 372660 452512
rect 368565 452507 368631 452510
rect 369485 452507 369551 452510
rect 372613 452508 372660 452510
rect 372724 452508 372730 452572
rect 374085 452570 374132 452572
rect 374040 452568 374132 452570
rect 374040 452512 374090 452568
rect 374040 452510 374132 452512
rect 374085 452508 374132 452510
rect 374196 452508 374202 452572
rect 372613 452507 372679 452508
rect 374085 452507 374151 452508
rect 343582 452100 343588 452164
rect 343652 452162 343658 452164
rect 361665 452162 361731 452165
rect 343652 452160 361731 452162
rect 343652 452104 361670 452160
rect 361726 452104 361731 452160
rect 343652 452102 361731 452104
rect 343652 452100 343658 452102
rect 361665 452099 361731 452102
rect 278630 451828 278636 451892
rect 278700 451890 278706 451892
rect 345565 451890 345631 451893
rect 278700 451888 345631 451890
rect 278700 451832 345570 451888
rect 345626 451832 345631 451888
rect 278700 451830 345631 451832
rect 278700 451828 278706 451830
rect 345565 451827 345631 451830
rect 340873 451754 340939 451757
rect 371417 451754 371483 451757
rect 340873 451752 371483 451754
rect 340873 451696 340878 451752
rect 340934 451696 371422 451752
rect 371478 451696 371483 451752
rect 340873 451694 371483 451696
rect 340873 451691 340939 451694
rect 371417 451691 371483 451694
rect 300117 451618 300183 451621
rect 345933 451618 345999 451621
rect 300117 451616 345999 451618
rect 300117 451560 300122 451616
rect 300178 451560 345938 451616
rect 345994 451560 345999 451616
rect 300117 451558 345999 451560
rect 300117 451555 300183 451558
rect 345933 451555 345999 451558
rect 357382 451556 357388 451620
rect 357452 451618 357458 451620
rect 358629 451618 358695 451621
rect 357452 451616 358695 451618
rect 357452 451560 358634 451616
rect 358690 451560 358695 451616
rect 357452 451558 358695 451560
rect 357452 451556 357458 451558
rect 358629 451555 358695 451558
rect 280705 451482 280771 451485
rect 345197 451482 345263 451485
rect 280705 451480 345263 451482
rect 280705 451424 280710 451480
rect 280766 451424 345202 451480
rect 345258 451424 345263 451480
rect 280705 451422 345263 451424
rect 280705 451419 280771 451422
rect 345197 451419 345263 451422
rect 346342 451420 346348 451484
rect 346412 451482 346418 451484
rect 368565 451482 368631 451485
rect 346412 451480 368631 451482
rect 346412 451424 368570 451480
rect 368626 451424 368631 451480
rect 346412 451422 368631 451424
rect 346412 451420 346418 451422
rect 368565 451419 368631 451422
rect 368974 451420 368980 451484
rect 369044 451482 369050 451484
rect 373993 451482 374059 451485
rect 369044 451480 374059 451482
rect 369044 451424 373998 451480
rect 374054 451424 374059 451480
rect 369044 451422 374059 451424
rect 369044 451420 369050 451422
rect 373993 451419 374059 451422
rect 347630 451284 347636 451348
rect 347700 451346 347706 451348
rect 352925 451346 352991 451349
rect 347700 451344 352991 451346
rect 347700 451288 352930 451344
rect 352986 451288 352991 451344
rect 347700 451286 352991 451288
rect 347700 451284 347706 451286
rect 352925 451283 352991 451286
rect 355174 451284 355180 451348
rect 355244 451346 355250 451348
rect 359549 451346 359615 451349
rect 355244 451344 359615 451346
rect 355244 451288 359554 451344
rect 359610 451288 359615 451344
rect 355244 451286 359615 451288
rect 355244 451284 355250 451286
rect 359549 451283 359615 451286
rect 375966 451284 375972 451348
rect 376036 451346 376042 451348
rect 378685 451346 378751 451349
rect 376036 451344 378751 451346
rect 376036 451288 378690 451344
rect 378746 451288 378751 451344
rect 376036 451286 378751 451288
rect 376036 451284 376042 451286
rect 378685 451283 378751 451286
rect 334985 450258 335051 450261
rect 370083 450258 370149 450261
rect 334985 450256 370149 450258
rect 334985 450200 334990 450256
rect 335046 450200 370088 450256
rect 370144 450200 370149 450256
rect 334985 450198 370149 450200
rect 334985 450195 335051 450198
rect 370083 450195 370149 450198
rect 314009 450122 314075 450125
rect 373395 450122 373461 450125
rect 314009 450120 373461 450122
rect 314009 450064 314014 450120
rect 314070 450064 373400 450120
rect 373456 450064 373461 450120
rect 314009 450062 373461 450064
rect 314009 450059 314075 450062
rect 373395 450059 373461 450062
rect 300209 449986 300275 449989
rect 360147 449986 360213 449989
rect 300209 449984 360213 449986
rect 300209 449928 300214 449984
rect 300270 449928 360152 449984
rect 360208 449928 360213 449984
rect 300209 449926 360213 449928
rect 300209 449923 300275 449926
rect 360147 449923 360213 449926
rect 339401 449714 339467 449717
rect 347267 449714 347333 449717
rect 339401 449712 347333 449714
rect -960 449578 480 449668
rect 339401 449656 339406 449712
rect 339462 449656 347272 449712
rect 347328 449656 347333 449712
rect 339401 449654 347333 449656
rect 339401 449651 339467 449654
rect 347267 449651 347333 449654
rect 3049 449578 3115 449581
rect 346531 449578 346597 449581
rect 371923 449578 371989 449581
rect -960 449576 3115 449578
rect -960 449520 3054 449576
rect 3110 449520 3115 449576
rect -960 449518 3115 449520
rect -960 449428 480 449518
rect 3049 449515 3115 449518
rect 340830 449576 346597 449578
rect 340830 449520 346536 449576
rect 346592 449520 346597 449576
rect 340830 449518 346597 449520
rect 340830 449306 340890 449518
rect 346531 449515 346597 449518
rect 354630 449576 371989 449578
rect 354630 449520 371928 449576
rect 371984 449520 371989 449576
rect 354630 449518 371989 449520
rect 343950 449380 343956 449444
rect 344020 449442 344026 449444
rect 344461 449442 344527 449445
rect 344020 449440 344527 449442
rect 344020 449384 344466 449440
rect 344522 449384 344527 449440
rect 344020 449382 344527 449384
rect 344020 449380 344026 449382
rect 344461 449379 344527 449382
rect 345197 449444 345263 449445
rect 345197 449440 345244 449444
rect 345308 449442 345314 449444
rect 349337 449442 349403 449445
rect 353385 449444 353451 449445
rect 349654 449442 349660 449444
rect 345197 449384 345202 449440
rect 345197 449380 345244 449384
rect 345308 449382 345354 449442
rect 349337 449440 349660 449442
rect 349337 449384 349342 449440
rect 349398 449384 349660 449440
rect 349337 449382 349660 449384
rect 345308 449380 345314 449382
rect 345197 449379 345263 449380
rect 349337 449379 349403 449382
rect 349654 449380 349660 449382
rect 349724 449380 349730 449444
rect 353334 449442 353340 449444
rect 353294 449382 353340 449442
rect 353404 449440 353451 449444
rect 353446 449384 353451 449440
rect 353334 449380 353340 449382
rect 353404 449380 353451 449384
rect 353385 449379 353451 449380
rect 335310 449246 340890 449306
rect 343955 449306 344021 449309
rect 344870 449306 344876 449308
rect 343955 449304 344876 449306
rect 343955 449248 343960 449304
rect 344016 449248 344876 449304
rect 343955 449246 344876 449248
rect 281073 449170 281139 449173
rect 335310 449170 335370 449246
rect 343955 449243 344021 449246
rect 344870 449244 344876 449246
rect 344940 449244 344946 449308
rect 346899 449304 346965 449309
rect 346899 449248 346904 449304
rect 346960 449248 346965 449304
rect 346899 449243 346965 449248
rect 281073 449168 335370 449170
rect 281073 449112 281078 449168
rect 281134 449112 335370 449168
rect 281073 449110 335370 449112
rect 281073 449107 281139 449110
rect 286317 449034 286383 449037
rect 346902 449034 346962 449243
rect 286317 449032 346962 449034
rect 286317 448976 286322 449032
rect 286378 448976 346962 449032
rect 286317 448974 346962 448976
rect 286317 448971 286383 448974
rect 312537 448898 312603 448901
rect 354630 448898 354690 449518
rect 371923 449515 371989 449518
rect 357566 449380 357572 449444
rect 357636 449442 357642 449444
rect 358077 449442 358143 449445
rect 357636 449440 358143 449442
rect 357636 449384 358082 449440
rect 358138 449384 358143 449440
rect 357636 449382 358143 449384
rect 357636 449380 357642 449382
rect 358077 449379 358143 449382
rect 370446 449380 370452 449444
rect 370516 449442 370522 449444
rect 370589 449442 370655 449445
rect 370516 449440 370655 449442
rect 370516 449384 370594 449440
rect 370650 449384 370655 449440
rect 370516 449382 370655 449384
rect 370516 449380 370522 449382
rect 370589 449379 370655 449382
rect 371550 449380 371556 449444
rect 371620 449442 371626 449444
rect 372061 449442 372127 449445
rect 371620 449440 372127 449442
rect 371620 449384 372066 449440
rect 372122 449384 372127 449440
rect 371620 449382 372127 449384
rect 371620 449380 371626 449382
rect 372061 449379 372127 449382
rect 372654 449380 372660 449444
rect 372724 449442 372730 449444
rect 372797 449442 372863 449445
rect 372724 449440 372863 449442
rect 372724 449384 372802 449440
rect 372858 449384 372863 449440
rect 372724 449382 372863 449384
rect 372724 449380 372730 449382
rect 372797 449379 372863 449382
rect 374126 449380 374132 449444
rect 374196 449442 374202 449444
rect 375005 449442 375071 449445
rect 374196 449440 375071 449442
rect 374196 449384 375010 449440
rect 375066 449384 375071 449440
rect 374196 449382 375071 449384
rect 374196 449380 374202 449382
rect 375005 449379 375071 449382
rect 382222 449380 382228 449444
rect 382292 449442 382298 449444
rect 383101 449442 383167 449445
rect 382292 449440 383167 449442
rect 382292 449384 383106 449440
rect 383162 449384 383167 449440
rect 382292 449382 383167 449384
rect 382292 449380 382298 449382
rect 383101 449379 383167 449382
rect 383837 449444 383903 449445
rect 384297 449444 384363 449445
rect 383837 449440 383884 449444
rect 383948 449442 383954 449444
rect 384246 449442 384252 449444
rect 383837 449384 383842 449440
rect 383837 449380 383884 449384
rect 383948 449382 383994 449442
rect 384206 449382 384252 449442
rect 384316 449440 384363 449444
rect 384358 449384 384363 449440
rect 383948 449380 383954 449382
rect 384246 449380 384252 449382
rect 384316 449380 384363 449384
rect 385350 449380 385356 449444
rect 385420 449442 385426 449444
rect 385677 449442 385743 449445
rect 385420 449440 385743 449442
rect 385420 449384 385682 449440
rect 385738 449384 385743 449440
rect 385420 449382 385743 449384
rect 385420 449380 385426 449382
rect 383837 449379 383903 449380
rect 384297 449379 384363 449380
rect 385677 449379 385743 449382
rect 368979 449304 369045 449309
rect 368979 449248 368984 449304
rect 369040 449248 369045 449304
rect 368979 449243 369045 449248
rect 373942 449244 373948 449308
rect 374012 449306 374018 449308
rect 374867 449306 374933 449309
rect 374012 449304 374933 449306
rect 374012 449248 374872 449304
rect 374928 449248 374933 449304
rect 374012 449246 374933 449248
rect 374012 449244 374018 449246
rect 374867 449243 374933 449246
rect 382958 449244 382964 449308
rect 383028 449306 383034 449308
rect 385539 449306 385605 449309
rect 383028 449304 385605 449306
rect 383028 449248 385544 449304
rect 385600 449248 385605 449304
rect 383028 449246 385605 449248
rect 383028 449244 383034 449246
rect 385539 449243 385605 449246
rect 312537 448896 354690 448898
rect 312537 448840 312542 448896
rect 312598 448840 354690 448896
rect 312537 448838 354690 448840
rect 312537 448835 312603 448838
rect 340229 448626 340295 448629
rect 368982 448626 369042 449243
rect 340229 448624 369042 448626
rect 340229 448568 340234 448624
rect 340290 448568 369042 448624
rect 340229 448566 369042 448568
rect 340229 448563 340295 448566
rect 309777 447810 309843 447813
rect 346342 447810 346348 447812
rect 309777 447808 346348 447810
rect 309777 447752 309782 447808
rect 309838 447752 346348 447808
rect 309777 447750 346348 447752
rect 309777 447747 309843 447750
rect 346342 447748 346348 447750
rect 346412 447748 346418 447812
rect 301589 446450 301655 446453
rect 343582 446450 343588 446452
rect 301589 446448 343588 446450
rect 301589 446392 301594 446448
rect 301650 446392 343588 446448
rect 301589 446390 343588 446392
rect 301589 446387 301655 446390
rect 343582 446388 343588 446390
rect 343652 446388 343658 446452
rect 284477 444954 284543 444957
rect 343950 444954 343956 444956
rect 284477 444952 343956 444954
rect 284477 444896 284482 444952
rect 284538 444896 343956 444952
rect 284477 444894 343956 444896
rect 284477 444891 284543 444894
rect 343950 444892 343956 444894
rect 344020 444892 344026 444956
rect 583520 444668 584960 444908
rect 291929 439514 291995 439517
rect 342437 439514 342503 439517
rect 291929 439512 342503 439514
rect 291929 439456 291934 439512
rect 291990 439456 342442 439512
rect 342498 439456 342503 439512
rect 291929 439454 342503 439456
rect 291929 439451 291995 439454
rect 342437 439451 342503 439454
rect 340965 438290 341031 438293
rect 341885 438290 341951 438293
rect 340965 438288 341951 438290
rect 340965 438232 340970 438288
rect 341026 438232 341890 438288
rect 341946 438232 341951 438288
rect 340965 438230 341951 438232
rect 340965 438227 341031 438230
rect 341885 438227 341951 438230
rect 340965 436794 341031 436797
rect 341793 436794 341859 436797
rect 340965 436792 341859 436794
rect -960 436508 480 436748
rect 340965 436736 340970 436792
rect 341026 436736 341798 436792
rect 341854 436736 341859 436792
rect 340965 436734 341859 436736
rect 340965 436731 341031 436734
rect 341793 436731 341859 436734
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect 340965 428498 341031 428501
rect 341701 428498 341767 428501
rect 340965 428496 341767 428498
rect 340965 428440 340970 428496
rect 341026 428440 341706 428496
rect 341762 428440 341767 428496
rect 340965 428438 341767 428440
rect 340965 428435 341031 428438
rect 341701 428435 341767 428438
rect -960 423602 480 423692
rect 3509 423602 3575 423605
rect -960 423600 3575 423602
rect -960 423544 3514 423600
rect 3570 423544 3575 423600
rect -960 423542 3575 423544
rect -960 423452 480 423542
rect 3509 423539 3575 423542
rect 580257 418298 580323 418301
rect 583520 418298 584960 418388
rect 580257 418296 584960 418298
rect 580257 418240 580262 418296
rect 580318 418240 584960 418296
rect 580257 418238 584960 418240
rect 580257 418235 580323 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3417 410546 3483 410549
rect -960 410544 3483 410546
rect -960 410488 3422 410544
rect 3478 410488 3483 410544
rect -960 410486 3483 410488
rect -960 410396 480 410486
rect 3417 410483 3483 410486
rect 340965 405786 341031 405789
rect 341609 405786 341675 405789
rect 340965 405784 341675 405786
rect 340965 405728 340970 405784
rect 341026 405728 341614 405784
rect 341670 405728 341675 405784
rect 340965 405726 341675 405728
rect 340965 405723 341031 405726
rect 341609 405723 341675 405726
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect 275921 403066 275987 403069
rect 342069 403066 342135 403069
rect 275921 403064 342135 403066
rect 275921 403008 275926 403064
rect 275982 403008 342074 403064
rect 342130 403008 342135 403064
rect 275921 403006 342135 403008
rect 275921 403003 275987 403006
rect 342069 403003 342135 403006
rect 266169 402114 266235 402117
rect 341977 402114 342043 402117
rect 266169 402112 342043 402114
rect 266169 402056 266174 402112
rect 266230 402056 341982 402112
rect 342038 402056 342043 402112
rect 266169 402054 342043 402056
rect 266169 402051 266235 402054
rect 341977 402051 342043 402054
rect 285029 401978 285095 401981
rect 345238 401978 345244 401980
rect 285029 401976 345244 401978
rect 285029 401920 285034 401976
rect 285090 401920 345244 401976
rect 285029 401918 345244 401920
rect 285029 401915 285095 401918
rect 345238 401916 345244 401918
rect 345308 401916 345314 401980
rect 280061 401842 280127 401845
rect 352782 401842 352788 401844
rect 280061 401840 352788 401842
rect 280061 401784 280066 401840
rect 280122 401784 352788 401840
rect 280061 401782 352788 401784
rect 280061 401779 280127 401782
rect 352782 401780 352788 401782
rect 352852 401780 352858 401844
rect 313917 401298 313983 401301
rect 368974 401298 368980 401300
rect 313917 401296 368980 401298
rect 313917 401240 313922 401296
rect 313978 401240 368980 401296
rect 313917 401238 368980 401240
rect 313917 401235 313983 401238
rect 368974 401236 368980 401238
rect 369044 401236 369050 401300
rect 319713 401162 319779 401165
rect 375966 401162 375972 401164
rect 319713 401160 375972 401162
rect 319713 401104 319718 401160
rect 319774 401104 375972 401160
rect 319713 401102 375972 401104
rect 319713 401099 319779 401102
rect 375966 401100 375972 401102
rect 376036 401100 376042 401164
rect 298921 401026 298987 401029
rect 357566 401026 357572 401028
rect 298921 401024 357572 401026
rect 298921 400968 298926 401024
rect 298982 400968 357572 401024
rect 298921 400966 357572 400968
rect 298921 400963 298987 400966
rect 357566 400964 357572 400966
rect 357636 400964 357642 401028
rect 293309 400890 293375 400893
rect 347630 400890 347636 400892
rect 293309 400888 347636 400890
rect 293309 400832 293314 400888
rect 293370 400832 347636 400888
rect 293309 400830 347636 400832
rect 293309 400827 293375 400830
rect 347630 400828 347636 400830
rect 347700 400890 347706 400892
rect 580717 400890 580783 400893
rect 347700 400888 580783 400890
rect 347700 400832 580722 400888
rect 580778 400832 580783 400888
rect 347700 400830 580783 400832
rect 347700 400828 347706 400830
rect 580717 400827 580783 400830
rect 341701 400754 341767 400757
rect 353518 400754 353524 400756
rect 341701 400752 353524 400754
rect 341701 400696 341706 400752
rect 341762 400696 353524 400752
rect 341701 400694 353524 400696
rect 341701 400691 341767 400694
rect 353518 400692 353524 400694
rect 353588 400692 353594 400756
rect 269021 400618 269087 400621
rect 343214 400618 343220 400620
rect 269021 400616 343220 400618
rect 269021 400560 269026 400616
rect 269082 400560 343220 400616
rect 269021 400558 343220 400560
rect 269021 400555 269087 400558
rect 343214 400556 343220 400558
rect 343284 400556 343290 400620
rect 348550 400556 348556 400620
rect 348620 400618 348626 400620
rect 354254 400618 354260 400620
rect 348620 400558 354260 400618
rect 348620 400556 348626 400558
rect 354254 400556 354260 400558
rect 354324 400556 354330 400620
rect 335905 400482 335971 400485
rect 385718 400482 385724 400484
rect 335905 400480 385724 400482
rect 335905 400424 335910 400480
rect 335966 400424 385724 400480
rect 335905 400422 385724 400424
rect 335905 400419 335971 400422
rect 385718 400420 385724 400422
rect 385788 400420 385794 400484
rect 336549 400346 336615 400349
rect 381302 400346 381308 400348
rect 336549 400344 381308 400346
rect 336549 400288 336554 400344
rect 336610 400288 381308 400344
rect 336549 400286 381308 400288
rect 336549 400283 336615 400286
rect 381302 400284 381308 400286
rect 381372 400284 381378 400348
rect 355174 400210 355180 400212
rect 335310 400150 355180 400210
rect 300301 400074 300367 400077
rect 335310 400074 335370 400150
rect 355174 400148 355180 400150
rect 355244 400148 355250 400212
rect 389541 400210 389607 400213
rect 367050 400150 379530 400210
rect 300301 400072 335370 400074
rect 300301 400016 300306 400072
rect 300362 400016 335370 400072
rect 300301 400014 335370 400016
rect 341609 400074 341675 400077
rect 344870 400074 344876 400076
rect 341609 400072 344876 400074
rect 341609 400016 341614 400072
rect 341670 400016 344876 400072
rect 341609 400014 344876 400016
rect 300301 400011 300367 400014
rect 341609 400011 341675 400014
rect 344870 400012 344876 400014
rect 344940 400074 344946 400076
rect 348550 400074 348556 400076
rect 344940 400014 348556 400074
rect 344940 400012 344946 400014
rect 348550 400012 348556 400014
rect 348620 400012 348626 400076
rect 351310 400012 351316 400076
rect 351380 400074 351386 400076
rect 357382 400074 357388 400076
rect 351380 400014 357388 400074
rect 351380 400012 351386 400014
rect 357382 400012 357388 400014
rect 357452 400012 357458 400076
rect 359230 400014 365730 400074
rect 323761 399938 323827 399941
rect 346526 399938 346532 399940
rect 323761 399936 346532 399938
rect 323761 399880 323766 399936
rect 323822 399880 346532 399936
rect 323761 399878 346532 399880
rect 323761 399875 323827 399878
rect 346526 399876 346532 399878
rect 346596 399876 346602 399940
rect 346715 399938 346781 399941
rect 347083 399940 347149 399941
rect 347819 399940 347885 399941
rect 346894 399938 346900 399940
rect 346715 399936 346900 399938
rect 346715 399880 346720 399936
rect 346776 399880 346900 399936
rect 346715 399878 346900 399880
rect 346715 399875 346781 399878
rect 346894 399876 346900 399878
rect 346964 399876 346970 399940
rect 347078 399876 347084 399940
rect 347148 399938 347154 399940
rect 347814 399938 347820 399940
rect 347148 399878 347240 399938
rect 347728 399878 347820 399938
rect 347148 399876 347154 399878
rect 347814 399876 347820 399878
rect 347884 399876 347890 399940
rect 348182 399876 348188 399940
rect 348252 399938 348258 399940
rect 348463 399938 348529 399941
rect 348252 399936 348529 399938
rect 348252 399880 348468 399936
rect 348524 399880 348529 399936
rect 348252 399878 348529 399880
rect 348252 399876 348258 399878
rect 347083 399875 347149 399876
rect 347819 399875 347885 399876
rect 348463 399875 348529 399878
rect 348734 399876 348740 399940
rect 348804 399938 348810 399940
rect 348923 399938 348989 399941
rect 348804 399936 348989 399938
rect 348804 399880 348928 399936
rect 348984 399880 348989 399936
rect 348804 399878 348989 399880
rect 348804 399876 348810 399878
rect 348923 399875 348989 399878
rect 349291 399938 349357 399941
rect 349838 399938 349844 399940
rect 349291 399936 349844 399938
rect 349291 399880 349296 399936
rect 349352 399880 349844 399936
rect 349291 399878 349844 399880
rect 349291 399875 349357 399878
rect 349838 399876 349844 399878
rect 349908 399876 349914 399940
rect 350206 399876 350212 399940
rect 350276 399938 350282 399940
rect 350855 399938 350921 399941
rect 350276 399936 350921 399938
rect 350276 399880 350860 399936
rect 350916 399880 350921 399936
rect 350276 399878 350921 399880
rect 350276 399876 350282 399878
rect 350855 399875 350921 399878
rect 351126 399876 351132 399940
rect 351196 399938 351202 399940
rect 351591 399938 351657 399941
rect 351196 399936 351657 399938
rect 351196 399880 351596 399936
rect 351652 399880 351657 399936
rect 351196 399878 351657 399880
rect 351196 399876 351202 399878
rect 351591 399875 351657 399878
rect 352414 399876 352420 399940
rect 352484 399938 352490 399940
rect 353247 399938 353313 399941
rect 352484 399936 353313 399938
rect 352484 399880 353252 399936
rect 353308 399880 353313 399936
rect 352484 399878 353313 399880
rect 352484 399876 352490 399878
rect 353247 399875 353313 399878
rect 353518 399876 353524 399940
rect 353588 399938 353594 399940
rect 353799 399938 353865 399941
rect 354351 399940 354417 399941
rect 354811 399940 354877 399941
rect 354300 399938 354306 399940
rect 353588 399936 353865 399938
rect 353588 399880 353804 399936
rect 353860 399880 353865 399936
rect 353588 399878 353865 399880
rect 354260 399878 354306 399938
rect 354370 399936 354417 399940
rect 354806 399938 354812 399940
rect 354412 399880 354417 399936
rect 353588 399876 353594 399878
rect 353799 399875 353865 399878
rect 354300 399876 354306 399878
rect 354370 399876 354417 399880
rect 354720 399878 354812 399938
rect 354806 399876 354812 399878
rect 354876 399876 354882 399940
rect 354990 399876 354996 399940
rect 355060 399938 355066 399940
rect 355271 399938 355337 399941
rect 355060 399936 355337 399938
rect 355060 399880 355276 399936
rect 355332 399880 355337 399936
rect 355060 399878 355337 399880
rect 355060 399876 355066 399878
rect 354351 399875 354417 399876
rect 354811 399875 354877 399876
rect 355271 399875 355337 399878
rect 356462 399876 356468 399940
rect 356532 399938 356538 399940
rect 356651 399938 356717 399941
rect 356532 399936 356717 399938
rect 356532 399880 356656 399936
rect 356712 399880 356717 399936
rect 356532 399878 356717 399880
rect 356532 399876 356538 399878
rect 356651 399875 356717 399878
rect 356830 399876 356836 399940
rect 356900 399938 356906 399940
rect 357111 399938 357177 399941
rect 356900 399936 357177 399938
rect 356900 399880 357116 399936
rect 357172 399880 357177 399936
rect 356900 399878 357177 399880
rect 356900 399876 356906 399878
rect 357111 399875 357177 399878
rect 357566 399876 357572 399940
rect 357636 399938 357642 399940
rect 357847 399938 357913 399941
rect 357636 399936 357913 399938
rect 357636 399880 357852 399936
rect 357908 399880 357913 399936
rect 357636 399878 357913 399880
rect 357636 399876 357642 399878
rect 357847 399875 357913 399878
rect 358118 399876 358124 399940
rect 358188 399938 358194 399940
rect 358399 399938 358465 399941
rect 358188 399936 358465 399938
rect 358188 399880 358404 399936
rect 358460 399880 358465 399936
rect 358188 399878 358465 399880
rect 358188 399876 358194 399878
rect 358399 399875 358465 399878
rect 358670 399876 358676 399940
rect 358740 399938 358746 399940
rect 359038 399938 359044 399940
rect 358740 399878 359044 399938
rect 358740 399876 358746 399878
rect 359038 399876 359044 399878
rect 359108 399876 359114 399940
rect 298737 399802 298803 399805
rect 346761 399804 346827 399805
rect 346342 399802 346348 399804
rect 298737 399800 346348 399802
rect 298737 399744 298742 399800
rect 298798 399744 346348 399800
rect 298737 399742 346348 399744
rect 298737 399739 298803 399742
rect 346342 399740 346348 399742
rect 346412 399740 346418 399804
rect 346710 399802 346716 399804
rect 346670 399742 346716 399802
rect 346780 399800 346827 399804
rect 346822 399744 346827 399800
rect 346710 399740 346716 399742
rect 346780 399740 346827 399744
rect 347262 399740 347268 399804
rect 347332 399802 347338 399804
rect 359230 399802 359290 400014
rect 359503 399938 359569 399941
rect 359774 399938 359780 399940
rect 359503 399936 359780 399938
rect 359503 399880 359508 399936
rect 359564 399880 359780 399936
rect 359503 399878 359780 399880
rect 359503 399875 359569 399878
rect 359774 399876 359780 399878
rect 359844 399876 359850 399940
rect 360055 399938 360121 399941
rect 360326 399938 360332 399940
rect 360055 399936 360332 399938
rect 360055 399880 360060 399936
rect 360116 399880 360332 399936
rect 360055 399878 360332 399880
rect 360055 399875 360121 399878
rect 360326 399876 360332 399878
rect 360396 399876 360402 399940
rect 361062 399876 361068 399940
rect 361132 399938 361138 399940
rect 361527 399938 361593 399941
rect 361132 399936 361593 399938
rect 361132 399880 361532 399936
rect 361588 399880 361593 399936
rect 361132 399878 361593 399880
rect 361132 399876 361138 399878
rect 361527 399875 361593 399878
rect 361987 399936 362053 399941
rect 363275 399940 363341 399941
rect 363270 399938 363276 399940
rect 361987 399880 361992 399936
rect 362048 399880 362053 399936
rect 361987 399875 362053 399880
rect 363184 399878 363276 399938
rect 363270 399876 363276 399878
rect 363340 399876 363346 399940
rect 363643 399938 363709 399941
rect 363822 399938 363828 399940
rect 363643 399936 363828 399938
rect 363643 399880 363648 399936
rect 363704 399880 363828 399936
rect 363643 399878 363828 399880
rect 363275 399875 363341 399876
rect 363643 399875 363709 399878
rect 363822 399876 363828 399878
rect 363892 399876 363898 399940
rect 364195 399938 364261 399941
rect 364014 399936 364261 399938
rect 364014 399880 364200 399936
rect 364256 399880 364261 399936
rect 364014 399878 364261 399880
rect 347332 399742 359290 399802
rect 347332 399740 347338 399742
rect 359406 399740 359412 399804
rect 359476 399802 359482 399804
rect 359779 399802 359845 399805
rect 359476 399800 359845 399802
rect 359476 399744 359784 399800
rect 359840 399744 359845 399800
rect 359476 399742 359845 399744
rect 359476 399740 359482 399742
rect 346761 399739 346827 399740
rect 359779 399739 359845 399742
rect 360510 399740 360516 399804
rect 360580 399802 360586 399804
rect 360883 399802 360949 399805
rect 360580 399800 360949 399802
rect 360580 399744 360888 399800
rect 360944 399744 360949 399800
rect 360580 399742 360949 399744
rect 360580 399740 360586 399742
rect 360883 399739 360949 399742
rect 361246 399740 361252 399804
rect 361316 399802 361322 399804
rect 361990 399802 362050 399875
rect 361316 399742 362050 399802
rect 361316 399740 361322 399742
rect 362902 399740 362908 399804
rect 362972 399802 362978 399804
rect 364014 399802 364074 399878
rect 364195 399875 364261 399878
rect 364374 399876 364380 399940
rect 364444 399938 364450 399940
rect 364747 399938 364813 399941
rect 364444 399936 364813 399938
rect 364444 399880 364752 399936
rect 364808 399880 364813 399936
rect 364444 399878 364813 399880
rect 364444 399876 364450 399878
rect 364747 399875 364813 399878
rect 364926 399876 364932 399940
rect 364996 399938 365002 399940
rect 365299 399938 365365 399941
rect 364996 399936 365365 399938
rect 364996 399880 365304 399936
rect 365360 399880 365365 399936
rect 364996 399878 365365 399880
rect 365670 399938 365730 400014
rect 367050 399938 367110 400150
rect 368422 400012 368428 400076
rect 368492 400074 368498 400076
rect 374126 400074 374132 400076
rect 368492 400014 369778 400074
rect 368492 400012 368498 400014
rect 369718 399941 369778 400014
rect 370822 400014 374132 400074
rect 367231 399938 367297 399941
rect 365670 399878 367110 399938
rect 367188 399936 367297 399938
rect 367188 399880 367236 399936
rect 367292 399880 367297 399936
rect 364996 399876 365002 399878
rect 365299 399875 365365 399878
rect 367188 399875 367297 399880
rect 367599 399938 367665 399941
rect 367599 399936 367708 399938
rect 367599 399880 367604 399936
rect 367660 399880 367708 399936
rect 367599 399875 367708 399880
rect 368054 399876 368060 399940
rect 368124 399938 368130 399940
rect 368703 399938 368769 399941
rect 369163 399940 369229 399941
rect 369531 399940 369597 399941
rect 369158 399938 369164 399940
rect 368124 399936 368769 399938
rect 368124 399880 368708 399936
rect 368764 399880 368769 399936
rect 368124 399878 368769 399880
rect 369072 399878 369164 399938
rect 368124 399876 368130 399878
rect 368703 399875 368769 399878
rect 369158 399876 369164 399878
rect 369228 399876 369234 399940
rect 369526 399938 369532 399940
rect 369440 399878 369532 399938
rect 369526 399876 369532 399878
rect 369596 399876 369602 399940
rect 369715 399936 369781 399941
rect 369715 399880 369720 399936
rect 369776 399880 369781 399936
rect 369163 399875 369229 399876
rect 369531 399875 369597 399876
rect 369715 399875 369781 399880
rect 370078 399876 370084 399940
rect 370148 399938 370154 399940
rect 370359 399938 370425 399941
rect 370635 399940 370701 399941
rect 370630 399938 370636 399940
rect 370148 399936 370425 399938
rect 370148 399880 370364 399936
rect 370420 399880 370425 399936
rect 370148 399878 370425 399880
rect 370544 399878 370636 399938
rect 370148 399876 370154 399878
rect 370359 399875 370425 399878
rect 370630 399876 370636 399878
rect 370700 399876 370706 399940
rect 370635 399875 370701 399876
rect 362972 399742 364074 399802
rect 362972 399740 362978 399742
rect 364926 399740 364932 399804
rect 364996 399802 365002 399804
rect 365115 399802 365181 399805
rect 364996 399800 365181 399802
rect 364996 399744 365120 399800
rect 365176 399744 365181 399800
rect 364996 399742 365181 399744
rect 364996 399740 365002 399742
rect 365115 399739 365181 399742
rect 365294 399740 365300 399804
rect 365364 399802 365370 399804
rect 366035 399802 366101 399805
rect 365364 399800 366101 399802
rect 365364 399744 366040 399800
rect 366096 399744 366101 399800
rect 365364 399742 366101 399744
rect 365364 399740 365370 399742
rect 366035 399739 366101 399742
rect 366398 399740 366404 399804
rect 366468 399802 366474 399804
rect 367188 399802 367248 399875
rect 366468 399742 367248 399802
rect 367648 399802 367708 399875
rect 368238 399802 368244 399804
rect 367648 399742 368244 399802
rect 366468 399740 366474 399742
rect 368238 399740 368244 399742
rect 368308 399740 368314 399804
rect 368606 399740 368612 399804
rect 368676 399802 368682 399804
rect 370267 399802 370333 399805
rect 368676 399800 370333 399802
rect 368676 399744 370272 399800
rect 370328 399744 370333 399800
rect 368676 399742 370333 399744
rect 368676 399740 368682 399742
rect 370267 399739 370333 399742
rect 315297 399666 315363 399669
rect 370822 399666 370882 400014
rect 374126 400012 374132 400014
rect 374196 400012 374202 400076
rect 376518 400074 376524 400076
rect 375974 400014 376524 400074
rect 371463 399938 371529 399941
rect 371190 399936 371529 399938
rect 371003 399902 371069 399907
rect 371003 399846 371008 399902
rect 371064 399846 371069 399902
rect 371003 399841 371069 399846
rect 371190 399880 371468 399936
rect 371524 399880 371529 399936
rect 371190 399878 371529 399880
rect 315297 399664 370882 399666
rect 315297 399608 315302 399664
rect 315358 399608 370882 399664
rect 315297 399606 370882 399608
rect 315297 399603 315363 399606
rect 312813 399530 312879 399533
rect 346342 399530 346348 399532
rect 312813 399528 346348 399530
rect 312813 399472 312818 399528
rect 312874 399472 346348 399528
rect 312813 399470 346348 399472
rect 312813 399467 312879 399470
rect 346342 399468 346348 399470
rect 346412 399468 346418 399532
rect 347221 399530 347287 399533
rect 351269 399530 351335 399533
rect 347221 399528 351335 399530
rect 347221 399472 347226 399528
rect 347282 399472 351274 399528
rect 351330 399472 351335 399528
rect 347221 399470 351335 399472
rect 347221 399467 347287 399470
rect 351269 399467 351335 399470
rect 352782 399468 352788 399532
rect 352852 399530 352858 399532
rect 352925 399530 352991 399533
rect 352852 399528 352991 399530
rect 352852 399472 352930 399528
rect 352986 399472 352991 399528
rect 352852 399470 352991 399472
rect 352852 399468 352858 399470
rect 352925 399467 352991 399470
rect 353201 399530 353267 399533
rect 353334 399530 353340 399532
rect 353201 399528 353340 399530
rect 353201 399472 353206 399528
rect 353262 399472 353340 399528
rect 353201 399470 353340 399472
rect 353201 399467 353267 399470
rect 353334 399468 353340 399470
rect 353404 399468 353410 399532
rect 359038 399468 359044 399532
rect 359108 399530 359114 399532
rect 359181 399530 359247 399533
rect 359108 399528 359247 399530
rect 359108 399472 359186 399528
rect 359242 399472 359247 399528
rect 359108 399470 359247 399472
rect 359108 399468 359114 399470
rect 359181 399467 359247 399470
rect 360694 399468 360700 399532
rect 360764 399530 360770 399532
rect 364149 399530 364215 399533
rect 360764 399528 364215 399530
rect 360764 399472 364154 399528
rect 364210 399472 364215 399528
rect 360764 399470 364215 399472
rect 360764 399468 360770 399470
rect 364149 399467 364215 399470
rect 365069 399530 365135 399533
rect 370497 399532 370563 399533
rect 366582 399530 366588 399532
rect 365069 399528 366588 399530
rect 365069 399472 365074 399528
rect 365130 399472 366588 399528
rect 365069 399470 366588 399472
rect 365069 399467 365135 399470
rect 366582 399468 366588 399470
rect 366652 399468 366658 399532
rect 370446 399468 370452 399532
rect 370516 399530 370563 399532
rect 370516 399528 370608 399530
rect 370558 399472 370608 399528
rect 370516 399470 370608 399472
rect 370516 399468 370563 399470
rect 370497 399467 370563 399468
rect 342069 399394 342135 399397
rect 346853 399394 346919 399397
rect 342069 399392 346919 399394
rect 342069 399336 342074 399392
rect 342130 399336 346858 399392
rect 346914 399336 346919 399392
rect 342069 399334 346919 399336
rect 342069 399331 342135 399334
rect 346853 399331 346919 399334
rect 348918 399332 348924 399396
rect 348988 399394 348994 399396
rect 348988 399334 370514 399394
rect 348988 399332 348994 399334
rect 340873 399258 340939 399261
rect 340873 399256 343098 399258
rect 340873 399200 340878 399256
rect 340934 399200 343098 399256
rect 340873 399198 343098 399200
rect 340873 399195 340939 399198
rect 343038 399122 343098 399198
rect 343214 399196 343220 399260
rect 343284 399258 343290 399260
rect 344001 399258 344067 399261
rect 343284 399256 344067 399258
rect 343284 399200 344006 399256
rect 344062 399200 344067 399256
rect 343284 399198 344067 399200
rect 343284 399196 343290 399198
rect 344001 399195 344067 399198
rect 345657 399258 345723 399261
rect 353569 399258 353635 399261
rect 345657 399256 353635 399258
rect 345657 399200 345662 399256
rect 345718 399200 353574 399256
rect 353630 399200 353635 399256
rect 345657 399198 353635 399200
rect 345657 399195 345723 399198
rect 353569 399195 353635 399198
rect 354806 399196 354812 399260
rect 354876 399258 354882 399260
rect 355317 399258 355383 399261
rect 354876 399256 355383 399258
rect 354876 399200 355322 399256
rect 355378 399200 355383 399256
rect 354876 399198 355383 399200
rect 354876 399196 354882 399198
rect 355317 399195 355383 399198
rect 358854 399196 358860 399260
rect 358924 399258 358930 399260
rect 358997 399258 359063 399261
rect 369853 399258 369919 399261
rect 358924 399256 359063 399258
rect 358924 399200 359002 399256
rect 359058 399200 359063 399256
rect 358924 399198 359063 399200
rect 358924 399196 358930 399198
rect 358997 399195 359063 399198
rect 360150 399256 369919 399258
rect 360150 399200 369858 399256
rect 369914 399200 369919 399256
rect 360150 399198 369919 399200
rect 360150 399122 360210 399198
rect 369853 399195 369919 399198
rect 343038 399062 348434 399122
rect 287646 398924 287652 398988
rect 287716 398986 287722 398988
rect 344461 398986 344527 398989
rect 287716 398984 344527 398986
rect 287716 398928 344466 398984
rect 344522 398928 344527 398984
rect 287716 398926 344527 398928
rect 287716 398924 287722 398926
rect 344461 398923 344527 398926
rect 344645 398986 344711 398989
rect 346209 398986 346275 398989
rect 346669 398986 346735 398989
rect 344645 398984 344754 398986
rect 344645 398928 344650 398984
rect 344706 398928 344754 398984
rect 344645 398923 344754 398928
rect 346209 398984 346735 398986
rect 346209 398928 346214 398984
rect 346270 398928 346674 398984
rect 346730 398928 346735 398984
rect 346209 398926 346735 398928
rect 348374 398986 348434 399062
rect 354446 399062 360210 399122
rect 370454 399122 370514 399334
rect 370681 399258 370747 399261
rect 371006 399258 371066 399841
rect 371190 399533 371250 399878
rect 371463 399875 371529 399878
rect 371647 399938 371713 399941
rect 371647 399936 371756 399938
rect 371647 399880 371652 399936
rect 371708 399880 371756 399936
rect 373211 399936 373277 399941
rect 372015 399904 372081 399907
rect 371647 399875 371756 399880
rect 371141 399528 371250 399533
rect 371141 399472 371146 399528
rect 371202 399472 371250 399528
rect 371141 399470 371250 399472
rect 371141 399467 371207 399470
rect 371696 399394 371756 399875
rect 371374 399334 371756 399394
rect 371972 399902 372081 399904
rect 371972 399846 372020 399902
rect 372076 399846 372081 399902
rect 371972 399841 372081 399846
rect 372659 399902 372725 399907
rect 372659 399846 372664 399902
rect 372720 399846 372725 399902
rect 373211 399880 373216 399936
rect 373272 399880 373277 399936
rect 373211 399875 373277 399880
rect 373763 399936 373829 399941
rect 374775 399938 374841 399941
rect 375051 399940 375117 399941
rect 375046 399938 375052 399940
rect 373763 399880 373768 399936
rect 373824 399880 373829 399936
rect 373763 399875 373829 399880
rect 374318 399936 374841 399938
rect 374318 399880 374780 399936
rect 374836 399880 374841 399936
rect 374318 399878 374841 399880
rect 374960 399878 375052 399938
rect 372659 399841 372725 399846
rect 371374 399261 371434 399334
rect 370681 399256 371066 399258
rect 370681 399200 370686 399256
rect 370742 399200 371066 399256
rect 370681 399198 371066 399200
rect 371325 399256 371434 399261
rect 371325 399200 371330 399256
rect 371386 399200 371434 399256
rect 371325 399198 371434 399200
rect 371693 399258 371759 399261
rect 371972 399258 372032 399841
rect 372662 399530 372722 399841
rect 372889 399530 372955 399533
rect 372662 399528 372955 399530
rect 372662 399472 372894 399528
rect 372950 399472 372955 399528
rect 372662 399470 372955 399472
rect 372889 399467 372955 399470
rect 372705 399394 372771 399397
rect 372838 399394 372844 399396
rect 372705 399392 372844 399394
rect 372705 399336 372710 399392
rect 372766 399336 372844 399392
rect 372705 399334 372844 399336
rect 372705 399331 372771 399334
rect 372838 399332 372844 399334
rect 372908 399332 372914 399396
rect 371693 399256 372032 399258
rect 371693 399200 371698 399256
rect 371754 399200 372032 399256
rect 371693 399198 372032 399200
rect 373214 399258 373274 399875
rect 373766 399669 373826 399875
rect 373766 399664 373875 399669
rect 373766 399608 373814 399664
rect 373870 399608 373875 399664
rect 373766 399606 373875 399608
rect 373809 399603 373875 399606
rect 374177 399666 374243 399669
rect 374318 399666 374378 399878
rect 374775 399875 374841 399878
rect 375046 399876 375052 399878
rect 375116 399876 375122 399940
rect 375419 399936 375485 399941
rect 375787 399940 375853 399941
rect 375782 399938 375788 399940
rect 375419 399880 375424 399936
rect 375480 399880 375485 399936
rect 375051 399875 375117 399876
rect 375419 399875 375485 399880
rect 375696 399878 375788 399938
rect 375782 399876 375788 399878
rect 375852 399876 375858 399940
rect 375787 399875 375853 399876
rect 374177 399664 374378 399666
rect 374177 399608 374182 399664
rect 374238 399608 374378 399664
rect 374177 399606 374378 399608
rect 375422 399666 375482 399875
rect 375833 399802 375899 399805
rect 375974 399802 376034 400014
rect 376518 400012 376524 400014
rect 376588 400012 376594 400076
rect 377254 400012 377260 400076
rect 377324 400074 377330 400076
rect 379470 400074 379530 400150
rect 382782 400208 389607 400210
rect 382782 400152 389546 400208
rect 389602 400152 389607 400208
rect 382782 400150 389607 400152
rect 377324 400014 379070 400074
rect 379470 400014 381370 400074
rect 377324 400012 377330 400014
rect 376247 399938 376313 399941
rect 376707 399940 376773 399941
rect 375833 399800 376034 399802
rect 375833 399744 375838 399800
rect 375894 399744 376034 399800
rect 375833 399742 376034 399744
rect 376112 399936 376313 399938
rect 376112 399880 376252 399936
rect 376308 399880 376313 399936
rect 376112 399878 376313 399880
rect 375833 399739 375899 399742
rect 375557 399666 375623 399669
rect 375422 399664 375623 399666
rect 375422 399608 375562 399664
rect 375618 399608 375623 399664
rect 375422 399606 375623 399608
rect 376112 399666 376172 399878
rect 376247 399875 376313 399878
rect 376523 399902 376589 399907
rect 376523 399846 376528 399902
rect 376584 399846 376589 399902
rect 376702 399876 376708 399940
rect 376772 399938 376778 399940
rect 376983 399938 377049 399941
rect 378179 399938 378245 399941
rect 378731 399940 378797 399941
rect 378726 399938 378732 399940
rect 376772 399878 376864 399938
rect 376983 399936 377184 399938
rect 376983 399880 376988 399936
rect 377044 399880 377184 399936
rect 378136 399936 378245 399938
rect 376983 399878 377184 399880
rect 376772 399876 376778 399878
rect 376707 399875 376773 399876
rect 376983 399875 377049 399878
rect 376523 399841 376589 399846
rect 376526 399669 376586 399841
rect 377124 399669 377184 399878
rect 377995 399902 378061 399907
rect 377995 399846 378000 399902
rect 378056 399846 378061 399902
rect 377995 399841 378061 399846
rect 378136 399880 378184 399936
rect 378240 399880 378245 399936
rect 378136 399875 378245 399880
rect 378640 399878 378732 399938
rect 378726 399876 378732 399878
rect 378796 399876 378802 399940
rect 379010 399938 379070 400014
rect 379467 399938 379533 399941
rect 379743 399938 379809 399941
rect 379010 399936 379533 399938
rect 379010 399880 379472 399936
rect 379528 399880 379533 399936
rect 379010 399878 379533 399880
rect 378731 399875 378797 399876
rect 379467 399875 379533 399878
rect 379700 399936 379809 399938
rect 379700 399880 379748 399936
rect 379804 399880 379809 399936
rect 379700 399875 379809 399880
rect 379927 399938 379993 399941
rect 380198 399938 380204 399940
rect 379927 399936 380204 399938
rect 379927 399880 379932 399936
rect 379988 399880 380204 399936
rect 379927 399878 380204 399880
rect 379927 399875 379993 399878
rect 380198 399876 380204 399878
rect 380268 399876 380274 399940
rect 380571 399936 380637 399941
rect 380387 399902 380453 399907
rect 376293 399666 376359 399669
rect 376112 399664 376359 399666
rect 376112 399608 376298 399664
rect 376354 399608 376359 399664
rect 376112 399606 376359 399608
rect 376526 399664 376635 399669
rect 376526 399608 376574 399664
rect 376630 399608 376635 399664
rect 376526 399606 376635 399608
rect 374177 399603 374243 399606
rect 375557 399603 375623 399606
rect 376293 399603 376359 399606
rect 376569 399603 376635 399606
rect 377121 399664 377187 399669
rect 377121 399608 377126 399664
rect 377182 399608 377187 399664
rect 377121 399603 377187 399608
rect 374637 399530 374703 399533
rect 375281 399530 375347 399533
rect 377489 399530 377555 399533
rect 374637 399528 374746 399530
rect 374637 399472 374642 399528
rect 374698 399472 374746 399528
rect 374637 399467 374746 399472
rect 375281 399528 377555 399530
rect 375281 399472 375286 399528
rect 375342 399472 377494 399528
rect 377550 399472 377555 399528
rect 375281 399470 377555 399472
rect 375281 399467 375347 399470
rect 377489 399467 377555 399470
rect 373625 399258 373691 399261
rect 373214 399256 373691 399258
rect 373214 399200 373630 399256
rect 373686 399200 373691 399256
rect 373214 399198 373691 399200
rect 370681 399195 370747 399198
rect 371325 399195 371391 399198
rect 371693 399195 371759 399198
rect 373625 399195 373691 399198
rect 372654 399122 372660 399124
rect 370454 399062 372660 399122
rect 353385 398986 353451 398989
rect 348374 398984 353451 398986
rect 348374 398928 353390 398984
rect 353446 398928 353451 398984
rect 348374 398926 353451 398928
rect 346209 398923 346275 398926
rect 346669 398923 346735 398926
rect 353385 398923 353451 398926
rect 353886 398924 353892 398988
rect 353956 398986 353962 398988
rect 354446 398986 354506 399062
rect 372654 399060 372660 399062
rect 372724 399060 372730 399124
rect 374686 399122 374746 399467
rect 376886 399332 376892 399396
rect 376956 399394 376962 399396
rect 377998 399394 378058 399841
rect 378136 399805 378196 399875
rect 378133 399800 378199 399805
rect 378133 399744 378138 399800
rect 378194 399744 378199 399800
rect 378133 399739 378199 399744
rect 378455 399802 378521 399805
rect 378910 399802 378916 399804
rect 378455 399800 378916 399802
rect 378455 399744 378460 399800
rect 378516 399744 378916 399800
rect 378455 399742 378916 399744
rect 378455 399739 378521 399742
rect 378910 399740 378916 399742
rect 378980 399740 378986 399804
rect 378225 399666 378291 399669
rect 379700 399666 379760 399875
rect 380387 399846 380392 399902
rect 380448 399846 380453 399902
rect 380571 399880 380576 399936
rect 380632 399880 380637 399936
rect 380571 399875 380637 399880
rect 380847 399936 380913 399941
rect 380847 399880 380852 399936
rect 380908 399880 380913 399936
rect 380847 399875 380913 399880
rect 381031 399940 381097 399941
rect 381031 399936 381078 399940
rect 381142 399938 381148 399940
rect 381031 399880 381036 399936
rect 381031 399876 381078 399880
rect 381142 399878 381188 399938
rect 381142 399876 381148 399878
rect 381031 399875 381097 399876
rect 380387 399841 380453 399846
rect 378225 399664 379760 399666
rect 378225 399608 378230 399664
rect 378286 399608 379760 399664
rect 380203 399698 380269 399703
rect 380203 399642 380208 399698
rect 380264 399642 380269 399698
rect 380390 399669 380450 399841
rect 380203 399637 380269 399642
rect 380341 399664 380450 399669
rect 378225 399606 379760 399608
rect 378225 399603 378291 399606
rect 376956 399334 378058 399394
rect 376956 399332 376962 399334
rect 378174 399196 378180 399260
rect 378244 399258 378250 399260
rect 378593 399258 378659 399261
rect 378244 399256 378659 399258
rect 378244 399200 378598 399256
rect 378654 399200 378659 399256
rect 378244 399198 378659 399200
rect 378244 399196 378250 399198
rect 378593 399195 378659 399198
rect 379646 399196 379652 399260
rect 379716 399258 379722 399260
rect 380206 399258 380266 399637
rect 380341 399608 380346 399664
rect 380402 399608 380450 399664
rect 380341 399606 380450 399608
rect 380574 399669 380634 399875
rect 380850 399805 380910 399875
rect 380801 399800 380910 399805
rect 380801 399744 380806 399800
rect 380862 399744 380910 399800
rect 380801 399742 380910 399744
rect 381123 399800 381189 399805
rect 381123 399744 381128 399800
rect 381184 399744 381189 399800
rect 380801 399739 380867 399742
rect 381123 399739 381189 399744
rect 381310 399802 381370 400014
rect 382782 399941 382842 400150
rect 389541 400147 389607 400150
rect 384982 400012 384988 400076
rect 385052 400074 385058 400076
rect 390645 400074 390711 400077
rect 385052 400014 386338 400074
rect 385052 400012 385058 400014
rect 386278 399941 386338 400014
rect 386646 400072 390711 400074
rect 386646 400016 390650 400072
rect 390706 400016 390711 400072
rect 386646 400014 390711 400016
rect 386646 399941 386706 400014
rect 390645 400011 390711 400014
rect 381486 399876 381492 399940
rect 381556 399938 381562 399940
rect 382319 399938 382385 399941
rect 381556 399936 382385 399938
rect 381556 399880 382324 399936
rect 382380 399880 382385 399936
rect 381556 399878 382385 399880
rect 381556 399876 381562 399878
rect 382319 399875 382385 399878
rect 382779 399936 382845 399941
rect 382779 399880 382784 399936
rect 382840 399880 382845 399936
rect 383147 399936 383213 399941
rect 383791 399938 383857 399941
rect 382779 399875 382845 399880
rect 382963 399902 383029 399907
rect 382963 399846 382968 399902
rect 383024 399846 383029 399902
rect 383147 399880 383152 399936
rect 383208 399880 383213 399936
rect 383147 399875 383213 399880
rect 383610 399936 383857 399938
rect 383610 399880 383796 399936
rect 383852 399880 383857 399936
rect 385355 399936 385421 399941
rect 385815 399938 385881 399941
rect 383610 399878 383857 399880
rect 382963 399841 383029 399846
rect 382222 399802 382228 399804
rect 381310 399742 382228 399802
rect 382222 399740 382228 399742
rect 382292 399740 382298 399804
rect 380574 399664 380683 399669
rect 380574 399608 380622 399664
rect 380678 399608 380683 399664
rect 380574 399606 380683 399608
rect 380341 399603 380407 399606
rect 380617 399603 380683 399606
rect 379716 399198 380266 399258
rect 381126 399258 381186 399739
rect 381261 399668 381327 399669
rect 381261 399664 381308 399668
rect 381372 399666 381378 399668
rect 381261 399608 381266 399664
rect 381261 399604 381308 399608
rect 381372 399606 381418 399666
rect 381372 399604 381378 399606
rect 381670 399604 381676 399668
rect 381740 399666 381746 399668
rect 382966 399666 383026 399841
rect 383150 399805 383210 399875
rect 383150 399800 383259 399805
rect 383150 399744 383198 399800
rect 383254 399744 383259 399800
rect 383150 399742 383259 399744
rect 383610 399802 383670 399878
rect 383791 399875 383857 399878
rect 384067 399902 384133 399907
rect 384067 399846 384072 399902
rect 384128 399846 384133 399902
rect 384067 399841 384133 399846
rect 384435 399902 384501 399907
rect 384435 399846 384440 399902
rect 384496 399846 384501 399902
rect 384435 399841 384501 399846
rect 384987 399902 385053 399907
rect 384987 399846 384992 399902
rect 385048 399846 385053 399902
rect 385355 399880 385360 399936
rect 385416 399880 385421 399936
rect 385355 399875 385421 399880
rect 385542 399936 385881 399938
rect 385542 399880 385820 399936
rect 385876 399880 385881 399936
rect 385542 399878 385881 399880
rect 384987 399841 385053 399846
rect 383745 399802 383811 399805
rect 383610 399800 383811 399802
rect 383610 399744 383750 399800
rect 383806 399744 383811 399800
rect 383610 399742 383811 399744
rect 383193 399739 383259 399742
rect 383745 399739 383811 399742
rect 381740 399606 383026 399666
rect 381740 399604 381746 399606
rect 381261 399603 381327 399604
rect 381629 399258 381695 399261
rect 384070 399258 384130 399841
rect 384438 399394 384498 399841
rect 381126 399256 381695 399258
rect 381126 399200 381634 399256
rect 381690 399200 381695 399256
rect 381126 399198 381695 399200
rect 379716 399196 379722 399198
rect 381629 399195 381695 399198
rect 383886 399198 384130 399258
rect 384254 399334 384498 399394
rect 374913 399122 374979 399125
rect 374686 399120 374979 399122
rect 374686 399064 374918 399120
rect 374974 399064 374979 399120
rect 374686 399062 374979 399064
rect 374913 399059 374979 399062
rect 353956 398926 354506 398986
rect 353956 398924 353962 398926
rect 359038 398924 359044 398988
rect 359108 398986 359114 398988
rect 360326 398986 360332 398988
rect 359108 398926 360332 398986
rect 359108 398924 359114 398926
rect 360326 398924 360332 398926
rect 360396 398924 360402 398988
rect 383886 398986 383946 399198
rect 384113 399122 384179 399125
rect 384254 399122 384314 399334
rect 384430 399196 384436 399260
rect 384500 399258 384506 399260
rect 384849 399258 384915 399261
rect 384500 399256 384915 399258
rect 384500 399200 384854 399256
rect 384910 399200 384915 399256
rect 384500 399198 384915 399200
rect 384990 399258 385050 399841
rect 385217 399530 385283 399533
rect 385358 399530 385418 399875
rect 385542 399533 385602 399878
rect 385815 399875 385881 399878
rect 386275 399936 386341 399941
rect 386275 399880 386280 399936
rect 386336 399880 386341 399936
rect 386275 399875 386341 399880
rect 386643 399936 386709 399941
rect 386643 399880 386648 399936
rect 386704 399880 386709 399936
rect 386643 399875 386709 399880
rect 386827 399936 386893 399941
rect 387103 399938 387169 399941
rect 386827 399880 386832 399936
rect 386888 399880 386893 399936
rect 386827 399875 386893 399880
rect 387060 399936 387169 399938
rect 387060 399880 387108 399936
rect 387164 399880 387169 399936
rect 387060 399875 387169 399880
rect 385718 399604 385724 399668
rect 385788 399666 385794 399668
rect 386137 399666 386203 399669
rect 385788 399664 386203 399666
rect 385788 399608 386142 399664
rect 386198 399608 386203 399664
rect 385788 399606 386203 399608
rect 385788 399604 385794 399606
rect 386137 399603 386203 399606
rect 386505 399666 386571 399669
rect 386830 399666 386890 399875
rect 386505 399664 386890 399666
rect 386505 399608 386510 399664
rect 386566 399608 386890 399664
rect 386505 399606 386890 399608
rect 386505 399603 386571 399606
rect 385217 399528 385418 399530
rect 385217 399472 385222 399528
rect 385278 399472 385418 399528
rect 385217 399470 385418 399472
rect 385493 399528 385602 399533
rect 385493 399472 385498 399528
rect 385554 399472 385602 399528
rect 385493 399470 385602 399472
rect 386873 399530 386939 399533
rect 387060 399530 387120 399875
rect 386873 399528 387120 399530
rect 386873 399472 386878 399528
rect 386934 399472 387120 399528
rect 386873 399470 387120 399472
rect 385217 399467 385283 399470
rect 385493 399467 385559 399470
rect 386873 399467 386939 399470
rect 384990 399198 385970 399258
rect 384500 399196 384506 399198
rect 384849 399195 384915 399198
rect 384113 399120 384314 399122
rect 384113 399064 384118 399120
rect 384174 399064 384314 399120
rect 384113 399062 384314 399064
rect 384113 399059 384179 399062
rect 384941 398986 385007 398989
rect 383886 398984 385007 398986
rect 383886 398928 384946 398984
rect 385002 398928 385007 398984
rect 383886 398926 385007 398928
rect 384941 398923 385007 398926
rect 293166 398788 293172 398852
rect 293236 398850 293242 398852
rect 340873 398850 340939 398853
rect 293236 398848 340939 398850
rect 293236 398792 340878 398848
rect 340934 398792 340939 398848
rect 293236 398790 340939 398792
rect 293236 398788 293242 398790
rect 340873 398787 340939 398790
rect 341057 398850 341123 398853
rect 344694 398850 344754 398923
rect 385910 398853 385970 399198
rect 341057 398848 344754 398850
rect 341057 398792 341062 398848
rect 341118 398792 344754 398848
rect 341057 398790 344754 398792
rect 341057 398787 341123 398790
rect 346342 398788 346348 398852
rect 346412 398850 346418 398852
rect 348918 398850 348924 398852
rect 346412 398790 348924 398850
rect 346412 398788 346418 398790
rect 348918 398788 348924 398790
rect 348988 398788 348994 398852
rect 349153 398850 349219 398853
rect 355685 398850 355751 398853
rect 349153 398848 355751 398850
rect 349153 398792 349158 398848
rect 349214 398792 355690 398848
rect 355746 398792 355751 398848
rect 349153 398790 355751 398792
rect 349153 398787 349219 398790
rect 355685 398787 355751 398790
rect 360326 398788 360332 398852
rect 360396 398850 360402 398852
rect 361481 398850 361547 398853
rect 372521 398850 372587 398853
rect 360396 398848 361547 398850
rect 360396 398792 361486 398848
rect 361542 398792 361547 398848
rect 360396 398790 361547 398792
rect 360396 398788 360402 398790
rect 361481 398787 361547 398790
rect 372478 398848 372587 398850
rect 372478 398792 372526 398848
rect 372582 398792 372587 398848
rect 372478 398787 372587 398792
rect 374453 398852 374519 398853
rect 374453 398848 374500 398852
rect 374564 398850 374570 398852
rect 374453 398792 374458 398848
rect 374453 398788 374500 398792
rect 374564 398790 374610 398850
rect 385861 398848 385970 398853
rect 385861 398792 385866 398848
rect 385922 398792 385970 398848
rect 385861 398790 385970 398792
rect 374564 398788 374570 398790
rect 374453 398787 374519 398788
rect 385861 398787 385927 398790
rect 347405 398714 347471 398717
rect 340830 398712 347471 398714
rect 340830 398656 347410 398712
rect 347466 398656 347471 398712
rect 340830 398654 347471 398656
rect 340830 398578 340890 398654
rect 347405 398651 347471 398654
rect 366541 398716 366607 398717
rect 370037 398716 370103 398717
rect 366541 398712 366588 398716
rect 366652 398714 366658 398716
rect 370037 398714 370084 398716
rect 366541 398656 366546 398712
rect 366541 398652 366588 398656
rect 366652 398654 366698 398714
rect 369992 398712 370084 398714
rect 369992 398656 370042 398712
rect 369992 398654 370084 398656
rect 366652 398652 366658 398654
rect 370037 398652 370084 398654
rect 370148 398652 370154 398716
rect 372245 398714 372311 398717
rect 372478 398714 372538 398787
rect 372245 398712 372538 398714
rect 372245 398656 372250 398712
rect 372306 398656 372538 398712
rect 372245 398654 372538 398656
rect 366541 398651 366607 398652
rect 370037 398651 370103 398652
rect 372245 398651 372311 398654
rect 380750 398652 380756 398716
rect 380820 398714 380826 398716
rect 381486 398714 381492 398716
rect 380820 398654 381492 398714
rect 380820 398652 380826 398654
rect 381486 398652 381492 398654
rect 381556 398652 381562 398716
rect 335310 398518 340890 398578
rect 330477 398442 330543 398445
rect 335310 398442 335370 398518
rect 346526 398516 346532 398580
rect 346596 398578 346602 398580
rect 351310 398578 351316 398580
rect 346596 398518 351316 398578
rect 346596 398516 346602 398518
rect 351310 398516 351316 398518
rect 351380 398516 351386 398580
rect 364742 398516 364748 398580
rect 364812 398578 364818 398580
rect 368657 398578 368723 398581
rect 364812 398576 368723 398578
rect 364812 398520 368662 398576
rect 368718 398520 368723 398576
rect 364812 398518 368723 398520
rect 364812 398516 364818 398518
rect 368657 398515 368723 398518
rect 370078 398516 370084 398580
rect 370148 398578 370154 398580
rect 370589 398578 370655 398581
rect 370148 398576 370655 398578
rect 370148 398520 370594 398576
rect 370650 398520 370655 398576
rect 370148 398518 370655 398520
rect 370148 398516 370154 398518
rect 370589 398515 370655 398518
rect 330477 398440 335370 398442
rect 330477 398384 330482 398440
rect 330538 398384 335370 398440
rect 330477 398382 335370 398384
rect 330477 398379 330543 398382
rect 349286 398380 349292 398444
rect 349356 398442 349362 398444
rect 349981 398442 350047 398445
rect 349356 398440 350047 398442
rect 349356 398384 349986 398440
rect 350042 398384 350047 398440
rect 349356 398382 350047 398384
rect 349356 398380 349362 398382
rect 349981 398379 350047 398382
rect 352046 398380 352052 398444
rect 352116 398442 352122 398444
rect 352281 398442 352347 398445
rect 370221 398442 370287 398445
rect 370589 398444 370655 398445
rect 370589 398442 370636 398444
rect 352116 398440 352347 398442
rect 352116 398384 352286 398440
rect 352342 398384 352347 398440
rect 352116 398382 352347 398384
rect 352116 398380 352122 398382
rect 352281 398379 352347 398382
rect 364566 398440 370287 398442
rect 364566 398384 370226 398440
rect 370282 398384 370287 398440
rect 364566 398382 370287 398384
rect 370544 398440 370636 398442
rect 370544 398384 370594 398440
rect 370544 398382 370636 398384
rect 302969 398306 303035 398309
rect 341057 398306 341123 398309
rect 302969 398304 341123 398306
rect 302969 398248 302974 398304
rect 303030 398248 341062 398304
rect 341118 398248 341123 398304
rect 302969 398246 341123 398248
rect 302969 398243 303035 398246
rect 341057 398243 341123 398246
rect 341425 398306 341491 398309
rect 349981 398306 350047 398309
rect 356830 398306 356836 398308
rect 341425 398304 350047 398306
rect 341425 398248 341430 398304
rect 341486 398248 349986 398304
rect 350042 398248 350047 398304
rect 341425 398246 350047 398248
rect 341425 398243 341491 398246
rect 349981 398243 350047 398246
rect 356654 398246 356836 398306
rect 356654 398173 356714 398246
rect 356830 398244 356836 398246
rect 356900 398244 356906 398308
rect 295333 398170 295399 398173
rect 342805 398170 342871 398173
rect 347865 398170 347931 398173
rect 295333 398168 342871 398170
rect 295333 398112 295338 398168
rect 295394 398112 342810 398168
rect 342866 398112 342871 398168
rect 295333 398110 342871 398112
rect 295333 398107 295399 398110
rect 342805 398107 342871 398110
rect 344464 398168 347931 398170
rect 344464 398112 347870 398168
rect 347926 398112 347931 398168
rect 344464 398110 347931 398112
rect 356654 398168 356763 398173
rect 356654 398112 356702 398168
rect 356758 398112 356763 398168
rect 356654 398110 356763 398112
rect 270309 398034 270375 398037
rect 344464 398034 344524 398110
rect 347865 398107 347931 398110
rect 356697 398107 356763 398110
rect 356830 398108 356836 398172
rect 356900 398170 356906 398172
rect 356900 398110 363338 398170
rect 356900 398108 356906 398110
rect 270309 398032 344524 398034
rect 270309 397976 270314 398032
rect 270370 397976 344524 398032
rect 270309 397974 344524 397976
rect 270309 397971 270375 397974
rect 345238 397972 345244 398036
rect 345308 398034 345314 398036
rect 345841 398034 345907 398037
rect 345308 398032 345907 398034
rect 345308 397976 345846 398032
rect 345902 397976 345907 398032
rect 345308 397974 345907 397976
rect 345308 397972 345314 397974
rect 345841 397971 345907 397974
rect 350758 397972 350764 398036
rect 350828 398034 350834 398036
rect 351821 398034 351887 398037
rect 350828 398032 351887 398034
rect 350828 397976 351826 398032
rect 351882 397976 351887 398032
rect 350828 397974 351887 397976
rect 350828 397972 350834 397974
rect 351821 397971 351887 397974
rect 355358 397972 355364 398036
rect 355428 398034 355434 398036
rect 355428 397974 357450 398034
rect 355428 397972 355434 397974
rect 339217 397898 339283 397901
rect 349797 397898 349863 397901
rect 339217 397896 345674 397898
rect 339217 397840 339222 397896
rect 339278 397840 345674 397896
rect 339217 397838 345674 397840
rect 339217 397835 339283 397838
rect -960 397490 480 397580
rect 3417 397490 3483 397493
rect -960 397488 3483 397490
rect -960 397432 3422 397488
rect 3478 397432 3483 397488
rect -960 397430 3483 397432
rect 345614 397490 345674 397838
rect 347270 397896 349863 397898
rect 347270 397840 349802 397896
rect 349858 397840 349863 397896
rect 347270 397838 349863 397840
rect 347270 397765 347330 397838
rect 349797 397835 349863 397838
rect 350574 397836 350580 397900
rect 350644 397898 350650 397900
rect 351085 397898 351151 397901
rect 350644 397896 351151 397898
rect 350644 397840 351090 397896
rect 351146 397840 351151 397896
rect 350644 397838 351151 397840
rect 357390 397898 357450 397974
rect 362718 397972 362724 398036
rect 362788 398034 362794 398036
rect 362861 398034 362927 398037
rect 362788 398032 362927 398034
rect 362788 397976 362866 398032
rect 362922 397976 362927 398032
rect 362788 397974 362927 397976
rect 363278 398034 363338 398110
rect 363454 398108 363460 398172
rect 363524 398170 363530 398172
rect 364566 398170 364626 398382
rect 370221 398379 370287 398382
rect 370589 398380 370636 398382
rect 370700 398380 370706 398444
rect 376702 398380 376708 398444
rect 376772 398442 376778 398444
rect 380801 398442 380867 398445
rect 376772 398440 380867 398442
rect 376772 398384 380806 398440
rect 380862 398384 380867 398440
rect 376772 398382 380867 398384
rect 376772 398380 376778 398382
rect 370589 398379 370655 398380
rect 380801 398379 380867 398382
rect 383694 398380 383700 398444
rect 383764 398442 383770 398444
rect 384573 398442 384639 398445
rect 383764 398440 384639 398442
rect 383764 398384 384578 398440
rect 384634 398384 384639 398440
rect 383764 398382 384639 398384
rect 383764 398380 383770 398382
rect 384573 398379 384639 398382
rect 372654 398244 372660 398308
rect 372724 398306 372730 398308
rect 373349 398306 373415 398309
rect 372724 398304 373415 398306
rect 372724 398248 373354 398304
rect 373410 398248 373415 398304
rect 372724 398246 373415 398248
rect 372724 398244 372730 398246
rect 373349 398243 373415 398246
rect 383285 398306 383351 398309
rect 388253 398306 388319 398309
rect 383285 398304 388319 398306
rect 383285 398248 383290 398304
rect 383346 398248 388258 398304
rect 388314 398248 388319 398304
rect 383285 398246 388319 398248
rect 383285 398243 383351 398246
rect 388253 398243 388319 398246
rect 363524 398110 364626 398170
rect 363524 398108 363530 398110
rect 367318 398108 367324 398172
rect 367388 398170 367394 398172
rect 367461 398170 367527 398173
rect 367388 398168 367527 398170
rect 367388 398112 367466 398168
rect 367522 398112 367527 398168
rect 367388 398110 367527 398112
rect 367388 398108 367394 398110
rect 367461 398107 367527 398110
rect 367686 398108 367692 398172
rect 367756 398170 367762 398172
rect 372981 398170 373047 398173
rect 367756 398168 373047 398170
rect 367756 398112 372986 398168
rect 373042 398112 373047 398168
rect 367756 398110 373047 398112
rect 367756 398108 367762 398110
rect 372981 398107 373047 398110
rect 382089 398170 382155 398173
rect 384665 398170 384731 398173
rect 382089 398168 384731 398170
rect 382089 398112 382094 398168
rect 382150 398112 384670 398168
rect 384726 398112 384731 398168
rect 382089 398110 384731 398112
rect 382089 398107 382155 398110
rect 384665 398107 384731 398110
rect 367829 398034 367895 398037
rect 368289 398036 368355 398037
rect 363278 398032 367895 398034
rect 363278 397976 367834 398032
rect 367890 397976 367895 398032
rect 363278 397974 367895 397976
rect 362788 397972 362794 397974
rect 362861 397971 362927 397974
rect 367829 397971 367895 397974
rect 368238 397972 368244 398036
rect 368308 398034 368355 398036
rect 368308 398032 368400 398034
rect 368350 397976 368400 398032
rect 368308 397974 368400 397976
rect 368308 397972 368355 397974
rect 368974 397972 368980 398036
rect 369044 398034 369050 398036
rect 374269 398034 374335 398037
rect 369044 398032 374335 398034
rect 369044 397976 374274 398032
rect 374330 397976 374335 398032
rect 369044 397974 374335 397976
rect 369044 397972 369050 397974
rect 368289 397971 368355 397972
rect 374269 397971 374335 397974
rect 379513 398034 379579 398037
rect 382641 398034 382707 398037
rect 379513 398032 382707 398034
rect 379513 397976 379518 398032
rect 379574 397976 382646 398032
rect 382702 397976 382707 398032
rect 379513 397974 382707 397976
rect 379513 397971 379579 397974
rect 382641 397971 382707 397974
rect 384021 398034 384087 398037
rect 392117 398034 392183 398037
rect 384021 398032 392183 398034
rect 384021 397976 384026 398032
rect 384082 397976 392122 398032
rect 392178 397976 392183 398032
rect 384021 397974 392183 397976
rect 384021 397971 384087 397974
rect 392117 397971 392183 397974
rect 365294 397898 365300 397900
rect 357390 397838 365300 397898
rect 350644 397836 350650 397838
rect 351085 397835 351151 397838
rect 365294 397836 365300 397838
rect 365364 397836 365370 397900
rect 368749 397898 368815 397901
rect 369526 397898 369532 397900
rect 368749 397896 369532 397898
rect 368749 397840 368754 397896
rect 368810 397840 369532 397896
rect 368749 397838 369532 397840
rect 368749 397835 368815 397838
rect 369526 397836 369532 397838
rect 369596 397836 369602 397900
rect 369894 397836 369900 397900
rect 369964 397898 369970 397900
rect 371049 397898 371115 397901
rect 369964 397896 371115 397898
rect 369964 397840 371054 397896
rect 371110 397840 371115 397896
rect 369964 397838 371115 397840
rect 369964 397836 369970 397838
rect 371049 397835 371115 397838
rect 372705 397898 372771 397901
rect 372838 397898 372844 397900
rect 372705 397896 372844 397898
rect 372705 397840 372710 397896
rect 372766 397840 372844 397896
rect 372705 397838 372844 397840
rect 372705 397835 372771 397838
rect 372838 397836 372844 397838
rect 372908 397836 372914 397900
rect 382774 397836 382780 397900
rect 382844 397898 382850 397900
rect 386045 397898 386111 397901
rect 382844 397896 386111 397898
rect 382844 397840 386050 397896
rect 386106 397840 386111 397896
rect 382844 397838 386111 397840
rect 382844 397836 382850 397838
rect 386045 397835 386111 397838
rect 347221 397760 347330 397765
rect 361481 397762 361547 397765
rect 347221 397704 347226 397760
rect 347282 397704 347330 397760
rect 347221 397702 347330 397704
rect 350582 397760 361547 397762
rect 350582 397704 361486 397760
rect 361542 397704 361547 397760
rect 350582 397702 361547 397704
rect 347221 397699 347287 397702
rect 347998 397564 348004 397628
rect 348068 397626 348074 397628
rect 348601 397626 348667 397629
rect 348068 397624 348667 397626
rect 348068 397568 348606 397624
rect 348662 397568 348667 397624
rect 348068 397566 348667 397568
rect 348068 397564 348074 397566
rect 348601 397563 348667 397566
rect 349981 397626 350047 397629
rect 350582 397626 350642 397702
rect 361481 397699 361547 397702
rect 370262 397700 370268 397764
rect 370332 397762 370338 397764
rect 370773 397762 370839 397765
rect 370332 397760 370839 397762
rect 370332 397704 370778 397760
rect 370834 397704 370839 397760
rect 370332 397702 370839 397704
rect 370332 397700 370338 397702
rect 370773 397699 370839 397702
rect 358813 397626 358879 397629
rect 349981 397624 350642 397626
rect 349981 397568 349986 397624
rect 350042 397568 350642 397624
rect 349981 397566 350642 397568
rect 350766 397624 358879 397626
rect 350766 397568 358818 397624
rect 358874 397568 358879 397624
rect 350766 397566 358879 397568
rect 349981 397563 350047 397566
rect 350766 397490 350826 397566
rect 358813 397563 358879 397566
rect 369158 397564 369164 397628
rect 369228 397626 369234 397628
rect 373073 397626 373139 397629
rect 369228 397624 373139 397626
rect 369228 397568 373078 397624
rect 373134 397568 373139 397624
rect 369228 397566 373139 397568
rect 369228 397564 369234 397566
rect 373073 397563 373139 397566
rect 376753 397626 376819 397629
rect 382089 397626 382155 397629
rect 376753 397624 382155 397626
rect 376753 397568 376758 397624
rect 376814 397568 382094 397624
rect 382150 397568 382155 397624
rect 376753 397566 382155 397568
rect 376753 397563 376819 397566
rect 382089 397563 382155 397566
rect 382222 397564 382228 397628
rect 382292 397626 382298 397628
rect 383469 397626 383535 397629
rect 382292 397624 383535 397626
rect 382292 397568 383474 397624
rect 383530 397568 383535 397624
rect 382292 397566 383535 397568
rect 382292 397564 382298 397566
rect 383469 397563 383535 397566
rect 345614 397430 350826 397490
rect -960 397340 480 397430
rect 3417 397427 3483 397430
rect 351862 397428 351868 397492
rect 351932 397490 351938 397492
rect 353017 397490 353083 397493
rect 353293 397492 353359 397493
rect 353293 397490 353340 397492
rect 351932 397488 353083 397490
rect 351932 397432 353022 397488
rect 353078 397432 353083 397488
rect 351932 397430 353083 397432
rect 353248 397488 353340 397490
rect 353248 397432 353298 397488
rect 353248 397430 353340 397432
rect 351932 397428 351938 397430
rect 353017 397427 353083 397430
rect 353293 397428 353340 397430
rect 353404 397428 353410 397492
rect 357382 397428 357388 397492
rect 357452 397490 357458 397492
rect 357985 397490 358051 397493
rect 357452 397488 358051 397490
rect 357452 397432 357990 397488
rect 358046 397432 358051 397488
rect 357452 397430 358051 397432
rect 357452 397428 357458 397430
rect 353293 397427 353359 397428
rect 357985 397427 358051 397430
rect 371366 397428 371372 397492
rect 371436 397490 371442 397492
rect 372429 397490 372495 397493
rect 371436 397488 372495 397490
rect 371436 397432 372434 397488
rect 372490 397432 372495 397488
rect 371436 397430 372495 397432
rect 371436 397428 371442 397430
rect 372429 397427 372495 397430
rect 373206 397428 373212 397492
rect 373276 397490 373282 397492
rect 374821 397490 374887 397493
rect 373276 397488 374887 397490
rect 373276 397432 374826 397488
rect 374882 397432 374887 397488
rect 373276 397430 374887 397432
rect 373276 397428 373282 397430
rect 374821 397427 374887 397430
rect 378358 397428 378364 397492
rect 378428 397490 378434 397492
rect 379145 397490 379211 397493
rect 378428 397488 379211 397490
rect 378428 397432 379150 397488
rect 379206 397432 379211 397488
rect 378428 397430 379211 397432
rect 378428 397428 378434 397430
rect 379145 397427 379211 397430
rect 380934 397428 380940 397492
rect 381004 397490 381010 397492
rect 382181 397490 382247 397493
rect 381004 397488 382247 397490
rect 381004 397432 382186 397488
rect 382242 397432 382247 397488
rect 381004 397430 382247 397432
rect 381004 397428 381010 397430
rect 382181 397427 382247 397430
rect 331949 397354 332015 397357
rect 348325 397354 348391 397357
rect 331949 397352 348391 397354
rect 331949 397296 331954 397352
rect 332010 397296 348330 397352
rect 348386 397296 348391 397352
rect 331949 397294 348391 397296
rect 331949 397291 332015 397294
rect 348325 397291 348391 397294
rect 363638 397292 363644 397356
rect 363708 397354 363714 397356
rect 366357 397354 366423 397357
rect 366633 397356 366699 397357
rect 367185 397356 367251 397357
rect 366582 397354 366588 397356
rect 363708 397352 366423 397354
rect 363708 397296 366362 397352
rect 366418 397296 366423 397352
rect 363708 397294 366423 397296
rect 366542 397294 366588 397354
rect 366652 397352 366699 397356
rect 367134 397354 367140 397356
rect 366694 397296 366699 397352
rect 363708 397292 363714 397294
rect 366357 397291 366423 397294
rect 366582 397292 366588 397294
rect 366652 397292 366699 397296
rect 367094 397294 367140 397354
rect 367204 397352 367251 397356
rect 367246 397296 367251 397352
rect 367134 397292 367140 397294
rect 367204 397292 367251 397296
rect 366633 397291 366699 397292
rect 367185 397291 367251 397292
rect 330753 397218 330819 397221
rect 355961 397218 356027 397221
rect 330753 397216 356027 397218
rect 330753 397160 330758 397216
rect 330814 397160 355966 397216
rect 356022 397160 356027 397216
rect 330753 397158 356027 397160
rect 330753 397155 330819 397158
rect 355961 397155 356027 397158
rect 356646 397156 356652 397220
rect 356716 397218 356722 397220
rect 364742 397218 364748 397220
rect 356716 397158 364748 397218
rect 356716 397156 356722 397158
rect 364742 397156 364748 397158
rect 364812 397156 364818 397220
rect 318558 397020 318564 397084
rect 318628 397082 318634 397084
rect 378041 397082 378107 397085
rect 318628 397080 378107 397082
rect 318628 397024 378046 397080
rect 378102 397024 378107 397080
rect 318628 397022 378107 397024
rect 318628 397020 318634 397022
rect 378041 397019 378107 397022
rect 315798 396884 315804 396948
rect 315868 396946 315874 396948
rect 375782 396946 375788 396948
rect 315868 396886 375788 396946
rect 315868 396884 315874 396886
rect 375782 396884 375788 396886
rect 375852 396884 375858 396948
rect 380198 396884 380204 396948
rect 380268 396946 380274 396948
rect 390829 396946 390895 396949
rect 380268 396944 390895 396946
rect 380268 396888 390834 396944
rect 390890 396888 390895 396944
rect 380268 396886 390895 396888
rect 380268 396884 380274 396886
rect 390829 396883 390895 396886
rect 260741 396810 260807 396813
rect 343357 396810 343423 396813
rect 260741 396808 343423 396810
rect 260741 396752 260746 396808
rect 260802 396752 343362 396808
rect 343418 396752 343423 396808
rect 260741 396750 343423 396752
rect 260741 396747 260807 396750
rect 343357 396747 343423 396750
rect 349245 396810 349311 396813
rect 350206 396810 350212 396812
rect 349245 396808 350212 396810
rect 349245 396752 349250 396808
rect 349306 396752 350212 396808
rect 349245 396750 350212 396752
rect 349245 396747 349311 396750
rect 350206 396748 350212 396750
rect 350276 396748 350282 396812
rect 350717 396810 350783 396813
rect 350942 396810 350948 396812
rect 350717 396808 350948 396810
rect 350717 396752 350722 396808
rect 350778 396752 350948 396808
rect 350717 396750 350948 396752
rect 350717 396747 350783 396750
rect 350942 396748 350948 396750
rect 351012 396748 351018 396812
rect 357934 396748 357940 396812
rect 358004 396810 358010 396812
rect 361062 396810 361068 396812
rect 358004 396750 361068 396810
rect 358004 396748 358010 396750
rect 361062 396748 361068 396750
rect 361132 396748 361138 396812
rect 266261 396674 266327 396677
rect 347773 396674 347839 396677
rect 354949 396676 355015 396677
rect 354949 396674 354996 396676
rect 266261 396672 347839 396674
rect 266261 396616 266266 396672
rect 266322 396616 347778 396672
rect 347834 396616 347839 396672
rect 266261 396614 347839 396616
rect 354904 396672 354996 396674
rect 354904 396616 354954 396672
rect 354904 396614 354996 396616
rect 266261 396611 266327 396614
rect 347773 396611 347839 396614
rect 354949 396612 354996 396614
rect 355060 396612 355066 396676
rect 358353 396674 358419 396677
rect 373942 396674 373948 396676
rect 358353 396672 373948 396674
rect 358353 396616 358358 396672
rect 358414 396616 373948 396672
rect 358353 396614 373948 396616
rect 354949 396611 355015 396612
rect 358353 396611 358419 396614
rect 373942 396612 373948 396614
rect 374012 396612 374018 396676
rect 330569 396538 330635 396541
rect 352557 396538 352623 396541
rect 330569 396536 352623 396538
rect 330569 396480 330574 396536
rect 330630 396480 352562 396536
rect 352618 396480 352623 396536
rect 330569 396478 352623 396480
rect 330569 396475 330635 396478
rect 352557 396475 352623 396478
rect 359273 396538 359339 396541
rect 359406 396538 359412 396540
rect 359273 396536 359412 396538
rect 359273 396480 359278 396536
rect 359334 396480 359412 396536
rect 359273 396478 359412 396480
rect 359273 396475 359339 396478
rect 359406 396476 359412 396478
rect 359476 396476 359482 396540
rect 345013 396132 345079 396133
rect 345013 396128 345060 396132
rect 345124 396130 345130 396132
rect 345013 396072 345018 396128
rect 345013 396068 345060 396072
rect 345124 396070 345170 396130
rect 345124 396068 345130 396070
rect 357014 396068 357020 396132
rect 357084 396130 357090 396132
rect 368054 396130 368060 396132
rect 357084 396070 368060 396130
rect 357084 396068 357090 396070
rect 368054 396068 368060 396070
rect 368124 396068 368130 396132
rect 385166 396068 385172 396132
rect 385236 396130 385242 396132
rect 385585 396130 385651 396133
rect 385236 396128 385651 396130
rect 385236 396072 385590 396128
rect 385646 396072 385651 396128
rect 385236 396070 385651 396072
rect 385236 396068 385242 396070
rect 345013 396067 345079 396068
rect 385585 396067 385651 396070
rect 283414 395932 283420 395996
rect 283484 395994 283490 395996
rect 304993 395994 305059 395997
rect 283484 395992 305059 395994
rect 283484 395936 304998 395992
rect 305054 395936 305059 395992
rect 283484 395934 305059 395936
rect 283484 395932 283490 395934
rect 304993 395931 305059 395934
rect 313038 395932 313044 395996
rect 313108 395994 313114 395996
rect 365161 395994 365227 395997
rect 367185 395994 367251 395997
rect 313108 395934 350550 395994
rect 313108 395932 313114 395934
rect 273989 395858 274055 395861
rect 335813 395858 335879 395861
rect 273989 395856 335879 395858
rect 273989 395800 273994 395856
rect 274050 395800 335818 395856
rect 335874 395800 335879 395856
rect 273989 395798 335879 395800
rect 273989 395795 274055 395798
rect 335813 395795 335879 395798
rect 343582 395796 343588 395860
rect 343652 395858 343658 395860
rect 344185 395858 344251 395861
rect 343652 395856 344251 395858
rect 343652 395800 344190 395856
rect 344246 395800 344251 395856
rect 343652 395798 344251 395800
rect 350490 395858 350550 395934
rect 365161 395992 367251 395994
rect 365161 395936 365166 395992
rect 365222 395936 367190 395992
rect 367246 395936 367251 395992
rect 365161 395934 367251 395936
rect 365161 395931 365227 395934
rect 367185 395931 367251 395934
rect 372705 395858 372771 395861
rect 350490 395856 372771 395858
rect 350490 395800 372710 395856
rect 372766 395800 372771 395856
rect 350490 395798 372771 395800
rect 343652 395796 343658 395798
rect 344185 395795 344251 395798
rect 372705 395795 372771 395798
rect 271413 395722 271479 395725
rect 347497 395722 347563 395725
rect 271413 395720 347563 395722
rect 271413 395664 271418 395720
rect 271474 395664 347502 395720
rect 347558 395664 347563 395720
rect 271413 395662 347563 395664
rect 271413 395659 271479 395662
rect 347497 395659 347563 395662
rect 363270 395660 363276 395724
rect 363340 395722 363346 395724
rect 369025 395722 369091 395725
rect 363340 395720 369091 395722
rect 363340 395664 369030 395720
rect 369086 395664 369091 395720
rect 363340 395662 369091 395664
rect 363340 395660 363346 395662
rect 369025 395659 369091 395662
rect 277117 395586 277183 395589
rect 354305 395586 354371 395589
rect 277117 395584 354371 395586
rect 277117 395528 277122 395584
rect 277178 395528 354310 395584
rect 354366 395528 354371 395584
rect 277117 395526 354371 395528
rect 277117 395523 277183 395526
rect 354305 395523 354371 395526
rect 355174 395524 355180 395588
rect 355244 395586 355250 395588
rect 364057 395586 364123 395589
rect 355244 395584 364123 395586
rect 355244 395528 364062 395584
rect 364118 395528 364123 395584
rect 355244 395526 364123 395528
rect 355244 395524 355250 395526
rect 364057 395523 364123 395526
rect 266997 395450 267063 395453
rect 342253 395450 342319 395453
rect 266997 395448 342319 395450
rect 266997 395392 267002 395448
rect 267058 395392 342258 395448
rect 342314 395392 342319 395448
rect 266997 395390 342319 395392
rect 266997 395387 267063 395390
rect 342253 395387 342319 395390
rect 346117 395450 346183 395453
rect 347078 395450 347084 395452
rect 346117 395448 347084 395450
rect 346117 395392 346122 395448
rect 346178 395392 347084 395448
rect 346117 395390 347084 395392
rect 346117 395387 346183 395390
rect 347078 395388 347084 395390
rect 347148 395388 347154 395452
rect 347814 395388 347820 395452
rect 347884 395450 347890 395452
rect 348141 395450 348207 395453
rect 347884 395448 348207 395450
rect 347884 395392 348146 395448
rect 348202 395392 348207 395448
rect 347884 395390 348207 395392
rect 347884 395388 347890 395390
rect 348141 395387 348207 395390
rect 349838 395388 349844 395452
rect 349908 395450 349914 395452
rect 349981 395450 350047 395453
rect 349908 395448 350047 395450
rect 349908 395392 349986 395448
rect 350042 395392 350047 395448
rect 349908 395390 350047 395392
rect 349908 395388 349914 395390
rect 349981 395387 350047 395390
rect 359406 395388 359412 395452
rect 359476 395450 359482 395452
rect 364374 395450 364380 395452
rect 359476 395390 364380 395450
rect 359476 395388 359482 395390
rect 364374 395388 364380 395390
rect 364444 395388 364450 395452
rect 270401 395314 270467 395317
rect 354213 395314 354279 395317
rect 270401 395312 354279 395314
rect 270401 395256 270406 395312
rect 270462 395256 354218 395312
rect 354274 395256 354279 395312
rect 270401 395254 354279 395256
rect 270401 395251 270467 395254
rect 354213 395251 354279 395254
rect 358118 395252 358124 395316
rect 358188 395314 358194 395316
rect 358537 395314 358603 395317
rect 358188 395312 358603 395314
rect 358188 395256 358542 395312
rect 358598 395256 358603 395312
rect 358188 395254 358603 395256
rect 358188 395252 358194 395254
rect 358537 395251 358603 395254
rect 364374 395252 364380 395316
rect 364444 395314 364450 395316
rect 364517 395314 364583 395317
rect 364444 395312 364583 395314
rect 364444 395256 364522 395312
rect 364578 395256 364583 395312
rect 364444 395254 364583 395256
rect 364444 395252 364450 395254
rect 364517 395251 364583 395254
rect 374453 395314 374519 395317
rect 375046 395314 375052 395316
rect 374453 395312 375052 395314
rect 374453 395256 374458 395312
rect 374514 395256 375052 395312
rect 374453 395254 375052 395256
rect 374453 395251 374519 395254
rect 375046 395252 375052 395254
rect 375116 395252 375122 395316
rect 378317 395314 378383 395317
rect 378726 395314 378732 395316
rect 378317 395312 378732 395314
rect 378317 395256 378322 395312
rect 378378 395256 378732 395312
rect 378317 395254 378732 395256
rect 378317 395251 378383 395254
rect 378726 395252 378732 395254
rect 378796 395252 378802 395316
rect 378910 395252 378916 395316
rect 378980 395314 378986 395316
rect 379145 395314 379211 395317
rect 378980 395312 379211 395314
rect 378980 395256 379150 395312
rect 379206 395256 379211 395312
rect 378980 395254 379211 395256
rect 378980 395252 378986 395254
rect 379145 395251 379211 395254
rect 283598 395116 283604 395180
rect 283668 395178 283674 395180
rect 305085 395178 305151 395181
rect 283668 395176 305151 395178
rect 283668 395120 305090 395176
rect 305146 395120 305151 395176
rect 283668 395118 305151 395120
rect 283668 395116 283674 395118
rect 305085 395115 305151 395118
rect 334893 395178 334959 395181
rect 364701 395178 364767 395181
rect 334893 395176 364767 395178
rect 334893 395120 334898 395176
rect 334954 395120 364706 395176
rect 364762 395120 364767 395176
rect 334893 395118 364767 395120
rect 334893 395115 334959 395118
rect 364701 395115 364767 395118
rect 346393 395042 346459 395045
rect 346710 395042 346716 395044
rect 346393 395040 346716 395042
rect 346393 394984 346398 395040
rect 346454 394984 346716 395040
rect 346393 394982 346716 394984
rect 346393 394979 346459 394982
rect 346710 394980 346716 394982
rect 346780 394980 346786 395044
rect 347313 395042 347379 395045
rect 349102 395042 349108 395044
rect 347313 395040 349108 395042
rect 347313 394984 347318 395040
rect 347374 394984 349108 395040
rect 347313 394982 349108 394984
rect 347313 394979 347379 394982
rect 349102 394980 349108 394982
rect 349172 394980 349178 395044
rect 358997 395042 359063 395045
rect 359774 395042 359780 395044
rect 358997 395040 359780 395042
rect 358997 394984 359002 395040
rect 359058 394984 359780 395040
rect 358997 394982 359780 394984
rect 358997 394979 359063 394982
rect 359774 394980 359780 394982
rect 359844 394980 359850 395044
rect 364517 395042 364583 395045
rect 364926 395042 364932 395044
rect 364517 395040 364932 395042
rect 364517 394984 364522 395040
rect 364578 394984 364932 395040
rect 364517 394982 364932 394984
rect 364517 394979 364583 394982
rect 364926 394980 364932 394982
rect 364996 394980 365002 395044
rect 347865 394906 347931 394909
rect 348734 394906 348740 394908
rect 347865 394904 348740 394906
rect 347865 394848 347870 394904
rect 347926 394848 348740 394904
rect 347865 394846 348740 394848
rect 347865 394843 347931 394846
rect 348734 394844 348740 394846
rect 348804 394844 348810 394908
rect 295558 394436 295564 394500
rect 295628 394498 295634 394500
rect 356421 394498 356487 394501
rect 295628 394496 356487 394498
rect 295628 394440 356426 394496
rect 356482 394440 356487 394496
rect 295628 394438 356487 394440
rect 295628 394436 295634 394438
rect 356421 394435 356487 394438
rect 363229 394498 363295 394501
rect 363822 394498 363828 394500
rect 363229 394496 363828 394498
rect 363229 394440 363234 394496
rect 363290 394440 363828 394496
rect 363229 394438 363828 394440
rect 363229 394435 363295 394438
rect 363822 394436 363828 394438
rect 363892 394436 363898 394500
rect 286910 394300 286916 394364
rect 286980 394362 286986 394364
rect 343633 394362 343699 394365
rect 286980 394360 343699 394362
rect 286980 394304 343638 394360
rect 343694 394304 343699 394360
rect 286980 394302 343699 394304
rect 286980 394300 286986 394302
rect 343633 394299 343699 394302
rect 296110 394164 296116 394228
rect 296180 394226 296186 394228
rect 352005 394226 352071 394229
rect 296180 394224 352071 394226
rect 296180 394168 352010 394224
rect 352066 394168 352071 394224
rect 296180 394166 352071 394168
rect 296180 394164 296186 394166
rect 352005 394163 352071 394166
rect 268653 394090 268719 394093
rect 352046 394090 352052 394092
rect 268653 394088 352052 394090
rect 268653 394032 268658 394088
rect 268714 394032 352052 394088
rect 268653 394030 352052 394032
rect 268653 394027 268719 394030
rect 352046 394028 352052 394030
rect 352116 394028 352122 394092
rect 271689 393954 271755 393957
rect 358670 393954 358676 393956
rect 271689 393952 358676 393954
rect 271689 393896 271694 393952
rect 271750 393896 358676 393952
rect 271689 393894 358676 393896
rect 271689 393891 271755 393894
rect 358670 393892 358676 393894
rect 358740 393892 358746 393956
rect 370681 393954 370747 393957
rect 371366 393954 371372 393956
rect 370681 393952 371372 393954
rect 370681 393896 370686 393952
rect 370742 393896 371372 393952
rect 370681 393894 371372 393896
rect 370681 393891 370747 393894
rect 371366 393892 371372 393894
rect 371436 393892 371442 393956
rect 297950 393756 297956 393820
rect 298020 393818 298026 393820
rect 356881 393818 356947 393821
rect 298020 393816 356947 393818
rect 298020 393760 356886 393816
rect 356942 393760 356947 393816
rect 298020 393758 356947 393760
rect 298020 393756 298026 393758
rect 356881 393755 356947 393758
rect 296478 393620 296484 393684
rect 296548 393682 296554 393684
rect 355961 393682 356027 393685
rect 296548 393680 356027 393682
rect 296548 393624 355966 393680
rect 356022 393624 356027 393680
rect 296548 393622 356027 393624
rect 296548 393620 296554 393622
rect 355961 393619 356027 393622
rect 350625 393546 350691 393549
rect 351126 393546 351132 393548
rect 350625 393544 351132 393546
rect 350625 393488 350630 393544
rect 350686 393488 351132 393544
rect 350625 393486 351132 393488
rect 350625 393483 350691 393486
rect 351126 393484 351132 393486
rect 351196 393484 351202 393548
rect 380893 393546 380959 393549
rect 381118 393546 381124 393548
rect 380893 393544 381124 393546
rect 380893 393488 380898 393544
rect 380954 393488 381124 393544
rect 380893 393486 381124 393488
rect 380893 393483 380959 393486
rect 381118 393484 381124 393486
rect 381188 393484 381194 393548
rect 302182 393076 302188 393140
rect 302252 393138 302258 393140
rect 362769 393138 362835 393141
rect 302252 393136 362835 393138
rect 302252 393080 362774 393136
rect 362830 393080 362835 393136
rect 302252 393078 362835 393080
rect 302252 393076 302258 393078
rect 362769 393075 362835 393078
rect 301998 392940 302004 393004
rect 302068 393002 302074 393004
rect 361246 393002 361252 393004
rect 302068 392942 361252 393002
rect 302068 392940 302074 392942
rect 361246 392940 361252 392942
rect 361316 392940 361322 393004
rect 297030 392804 297036 392868
rect 297100 392866 297106 392868
rect 357566 392866 357572 392868
rect 297100 392806 357572 392866
rect 297100 392804 297106 392806
rect 357566 392804 357572 392806
rect 357636 392804 357642 392868
rect 285121 392730 285187 392733
rect 364333 392730 364399 392733
rect 285121 392728 364399 392730
rect 285121 392672 285126 392728
rect 285182 392672 364338 392728
rect 364394 392672 364399 392728
rect 285121 392670 364399 392672
rect 285121 392667 285187 392670
rect 364333 392667 364399 392670
rect 368473 392730 368539 392733
rect 368606 392730 368612 392732
rect 368473 392728 368612 392730
rect 368473 392672 368478 392728
rect 368534 392672 368612 392728
rect 368473 392670 368612 392672
rect 368473 392667 368539 392670
rect 368606 392668 368612 392670
rect 368676 392668 368682 392732
rect 271781 392594 271847 392597
rect 360510 392594 360516 392596
rect 271781 392592 360516 392594
rect 271781 392536 271786 392592
rect 271842 392536 360516 392592
rect 271781 392534 360516 392536
rect 271781 392531 271847 392534
rect 360510 392532 360516 392534
rect 360580 392532 360586 392596
rect 298502 392396 298508 392460
rect 298572 392458 298578 392460
rect 357525 392458 357591 392461
rect 298572 392456 357591 392458
rect 298572 392400 357530 392456
rect 357586 392400 357591 392456
rect 298572 392398 357591 392400
rect 298572 392396 298578 392398
rect 357525 392395 357591 392398
rect 292982 392260 292988 392324
rect 293052 392322 293058 392324
rect 353109 392322 353175 392325
rect 293052 392320 353175 392322
rect 293052 392264 353114 392320
rect 353170 392264 353175 392320
rect 293052 392262 353175 392264
rect 293052 392260 293058 392262
rect 353109 392259 353175 392262
rect 373993 392186 374059 392189
rect 374494 392186 374500 392188
rect 373993 392184 374500 392186
rect 373993 392128 373998 392184
rect 374054 392128 374500 392184
rect 373993 392126 374500 392128
rect 373993 392123 374059 392126
rect 374494 392124 374500 392126
rect 374564 392124 374570 392188
rect 285070 391852 285076 391916
rect 285140 391914 285146 391916
rect 309961 391914 310027 391917
rect 285140 391912 310027 391914
rect 285140 391856 309966 391912
rect 310022 391856 310027 391912
rect 285140 391854 310027 391856
rect 285140 391852 285146 391854
rect 309961 391851 310027 391854
rect 310278 391852 310284 391916
rect 310348 391914 310354 391916
rect 369393 391914 369459 391917
rect 310348 391912 369459 391914
rect 310348 391856 369398 391912
rect 369454 391856 369459 391912
rect 310348 391854 369459 391856
rect 310348 391852 310354 391854
rect 369393 391851 369459 391854
rect 295190 391716 295196 391780
rect 295260 391778 295266 391780
rect 353845 391778 353911 391781
rect 295260 391776 353911 391778
rect 295260 391720 353850 391776
rect 353906 391720 353911 391776
rect 295260 391718 353911 391720
rect 295260 391716 295266 391718
rect 353845 391715 353911 391718
rect 295006 391580 295012 391644
rect 295076 391642 295082 391644
rect 354029 391642 354095 391645
rect 295076 391640 354095 391642
rect 295076 391584 354034 391640
rect 354090 391584 354095 391640
rect 583520 391628 584960 391868
rect 295076 391582 354095 391584
rect 295076 391580 295082 391582
rect 354029 391579 354095 391582
rect 292798 391444 292804 391508
rect 292868 391506 292874 391508
rect 353753 391506 353819 391509
rect 292868 391504 353819 391506
rect 292868 391448 353758 391504
rect 353814 391448 353819 391504
rect 292868 391446 353819 391448
rect 292868 391444 292874 391446
rect 353753 391443 353819 391446
rect 275553 391370 275619 391373
rect 349286 391370 349292 391372
rect 275553 391368 349292 391370
rect 275553 391312 275558 391368
rect 275614 391312 349292 391368
rect 275553 391310 349292 391312
rect 275553 391307 275619 391310
rect 349286 391308 349292 391310
rect 349356 391308 349362 391372
rect 375414 391308 375420 391372
rect 375484 391370 375490 391372
rect 376017 391370 376083 391373
rect 375484 391368 376083 391370
rect 375484 391312 376022 391368
rect 376078 391312 376083 391368
rect 375484 391310 376083 391312
rect 375484 391308 375490 391310
rect 376017 391307 376083 391310
rect 266077 391234 266143 391237
rect 343725 391234 343791 391237
rect 266077 391232 343791 391234
rect 266077 391176 266082 391232
rect 266138 391176 343730 391232
rect 343786 391176 343791 391232
rect 266077 391174 343791 391176
rect 266077 391171 266143 391174
rect 343725 391171 343791 391174
rect 288934 391036 288940 391100
rect 289004 391098 289010 391100
rect 345105 391098 345171 391101
rect 289004 391096 345171 391098
rect 289004 391040 345110 391096
rect 345166 391040 345171 391096
rect 289004 391038 345171 391040
rect 289004 391036 289010 391038
rect 345105 391035 345171 391038
rect 307702 390628 307708 390692
rect 307772 390690 307778 390692
rect 307937 390690 308003 390693
rect 307772 390688 308003 390690
rect 307772 390632 307942 390688
rect 307998 390632 308003 390688
rect 307772 390630 308003 390632
rect 307772 390628 307778 390630
rect 307937 390627 308003 390630
rect 317270 390492 317276 390556
rect 317340 390554 317346 390556
rect 376661 390554 376727 390557
rect 317340 390552 376727 390554
rect 317340 390496 376666 390552
rect 376722 390496 376727 390552
rect 317340 390494 376727 390496
rect 317340 390492 317346 390494
rect 376661 390491 376727 390494
rect 320030 390356 320036 390420
rect 320100 390418 320106 390420
rect 380525 390418 380591 390421
rect 320100 390416 380591 390418
rect 320100 390360 380530 390416
rect 380586 390360 380591 390416
rect 320100 390358 380591 390360
rect 320100 390356 320106 390358
rect 380525 390355 380591 390358
rect 294638 390220 294644 390284
rect 294708 390282 294714 390284
rect 353293 390282 353359 390285
rect 294708 390280 353359 390282
rect 294708 390224 353298 390280
rect 353354 390224 353359 390280
rect 294708 390222 353359 390224
rect 294708 390220 294714 390222
rect 353293 390219 353359 390222
rect 354029 390282 354095 390285
rect 357014 390282 357020 390284
rect 354029 390280 357020 390282
rect 354029 390224 354034 390280
rect 354090 390224 357020 390280
rect 354029 390222 357020 390224
rect 354029 390219 354095 390222
rect 357014 390220 357020 390222
rect 357084 390220 357090 390284
rect 317086 390084 317092 390148
rect 317156 390146 317162 390148
rect 377857 390146 377923 390149
rect 317156 390144 377923 390146
rect 317156 390088 377862 390144
rect 377918 390088 377923 390144
rect 317156 390086 377923 390088
rect 317156 390084 317162 390086
rect 377857 390083 377923 390086
rect 260649 390010 260715 390013
rect 324221 390010 324287 390013
rect 260649 390008 324287 390010
rect 260649 389952 260654 390008
rect 260710 389952 324226 390008
rect 324282 389952 324287 390008
rect 260649 389950 324287 389952
rect 260649 389947 260715 389950
rect 324221 389947 324287 389950
rect 262029 389874 262095 389877
rect 346710 389874 346716 389876
rect 262029 389872 346716 389874
rect 262029 389816 262034 389872
rect 262090 389816 346716 389872
rect 262029 389814 346716 389816
rect 262029 389811 262095 389814
rect 346710 389812 346716 389814
rect 346780 389812 346786 389876
rect 294822 389676 294828 389740
rect 294892 389738 294898 389740
rect 354305 389738 354371 389741
rect 294892 389736 354371 389738
rect 294892 389680 354310 389736
rect 354366 389680 354371 389736
rect 294892 389678 354371 389680
rect 294892 389676 294898 389678
rect 354305 389675 354371 389678
rect 342253 389194 342319 389197
rect 348182 389194 348188 389196
rect 342253 389192 348188 389194
rect 342253 389136 342258 389192
rect 342314 389136 348188 389192
rect 342253 389134 348188 389136
rect 342253 389131 342319 389134
rect 348182 389132 348188 389134
rect 348252 389132 348258 389196
rect 344134 388996 344140 389060
rect 344204 389058 344210 389060
rect 383878 389058 383884 389060
rect 344204 388998 383884 389058
rect 344204 388996 344210 388998
rect 383878 388996 383884 388998
rect 383948 388996 383954 389060
rect 286358 388860 286364 388924
rect 286428 388922 286434 388924
rect 345381 388922 345447 388925
rect 286428 388920 345447 388922
rect 286428 388864 345386 388920
rect 345442 388864 345447 388920
rect 286428 388862 345447 388864
rect 286428 388860 286434 388862
rect 345381 388859 345447 388862
rect 288198 388724 288204 388788
rect 288268 388786 288274 388788
rect 348417 388786 348483 388789
rect 288268 388784 348483 388786
rect 288268 388728 348422 388784
rect 348478 388728 348483 388784
rect 288268 388726 348483 388728
rect 288268 388724 288274 388726
rect 348417 388723 348483 388726
rect 289486 388588 289492 388652
rect 289556 388650 289562 388652
rect 349521 388650 349587 388653
rect 289556 388648 349587 388650
rect 289556 388592 349526 388648
rect 349582 388592 349587 388648
rect 289556 388590 349587 388592
rect 289556 388588 289562 388590
rect 349521 388587 349587 388590
rect 272517 388514 272583 388517
rect 345238 388514 345244 388516
rect 272517 388512 345244 388514
rect 272517 388456 272522 388512
rect 272578 388456 345244 388512
rect 272517 388454 345244 388456
rect 272517 388451 272583 388454
rect 345238 388452 345244 388454
rect 345308 388452 345314 388516
rect 346209 388514 346275 388517
rect 385350 388514 385356 388516
rect 346209 388512 385356 388514
rect 346209 388456 346214 388512
rect 346270 388456 385356 388512
rect 346209 388454 385356 388456
rect 346209 388451 346275 388454
rect 385350 388452 385356 388454
rect 385420 388452 385426 388516
rect 259269 388378 259335 388381
rect 347998 388378 348004 388380
rect 259269 388376 348004 388378
rect 259269 388320 259274 388376
rect 259330 388320 348004 388376
rect 259269 388318 348004 388320
rect 259269 388315 259335 388318
rect 347998 388316 348004 388318
rect 348068 388316 348074 388380
rect 344645 388242 344711 388245
rect 363638 388242 363644 388244
rect 344645 388240 363644 388242
rect 344645 388184 344650 388240
rect 344706 388184 363644 388240
rect 344645 388182 363644 388184
rect 344645 388179 344711 388182
rect 363638 388180 363644 388182
rect 363708 388180 363714 388244
rect 312721 387698 312787 387701
rect 371550 387698 371556 387700
rect 312721 387696 371556 387698
rect 312721 387640 312726 387696
rect 312782 387640 371556 387696
rect 312721 387638 371556 387640
rect 312721 387635 312787 387638
rect 371550 387636 371556 387638
rect 371620 387636 371626 387700
rect 348417 387562 348483 387565
rect 356462 387562 356468 387564
rect 348417 387560 356468 387562
rect 348417 387504 348422 387560
rect 348478 387504 356468 387560
rect 348417 387502 356468 387504
rect 348417 387499 348483 387502
rect 356462 387500 356468 387502
rect 356532 387500 356538 387564
rect 283782 387364 283788 387428
rect 283852 387426 283858 387428
rect 343449 387426 343515 387429
rect 283852 387424 343515 387426
rect 283852 387368 343454 387424
rect 343510 387368 343515 387424
rect 283852 387366 343515 387368
rect 283852 387364 283858 387366
rect 343449 387363 343515 387366
rect 297582 387228 297588 387292
rect 297652 387290 297658 387292
rect 357801 387290 357867 387293
rect 297652 387288 357867 387290
rect 297652 387232 357806 387288
rect 357862 387232 357867 387288
rect 297652 387230 357867 387232
rect 297652 387228 297658 387230
rect 357801 387227 357867 387230
rect 269665 387154 269731 387157
rect 359038 387154 359044 387156
rect 269665 387152 359044 387154
rect 269665 387096 269670 387152
rect 269726 387096 359044 387152
rect 269665 387094 359044 387096
rect 269665 387091 269731 387094
rect 359038 387092 359044 387094
rect 359108 387092 359114 387156
rect 285438 386956 285444 387020
rect 285508 387018 285514 387020
rect 344185 387018 344251 387021
rect 577497 387018 577563 387021
rect 285508 387016 344251 387018
rect 285508 386960 344190 387016
rect 344246 386960 344251 387016
rect 285508 386958 344251 386960
rect 285508 386956 285514 386958
rect 344185 386955 344251 386958
rect 354630 387016 577563 387018
rect 354630 386960 577502 387016
rect 577558 386960 577563 387016
rect 354630 386958 577563 386960
rect 343030 386820 343036 386884
rect 343100 386882 343106 386884
rect 349654 386882 349660 386884
rect 343100 386822 349660 386882
rect 343100 386820 343106 386822
rect 349654 386820 349660 386822
rect 349724 386882 349730 386884
rect 354630 386882 354690 386958
rect 577497 386955 577563 386958
rect 349724 386822 354690 386882
rect 349724 386820 349730 386822
rect 342846 386684 342852 386748
rect 342916 386746 342922 386748
rect 380157 386746 380223 386749
rect 342916 386744 380223 386746
rect 342916 386688 380162 386744
rect 380218 386688 380223 386744
rect 342916 386686 380223 386688
rect 342916 386684 342922 386686
rect 380157 386683 380223 386686
rect 329373 386066 329439 386069
rect 368974 386066 368980 386068
rect 329373 386064 368980 386066
rect 329373 386008 329378 386064
rect 329434 386008 368980 386064
rect 329373 386006 368980 386008
rect 329373 386003 329439 386006
rect 368974 386004 368980 386006
rect 369044 386004 369050 386068
rect 330518 385868 330524 385932
rect 330588 385930 330594 385932
rect 381537 385930 381603 385933
rect 330588 385928 381603 385930
rect 330588 385872 381542 385928
rect 381598 385872 381603 385928
rect 330588 385870 381603 385872
rect 330588 385868 330594 385870
rect 381537 385867 381603 385870
rect 286542 385732 286548 385796
rect 286612 385794 286618 385796
rect 302969 385794 303035 385797
rect 286612 385792 303035 385794
rect 286612 385736 302974 385792
rect 303030 385736 303035 385792
rect 286612 385734 303035 385736
rect 286612 385732 286618 385734
rect 302969 385731 303035 385734
rect 324313 385794 324379 385797
rect 382958 385794 382964 385796
rect 324313 385792 382964 385794
rect 324313 385736 324318 385792
rect 324374 385736 382964 385792
rect 324313 385734 382964 385736
rect 324313 385731 324379 385734
rect 382958 385732 382964 385734
rect 383028 385732 383034 385796
rect 269573 385658 269639 385661
rect 353334 385658 353340 385660
rect 269573 385656 353340 385658
rect 269573 385600 269578 385656
rect 269634 385600 353340 385656
rect 269573 385598 353340 385600
rect 269573 385595 269639 385598
rect 353334 385596 353340 385598
rect 353404 385596 353410 385660
rect -960 384284 480 384524
rect 295926 384372 295932 384436
rect 295996 384434 296002 384436
rect 352281 384434 352347 384437
rect 295996 384432 352347 384434
rect 295996 384376 352286 384432
rect 352342 384376 352347 384432
rect 295996 384374 352347 384376
rect 295996 384372 296002 384374
rect 352281 384371 352347 384374
rect 279141 384298 279207 384301
rect 370262 384298 370268 384300
rect 279141 384296 370268 384298
rect 279141 384240 279146 384296
rect 279202 384240 370268 384296
rect 279141 384238 370268 384240
rect 279141 384235 279207 384238
rect 370262 384236 370268 384238
rect 370332 384236 370338 384300
rect 343265 383482 343331 383485
rect 355358 383482 355364 383484
rect 343265 383480 355364 383482
rect 343265 383424 343270 383480
rect 343326 383424 355364 383480
rect 343265 383422 355364 383424
rect 343265 383419 343331 383422
rect 355358 383420 355364 383422
rect 355428 383420 355434 383484
rect 347497 383346 347563 383349
rect 364558 383346 364564 383348
rect 347497 383344 364564 383346
rect 347497 383288 347502 383344
rect 347558 383288 364564 383344
rect 347497 383286 364564 383288
rect 347497 383283 347563 383286
rect 364558 383284 364564 383286
rect 364628 383284 364634 383348
rect 304942 383148 304948 383212
rect 305012 383210 305018 383212
rect 366265 383210 366331 383213
rect 305012 383208 366331 383210
rect 305012 383152 366270 383208
rect 366326 383152 366331 383208
rect 305012 383150 366331 383152
rect 305012 383148 305018 383150
rect 366265 383147 366331 383150
rect 272793 383074 272859 383077
rect 351862 383074 351868 383076
rect 272793 383072 351868 383074
rect 272793 383016 272798 383072
rect 272854 383016 351868 383072
rect 272793 383014 351868 383016
rect 272793 383011 272859 383014
rect 351862 383012 351868 383014
rect 351932 383012 351938 383076
rect 275461 382938 275527 382941
rect 356830 382938 356836 382940
rect 275461 382936 356836 382938
rect 275461 382880 275466 382936
rect 275522 382880 356836 382936
rect 275461 382878 356836 382880
rect 275461 382875 275527 382878
rect 356830 382876 356836 382878
rect 356900 382876 356906 382940
rect 285254 381788 285260 381852
rect 285324 381850 285330 381852
rect 300393 381850 300459 381853
rect 285324 381848 300459 381850
rect 285324 381792 300398 381848
rect 300454 381792 300459 381848
rect 285324 381790 300459 381792
rect 285324 381788 285330 381790
rect 300393 381787 300459 381790
rect 290958 381652 290964 381716
rect 291028 381714 291034 381716
rect 345841 381714 345907 381717
rect 291028 381712 345907 381714
rect 291028 381656 345846 381712
rect 345902 381656 345907 381712
rect 291028 381654 345907 381656
rect 291028 381652 291034 381654
rect 345841 381651 345907 381654
rect 299974 381516 299980 381580
rect 300044 381578 300050 381580
rect 357617 381578 357683 381581
rect 300044 381576 357683 381578
rect 300044 381520 357622 381576
rect 357678 381520 357683 381576
rect 300044 381518 357683 381520
rect 300044 381516 300050 381518
rect 357617 381515 357683 381518
rect 297398 380156 297404 380220
rect 297468 380218 297474 380220
rect 355593 380218 355659 380221
rect 297468 380216 355659 380218
rect 297468 380160 355598 380216
rect 355654 380160 355659 380216
rect 297468 380158 355659 380160
rect 297468 380156 297474 380158
rect 355593 380155 355659 380158
rect 290774 379340 290780 379404
rect 290844 379402 290850 379404
rect 348509 379402 348575 379405
rect 290844 379400 348575 379402
rect 290844 379344 348514 379400
rect 348570 379344 348575 379400
rect 290844 379342 348575 379344
rect 290844 379340 290850 379342
rect 348509 379339 348575 379342
rect 291878 379204 291884 379268
rect 291948 379266 291954 379268
rect 351453 379266 351519 379269
rect 291948 379264 351519 379266
rect 291948 379208 351458 379264
rect 351514 379208 351519 379264
rect 291948 379206 351519 379208
rect 291948 379204 291954 379206
rect 351453 379203 351519 379206
rect 292246 379068 292252 379132
rect 292316 379130 292322 379132
rect 350993 379130 351059 379133
rect 292316 379128 351059 379130
rect 292316 379072 350998 379128
rect 351054 379072 351059 379128
rect 292316 379070 351059 379072
rect 292316 379068 292322 379070
rect 350993 379067 351059 379070
rect 306966 378932 306972 378996
rect 307036 378994 307042 378996
rect 366582 378994 366588 378996
rect 307036 378934 366588 378994
rect 307036 378932 307042 378934
rect 366582 378932 366588 378934
rect 366652 378932 366658 378996
rect 289302 378796 289308 378860
rect 289372 378858 289378 378860
rect 349429 378858 349495 378861
rect 289372 378856 349495 378858
rect 289372 378800 349434 378856
rect 349490 378800 349495 378856
rect 289372 378798 349495 378800
rect 289372 378796 289378 378798
rect 349429 378795 349495 378798
rect 289118 378660 289124 378724
rect 289188 378722 289194 378724
rect 349981 378722 350047 378725
rect 289188 378720 350047 378722
rect 289188 378664 349986 378720
rect 350042 378664 350047 378720
rect 289188 378662 350047 378664
rect 289188 378660 289194 378662
rect 349981 378659 350047 378662
rect 580257 378450 580323 378453
rect 583520 378450 584960 378540
rect 580257 378448 584960 378450
rect 580257 378392 580262 378448
rect 580318 378392 584960 378448
rect 580257 378390 584960 378392
rect 580257 378387 580323 378390
rect 583520 378300 584960 378390
rect 314326 377708 314332 377772
rect 314396 377770 314402 377772
rect 374821 377770 374887 377773
rect 314396 377768 374887 377770
rect 314396 377712 374826 377768
rect 374882 377712 374887 377768
rect 314396 377710 374887 377712
rect 314396 377708 314402 377710
rect 374821 377707 374887 377710
rect 283966 377572 283972 377636
rect 284036 377634 284042 377636
rect 343582 377634 343588 377636
rect 284036 377574 343588 377634
rect 284036 377572 284042 377574
rect 343582 377572 343588 377574
rect 343652 377572 343658 377636
rect 349981 377634 350047 377637
rect 372654 377634 372660 377636
rect 349981 377632 372660 377634
rect 349981 377576 349986 377632
rect 350042 377576 372660 377632
rect 349981 377574 372660 377576
rect 349981 377571 350047 377574
rect 372654 377572 372660 377574
rect 372724 377572 372730 377636
rect 308990 377436 308996 377500
rect 309060 377498 309066 377500
rect 368841 377498 368907 377501
rect 309060 377496 368907 377498
rect 309060 377440 368846 377496
rect 368902 377440 368907 377496
rect 309060 377438 368907 377440
rect 309060 377436 309066 377438
rect 368841 377435 368907 377438
rect 292062 377300 292068 377364
rect 292132 377362 292138 377364
rect 352189 377362 352255 377365
rect 292132 377360 352255 377362
rect 292132 377304 352194 377360
rect 352250 377304 352255 377360
rect 292132 377302 352255 377304
rect 292132 377300 292138 377302
rect 352189 377299 352255 377302
rect 277894 375396 277900 375460
rect 277964 375458 277970 375460
rect 309777 375458 309843 375461
rect 277964 375456 309843 375458
rect 277964 375400 309782 375456
rect 309838 375400 309843 375456
rect 277964 375398 309843 375400
rect 277964 375396 277970 375398
rect 309777 375395 309843 375398
rect 306230 373492 306236 373556
rect 306300 373554 306306 373556
rect 364609 373554 364675 373557
rect 306300 373552 364675 373554
rect 306300 373496 364614 373552
rect 364670 373496 364675 373552
rect 306300 373494 364675 373496
rect 306300 373492 306306 373494
rect 364609 373491 364675 373494
rect 291694 373356 291700 373420
rect 291764 373418 291770 373420
rect 350901 373418 350967 373421
rect 291764 373416 350967 373418
rect 291764 373360 350906 373416
rect 350962 373360 350967 373416
rect 291764 373358 350967 373360
rect 291764 373356 291770 373358
rect 350901 373355 350967 373358
rect 307518 373220 307524 373284
rect 307588 373282 307594 373284
rect 367318 373282 367324 373284
rect 307588 373222 367324 373282
rect 307588 373220 307594 373222
rect 367318 373220 367324 373222
rect 367388 373220 367394 373284
rect 278446 372948 278452 373012
rect 278516 373010 278522 373012
rect 286685 373010 286751 373013
rect 278516 373008 286751 373010
rect 278516 372952 286690 373008
rect 286746 372952 286751 373008
rect 278516 372950 286751 372952
rect 278516 372948 278522 372950
rect 286685 372947 286751 372950
rect 222101 372874 222167 372877
rect 284569 372874 284635 372877
rect 222101 372872 284635 372874
rect 222101 372816 222106 372872
rect 222162 372816 284574 372872
rect 284630 372816 284635 372872
rect 222101 372814 284635 372816
rect 222101 372811 222167 372814
rect 284569 372811 284635 372814
rect 221222 372676 221228 372740
rect 221292 372738 221298 372740
rect 286041 372738 286107 372741
rect 221292 372736 286107 372738
rect 221292 372680 286046 372736
rect 286102 372680 286107 372736
rect 221292 372678 286107 372680
rect 221292 372676 221298 372678
rect 286041 372675 286107 372678
rect 290641 372330 290707 372333
rect 291837 372330 291903 372333
rect 324262 372330 324268 372332
rect 290641 372328 324268 372330
rect 290641 372272 290646 372328
rect 290702 372272 291842 372328
rect 291898 372272 324268 372328
rect 290641 372270 324268 372272
rect 290641 372267 290707 372270
rect 291837 372267 291903 372270
rect 324262 372268 324268 372270
rect 324332 372268 324338 372332
rect 281165 372194 281231 372197
rect 289997 372194 290063 372197
rect 281165 372192 290063 372194
rect 281165 372136 281170 372192
rect 281226 372136 290002 372192
rect 290058 372136 290063 372192
rect 281165 372134 290063 372136
rect 281165 372131 281231 372134
rect 289997 372131 290063 372134
rect 281441 372058 281507 372061
rect 293309 372058 293375 372061
rect 281441 372056 293375 372058
rect 281441 372000 281446 372056
rect 281502 372000 293314 372056
rect 293370 372000 293375 372056
rect 281441 371998 293375 372000
rect 281441 371995 281507 371998
rect 293309 371995 293375 371998
rect 282269 371924 282335 371925
rect 282269 371922 282316 371924
rect 282188 371920 282316 371922
rect 282380 371922 282386 371924
rect 297357 371922 297423 371925
rect 282380 371920 297423 371922
rect 282188 371864 282274 371920
rect 282380 371864 297362 371920
rect 297418 371864 297423 371920
rect 282188 371862 282316 371864
rect 282269 371860 282316 371862
rect 282380 371862 297423 371864
rect 282380 371860 282386 371862
rect 282269 371859 282335 371860
rect 297357 371859 297423 371862
rect 333973 371922 334039 371925
rect 344134 371922 344140 371924
rect 333973 371920 344140 371922
rect 333973 371864 333978 371920
rect 334034 371864 344140 371920
rect 333973 371862 344140 371864
rect 333973 371859 334039 371862
rect 344134 371860 344140 371862
rect 344204 371860 344210 371924
rect 281022 371724 281028 371788
rect 281092 371786 281098 371788
rect 310237 371786 310303 371789
rect 281092 371784 310303 371786
rect 281092 371728 310242 371784
rect 310298 371728 310303 371784
rect 281092 371726 310303 371728
rect 281092 371724 281098 371726
rect 310237 371723 310303 371726
rect 279366 371588 279372 371652
rect 279436 371650 279442 371652
rect 280705 371650 280771 371653
rect 279436 371648 280771 371650
rect 279436 371592 280710 371648
rect 280766 371592 280771 371648
rect 279436 371590 280771 371592
rect 279436 371588 279442 371590
rect 280705 371587 280771 371590
rect 280838 371588 280844 371652
rect 280908 371650 280914 371652
rect 310697 371650 310763 371653
rect 280908 371648 310763 371650
rect 280908 371592 310702 371648
rect 310758 371592 310763 371648
rect 280908 371590 310763 371592
rect 280908 371588 280914 371590
rect 310697 371587 310763 371590
rect -960 371378 480 371468
rect 276606 371452 276612 371516
rect 276676 371514 276682 371516
rect 289629 371514 289695 371517
rect 323158 371514 323164 371516
rect 276676 371512 323164 371514
rect 276676 371456 289634 371512
rect 289690 371456 323164 371512
rect 276676 371454 323164 371456
rect 276676 371452 276682 371454
rect 289629 371451 289695 371454
rect 323158 371452 323164 371454
rect 323228 371452 323234 371516
rect 3417 371378 3483 371381
rect -960 371376 3483 371378
rect -960 371320 3422 371376
rect 3478 371320 3483 371376
rect -960 371318 3483 371320
rect -960 371228 480 371318
rect 3417 371315 3483 371318
rect 242249 371378 242315 371381
rect 290641 371378 290707 371381
rect 242249 371376 290707 371378
rect 242249 371320 242254 371376
rect 242310 371320 290646 371376
rect 290702 371320 290707 371376
rect 242249 371318 290707 371320
rect 242249 371315 242315 371318
rect 290641 371315 290707 371318
rect 302969 370834 303035 370837
rect 324865 370834 324931 370837
rect 302969 370832 324931 370834
rect 302969 370776 302974 370832
rect 303030 370776 324870 370832
rect 324926 370776 324931 370832
rect 302969 370774 324931 370776
rect 302969 370771 303035 370774
rect 324865 370771 324931 370774
rect 289353 370698 289419 370701
rect 343030 370698 343036 370700
rect 289353 370696 343036 370698
rect 289353 370640 289358 370696
rect 289414 370640 343036 370696
rect 289353 370638 343036 370640
rect 289353 370635 289419 370638
rect 343030 370636 343036 370638
rect 343100 370636 343106 370700
rect 315614 370500 315620 370564
rect 315684 370562 315690 370564
rect 374545 370562 374611 370565
rect 315684 370560 374611 370562
rect 315684 370504 374550 370560
rect 374606 370504 374611 370560
rect 315684 370502 374611 370504
rect 315684 370500 315690 370502
rect 374545 370499 374611 370502
rect 253197 370426 253263 370429
rect 313549 370426 313615 370429
rect 253197 370424 313615 370426
rect 253197 370368 253202 370424
rect 253258 370368 313554 370424
rect 313610 370368 313615 370424
rect 253197 370366 313615 370368
rect 253197 370363 253263 370366
rect 313549 370363 313615 370366
rect 280654 370228 280660 370292
rect 280724 370290 280730 370292
rect 310605 370290 310671 370293
rect 280724 370288 310671 370290
rect 280724 370232 310610 370288
rect 310666 370232 310671 370288
rect 280724 370230 310671 370232
rect 280724 370228 280730 370230
rect 310605 370227 310671 370230
rect 224861 370154 224927 370157
rect 284937 370154 285003 370157
rect 224861 370152 285003 370154
rect 224861 370096 224866 370152
rect 224922 370096 284942 370152
rect 284998 370096 285003 370152
rect 224861 370094 285003 370096
rect 224861 370091 224927 370094
rect 284937 370091 285003 370094
rect 286041 370154 286107 370157
rect 300117 370154 300183 370157
rect 333094 370154 333100 370156
rect 286041 370152 333100 370154
rect 286041 370096 286046 370152
rect 286102 370096 300122 370152
rect 300178 370096 333100 370152
rect 286041 370094 333100 370096
rect 286041 370091 286107 370094
rect 300117 370091 300183 370094
rect 333094 370092 333100 370094
rect 333164 370092 333170 370156
rect 224217 370018 224283 370021
rect 284477 370018 284543 370021
rect 284845 370018 284911 370021
rect 331806 370018 331812 370020
rect 224217 370016 331812 370018
rect 224217 369960 224222 370016
rect 224278 369960 284482 370016
rect 284538 369960 284850 370016
rect 284906 369960 331812 370016
rect 224217 369958 331812 369960
rect 224217 369955 224283 369958
rect 284477 369955 284543 369958
rect 284845 369955 284911 369958
rect 331806 369956 331812 369958
rect 331876 369956 331882 370020
rect 282126 369820 282132 369884
rect 282196 369882 282202 369884
rect 302739 369882 302805 369885
rect 282196 369880 302805 369882
rect 282196 369824 302744 369880
rect 302800 369824 302805 369880
rect 282196 369822 302805 369824
rect 282196 369820 282202 369822
rect 302739 369819 302805 369822
rect 310697 369882 310763 369885
rect 311571 369882 311637 369885
rect 315849 369882 315915 369885
rect 310697 369880 311637 369882
rect 310697 369824 310702 369880
rect 310758 369824 311576 369880
rect 311632 369824 311637 369880
rect 310697 369822 311637 369824
rect 310697 369819 310763 369822
rect 311571 369819 311637 369822
rect 315806 369880 315915 369882
rect 315806 369824 315854 369880
rect 315910 369824 315915 369880
rect 315806 369819 315915 369824
rect 280429 369746 280495 369749
rect 288019 369746 288085 369749
rect 312077 369746 312143 369749
rect 280429 369744 288085 369746
rect 280429 369688 280434 369744
rect 280490 369688 288024 369744
rect 288080 369688 288085 369744
rect 280429 369686 288085 369688
rect 280429 369683 280495 369686
rect 288019 369683 288085 369686
rect 292530 369744 312143 369746
rect 292530 369688 312082 369744
rect 312138 369688 312143 369744
rect 292530 369686 312143 369688
rect 285075 369610 285141 369613
rect 287283 369612 287349 369613
rect 285622 369610 285628 369612
rect 285075 369608 285628 369610
rect 285075 369552 285080 369608
rect 285136 369552 285628 369608
rect 285075 369550 285628 369552
rect 285075 369547 285141 369550
rect 285622 369548 285628 369550
rect 285692 369548 285698 369612
rect 287278 369610 287284 369612
rect 287192 369550 287284 369610
rect 287278 369548 287284 369550
rect 287348 369548 287354 369612
rect 287283 369547 287349 369548
rect 276013 369474 276079 369477
rect 290089 369474 290155 369477
rect 276013 369472 290155 369474
rect 276013 369416 276018 369472
rect 276074 369416 290094 369472
rect 290150 369416 290155 369472
rect 276013 369414 290155 369416
rect 276013 369411 276079 369414
rect 290089 369411 290155 369414
rect 228357 369338 228423 369341
rect 279918 369338 279924 369340
rect 228357 369336 279924 369338
rect 228357 369280 228362 369336
rect 228418 369280 279924 369336
rect 228357 369278 279924 369280
rect 228357 369275 228423 369278
rect 279918 369276 279924 369278
rect 279988 369338 279994 369340
rect 280429 369338 280495 369341
rect 285811 369338 285877 369341
rect 287283 369340 287349 369341
rect 287278 369338 287284 369340
rect 279988 369336 280495 369338
rect 279988 369280 280434 369336
rect 280490 369280 280495 369336
rect 279988 369278 280495 369280
rect 279988 369276 279994 369278
rect 280429 369275 280495 369278
rect 282870 369336 285877 369338
rect 282870 369280 285816 369336
rect 285872 369280 285877 369336
rect 282870 369278 285877 369280
rect 287192 369278 287284 369338
rect 225597 369202 225663 369205
rect 278630 369202 278636 369204
rect 225597 369200 278636 369202
rect 225597 369144 225602 369200
rect 225658 369144 278636 369200
rect 225597 369142 278636 369144
rect 225597 369139 225663 369142
rect 278630 369140 278636 369142
rect 278700 369202 278706 369204
rect 281390 369202 281396 369204
rect 278700 369142 281396 369202
rect 278700 369140 278706 369142
rect 281390 369140 281396 369142
rect 281460 369202 281466 369204
rect 282870 369202 282930 369278
rect 285811 369275 285877 369278
rect 287278 369276 287284 369278
rect 287348 369276 287354 369340
rect 287283 369275 287349 369276
rect 281460 369142 282930 369202
rect 281460 369140 281466 369142
rect 251817 369066 251883 369069
rect 292530 369066 292590 369686
rect 312077 369683 312143 369686
rect 315430 369684 315436 369748
rect 315500 369746 315506 369748
rect 315806 369746 315866 369819
rect 315500 369686 315866 369746
rect 315500 369684 315506 369686
rect 311014 369548 311020 369612
rect 311084 369610 311090 369612
rect 311801 369610 311867 369613
rect 311084 369608 311867 369610
rect 311084 369552 311806 369608
rect 311862 369552 311867 369608
rect 311084 369550 311867 369552
rect 311084 369548 311090 369550
rect 311801 369547 311867 369550
rect 313774 369548 313780 369612
rect 313844 369610 313850 369612
rect 314377 369610 314443 369613
rect 313844 369608 314443 369610
rect 313844 369552 314382 369608
rect 314438 369552 314443 369608
rect 313844 369550 314443 369552
rect 313844 369548 313850 369550
rect 314377 369547 314443 369550
rect 319294 369548 319300 369612
rect 319364 369610 319370 369612
rect 319897 369610 319963 369613
rect 319364 369608 319963 369610
rect 319364 369552 319902 369608
rect 319958 369552 319963 369608
rect 319364 369550 319963 369552
rect 319364 369548 319370 369550
rect 319897 369547 319963 369550
rect 320950 369548 320956 369612
rect 321020 369610 321026 369612
rect 321369 369610 321435 369613
rect 321020 369608 321435 369610
rect 321020 369552 321374 369608
rect 321430 369552 321435 369608
rect 321020 369550 321435 369552
rect 321020 369548 321026 369550
rect 321369 369547 321435 369550
rect 301446 369412 301452 369476
rect 301516 369474 301522 369476
rect 302141 369474 302207 369477
rect 301516 369472 302207 369474
rect 301516 369416 302146 369472
rect 302202 369416 302207 369472
rect 301516 369414 302207 369416
rect 301516 369412 301522 369414
rect 302141 369411 302207 369414
rect 302734 369412 302740 369476
rect 302804 369474 302810 369476
rect 303337 369474 303403 369477
rect 302804 369472 303403 369474
rect 302804 369416 303342 369472
rect 303398 369416 303403 369472
rect 302804 369414 303403 369416
rect 302804 369412 302810 369414
rect 303337 369411 303403 369414
rect 311198 369412 311204 369476
rect 311268 369474 311274 369476
rect 311433 369474 311499 369477
rect 311268 369472 311499 369474
rect 311268 369416 311438 369472
rect 311494 369416 311499 369472
rect 311268 369414 311499 369416
rect 311268 369412 311274 369414
rect 311433 369411 311499 369414
rect 312486 369412 312492 369476
rect 312556 369474 312562 369476
rect 313181 369474 313247 369477
rect 312556 369472 313247 369474
rect 312556 369416 313186 369472
rect 313242 369416 313247 369472
rect 312556 369414 313247 369416
rect 312556 369412 312562 369414
rect 313181 369411 313247 369414
rect 313590 369412 313596 369476
rect 313660 369474 313666 369476
rect 314285 369474 314351 369477
rect 313660 369472 314351 369474
rect 313660 369416 314290 369472
rect 314346 369416 314351 369472
rect 313660 369414 314351 369416
rect 313660 369412 313666 369414
rect 314285 369411 314351 369414
rect 318006 369412 318012 369476
rect 318076 369474 318082 369476
rect 318701 369474 318767 369477
rect 318076 369472 318767 369474
rect 318076 369416 318706 369472
rect 318762 369416 318767 369472
rect 318076 369414 318767 369416
rect 318076 369412 318082 369414
rect 318701 369411 318767 369414
rect 319662 369412 319668 369476
rect 319732 369474 319738 369476
rect 319805 369474 319871 369477
rect 319732 369472 319871 369474
rect 319732 369416 319810 369472
rect 319866 369416 319871 369472
rect 319732 369414 319871 369416
rect 319732 369412 319738 369414
rect 319805 369411 319871 369414
rect 321134 369412 321140 369476
rect 321204 369474 321210 369476
rect 321277 369474 321343 369477
rect 321204 369472 321343 369474
rect 321204 369416 321282 369472
rect 321338 369416 321343 369472
rect 321204 369414 321343 369416
rect 321204 369412 321210 369414
rect 321277 369411 321343 369414
rect 308995 369336 309061 369341
rect 310099 369340 310165 369341
rect 310094 369338 310100 369340
rect 308995 369280 309000 369336
rect 309056 369280 309061 369336
rect 308995 369275 309061 369280
rect 310008 369278 310100 369338
rect 310094 369276 310100 369278
rect 310164 369276 310170 369340
rect 310099 369275 310165 369276
rect 251817 369064 292590 369066
rect 251817 369008 251822 369064
rect 251878 369008 292590 369064
rect 251817 369006 292590 369008
rect 251817 369003 251883 369006
rect 248413 368930 248479 368933
rect 308998 368930 309058 369275
rect 248413 368928 309058 368930
rect 248413 368872 248418 368928
rect 248474 368872 309058 368928
rect 248413 368870 309058 368872
rect 248413 368867 248479 368870
rect 285622 368732 285628 368796
rect 285692 368794 285698 368796
rect 334617 368794 334683 368797
rect 285692 368792 334683 368794
rect 285692 368736 334622 368792
rect 334678 368736 334683 368792
rect 285692 368734 334683 368736
rect 285692 368732 285698 368734
rect 334617 368731 334683 368734
rect 229921 368658 229987 368661
rect 276013 368658 276079 368661
rect 276381 368658 276447 368661
rect 229921 368656 276447 368658
rect 229921 368600 229926 368656
rect 229982 368600 276018 368656
rect 276074 368600 276386 368656
rect 276442 368600 276447 368656
rect 229921 368598 276447 368600
rect 229921 368595 229987 368598
rect 276013 368595 276079 368598
rect 276381 368595 276447 368598
rect 287278 368596 287284 368660
rect 287348 368658 287354 368660
rect 339401 368658 339467 368661
rect 341517 368658 341583 368661
rect 287348 368656 341583 368658
rect 287348 368600 339406 368656
rect 339462 368600 341522 368656
rect 341578 368600 341583 368656
rect 287348 368598 341583 368600
rect 287348 368596 287354 368598
rect 339401 368595 339467 368598
rect 341517 368595 341583 368598
rect 250437 368386 250503 368389
rect 310094 368386 310100 368388
rect 250437 368384 310100 368386
rect 250437 368328 250442 368384
rect 250498 368328 310100 368384
rect 250437 368326 310100 368328
rect 250437 368323 250503 368326
rect 310094 368324 310100 368326
rect 310164 368386 310170 368388
rect 334985 368386 335051 368389
rect 310164 368384 335051 368386
rect 310164 368328 334990 368384
rect 335046 368328 335051 368384
rect 310164 368326 335051 368328
rect 310164 368324 310170 368326
rect 334985 368323 335051 368326
rect 328361 366482 328427 366485
rect 580257 366482 580323 366485
rect 328361 366480 580323 366482
rect 328361 366424 328366 366480
rect 328422 366424 580262 366480
rect 580318 366424 580323 366480
rect 328361 366422 580323 366424
rect 328361 366419 328427 366422
rect 580257 366419 580323 366422
rect 324262 366284 324268 366348
rect 324332 366346 324338 366348
rect 580533 366346 580599 366349
rect 324332 366344 580599 366346
rect 324332 366288 580538 366344
rect 580594 366288 580599 366344
rect 324332 366286 580599 366288
rect 324332 366284 324338 366286
rect 580533 366283 580599 366286
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 323158 364924 323164 364988
rect 323228 364986 323234 364988
rect 580441 364986 580507 364989
rect 323228 364984 580507 364986
rect 323228 364928 580446 364984
rect 580502 364928 580507 364984
rect 583520 364972 584960 365062
rect 323228 364926 580507 364928
rect 323228 364924 323234 364926
rect 580441 364923 580507 364926
rect 250437 363626 250503 363629
rect 281022 363626 281028 363628
rect 250437 363624 281028 363626
rect 250437 363568 250442 363624
rect 250498 363568 281028 363624
rect 250437 363566 281028 363568
rect 250437 363563 250503 363566
rect 281022 363564 281028 363566
rect 281092 363564 281098 363628
rect 251909 362266 251975 362269
rect 280838 362266 280844 362268
rect 251909 362264 280844 362266
rect 251909 362208 251914 362264
rect 251970 362208 280844 362264
rect 251909 362206 280844 362208
rect 251909 362203 251975 362206
rect 280838 362204 280844 362206
rect 280908 362204 280914 362268
rect 243537 360906 243603 360909
rect 282269 360906 282335 360909
rect 243537 360904 282335 360906
rect 243537 360848 243542 360904
rect 243598 360848 282274 360904
rect 282330 360848 282335 360904
rect 243537 360846 282335 360848
rect 243537 360843 243603 360846
rect 282269 360843 282335 360846
rect 277669 358866 277735 358869
rect 278446 358866 278452 358868
rect 277669 358864 278452 358866
rect 277669 358808 277674 358864
rect 277730 358808 278452 358864
rect 277669 358806 278452 358808
rect 277669 358803 277735 358806
rect 278446 358804 278452 358806
rect 278516 358804 278522 358868
rect -960 358458 480 358548
rect 3141 358458 3207 358461
rect -960 358456 3207 358458
rect -960 358400 3146 358456
rect 3202 358400 3207 358456
rect -960 358398 3207 358400
rect -960 358308 480 358398
rect 3141 358395 3207 358398
rect 247769 358050 247835 358053
rect 282310 358050 282316 358052
rect 247769 358048 282316 358050
rect 247769 357992 247774 358048
rect 247830 357992 282316 358048
rect 247769 357990 282316 357992
rect 247769 357987 247835 357990
rect 282310 357988 282316 357990
rect 282380 357988 282386 358052
rect 327809 358050 327875 358053
rect 350942 358050 350948 358052
rect 327809 358048 350948 358050
rect 327809 357992 327814 358048
rect 327870 357992 350948 358048
rect 327809 357990 350948 357992
rect 327809 357987 327875 357990
rect 350942 357988 350948 357990
rect 351012 357988 351018 358052
rect 280705 356826 280771 356829
rect 281257 356826 281323 356829
rect 280705 356824 281323 356826
rect 280705 356768 280710 356824
rect 280766 356768 281262 356824
rect 281318 356768 281323 356824
rect 280705 356766 281323 356768
rect 280705 356763 280771 356766
rect 281257 356763 281323 356766
rect 323710 356628 323716 356692
rect 323780 356690 323786 356692
rect 383929 356690 383995 356693
rect 323780 356688 383995 356690
rect 323780 356632 383934 356688
rect 383990 356632 383995 356688
rect 323780 356630 383995 356632
rect 323780 356628 323786 356630
rect 383929 356627 383995 356630
rect 246389 353970 246455 353973
rect 282177 353970 282243 353973
rect 246389 353968 282243 353970
rect 246389 353912 246394 353968
rect 246450 353912 282182 353968
rect 282238 353912 282243 353968
rect 246389 353910 282243 353912
rect 246389 353907 246455 353910
rect 282177 353907 282243 353910
rect 580717 351930 580783 351933
rect 583520 351930 584960 352020
rect 580717 351928 584960 351930
rect 580717 351872 580722 351928
rect 580778 351872 584960 351928
rect 580717 351870 584960 351872
rect 580717 351867 580783 351870
rect 583520 351780 584960 351870
rect 280705 345810 280771 345813
rect 281073 345810 281139 345813
rect 280705 345808 281139 345810
rect 280705 345752 280710 345808
rect 280766 345752 281078 345808
rect 281134 345752 281139 345808
rect 280705 345750 281139 345752
rect 280705 345747 280771 345750
rect 281073 345747 281139 345750
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 323894 342892 323900 342956
rect 323964 342954 323970 342956
rect 382457 342954 382523 342957
rect 323964 342952 382523 342954
rect 323964 342896 382462 342952
rect 382518 342896 382523 342952
rect 323964 342894 382523 342896
rect 323964 342892 323970 342894
rect 382457 342891 382523 342894
rect 327901 341594 327967 341597
rect 374453 341594 374519 341597
rect 327901 341592 374519 341594
rect 327901 341536 327906 341592
rect 327962 341536 374458 341592
rect 374514 341536 374519 341592
rect 327901 341534 374519 341536
rect 327901 341531 327967 341534
rect 374453 341531 374519 341534
rect 325366 341396 325372 341460
rect 325436 341458 325442 341460
rect 385309 341458 385375 341461
rect 325436 341456 385375 341458
rect 325436 341400 385314 341456
rect 385370 341400 385375 341456
rect 325436 341398 385375 341400
rect 325436 341396 325442 341398
rect 385309 341395 385375 341398
rect 324630 340036 324636 340100
rect 324700 340098 324706 340100
rect 383745 340098 383811 340101
rect 324700 340096 383811 340098
rect 324700 340040 383750 340096
rect 383806 340040 383811 340096
rect 324700 340038 383811 340040
rect 324700 340036 324706 340038
rect 383745 340035 383811 340038
rect 583520 338452 584960 338692
rect 376518 338132 376524 338196
rect 376588 338194 376594 338196
rect 427813 338194 427879 338197
rect 376588 338192 427879 338194
rect 376588 338136 427818 338192
rect 427874 338136 427879 338192
rect 376588 338134 427879 338136
rect 376588 338132 376594 338134
rect 427813 338131 427879 338134
rect 380750 335412 380756 335476
rect 380820 335474 380826 335476
rect 513373 335474 513439 335477
rect 380820 335472 513439 335474
rect 380820 335416 513378 335472
rect 513434 335416 513439 335472
rect 380820 335414 513439 335416
rect 380820 335412 380826 335414
rect 513373 335411 513439 335414
rect 340505 334658 340571 334661
rect 380750 334658 380756 334660
rect 340505 334656 380756 334658
rect 340505 334600 340510 334656
rect 340566 334600 380756 334656
rect 340505 334598 380756 334600
rect 340505 334595 340571 334598
rect 380750 334596 380756 334598
rect 380820 334596 380826 334660
rect 327441 333298 327507 333301
rect 386873 333298 386939 333301
rect 327441 333296 386939 333298
rect 327441 333240 327446 333296
rect 327502 333240 386878 333296
rect 386934 333240 386939 333296
rect 327441 333238 386939 333240
rect 327441 333235 327507 333238
rect 386873 333235 386939 333238
rect -960 332196 480 332436
rect 329230 330516 329236 330580
rect 329300 330578 329306 330580
rect 379697 330578 379763 330581
rect 329300 330576 379763 330578
rect 329300 330520 379702 330576
rect 379758 330520 379763 330576
rect 329300 330518 379763 330520
rect 329300 330516 329306 330518
rect 379697 330515 379763 330518
rect 327533 330442 327599 330445
rect 386781 330442 386847 330445
rect 327533 330440 386847 330442
rect 327533 330384 327538 330440
rect 327594 330384 386786 330440
rect 386842 330384 386847 330440
rect 327533 330382 386847 330384
rect 327533 330379 327599 330382
rect 386781 330379 386847 330382
rect 327993 327722 328059 327725
rect 386689 327722 386755 327725
rect 327993 327720 386755 327722
rect 327993 327664 327998 327720
rect 328054 327664 386694 327720
rect 386750 327664 386755 327720
rect 327993 327662 386755 327664
rect 327993 327659 328059 327662
rect 386689 327659 386755 327662
rect 325366 327116 325372 327180
rect 325436 327178 325442 327180
rect 331213 327178 331279 327181
rect 325436 327176 331279 327178
rect 325436 327120 331218 327176
rect 331274 327120 331279 327176
rect 325436 327118 331279 327120
rect 325436 327116 325442 327118
rect 331213 327115 331279 327118
rect 338614 326300 338620 326364
rect 338684 326362 338690 326364
rect 380893 326362 380959 326365
rect 338684 326360 380959 326362
rect 338684 326304 380898 326360
rect 380954 326304 380959 326360
rect 338684 326302 380959 326304
rect 338684 326300 338690 326302
rect 380893 326299 380959 326302
rect 342345 325274 342411 325277
rect 370078 325274 370084 325276
rect 342345 325272 370084 325274
rect 342345 325216 342350 325272
rect 342406 325216 370084 325272
rect 342345 325214 370084 325216
rect 342345 325211 342411 325214
rect 370078 325212 370084 325214
rect 370148 325212 370154 325276
rect 580717 325274 580783 325277
rect 583520 325274 584960 325364
rect 580717 325272 584960 325274
rect 580717 325216 580722 325272
rect 580778 325216 584960 325272
rect 580717 325214 584960 325216
rect 580717 325211 580783 325214
rect 337929 325138 337995 325141
rect 378358 325138 378364 325140
rect 337929 325136 378364 325138
rect 337929 325080 337934 325136
rect 337990 325080 378364 325136
rect 337929 325078 378364 325080
rect 337929 325075 337995 325078
rect 378358 325076 378364 325078
rect 378428 325076 378434 325140
rect 583520 325124 584960 325214
rect 340873 325002 340939 325005
rect 382222 325002 382228 325004
rect 335310 325000 382228 325002
rect 335310 324944 340878 325000
rect 340934 324944 382228 325000
rect 335310 324942 382228 324944
rect 323526 324396 323532 324460
rect 323596 324458 323602 324460
rect 335310 324458 335370 324942
rect 340873 324939 340939 324942
rect 382222 324940 382228 324942
rect 382292 324940 382298 325004
rect 323596 324398 335370 324458
rect 323596 324396 323602 324398
rect 330293 323778 330359 323781
rect 385769 323778 385835 323781
rect 330293 323776 385835 323778
rect 330293 323720 330298 323776
rect 330354 323720 385774 323776
rect 385830 323720 385835 323776
rect 330293 323718 385835 323720
rect 330293 323715 330359 323718
rect 385769 323715 385835 323718
rect 230013 323642 230079 323645
rect 276606 323642 276612 323644
rect 230013 323640 276612 323642
rect 230013 323584 230018 323640
rect 230074 323584 276612 323640
rect 230013 323582 276612 323584
rect 230013 323579 230079 323582
rect 276606 323580 276612 323582
rect 276676 323580 276682 323644
rect 324078 323580 324084 323644
rect 324148 323642 324154 323644
rect 384941 323642 385007 323645
rect 324148 323640 385007 323642
rect 324148 323584 384946 323640
rect 385002 323584 385007 323640
rect 324148 323582 385007 323584
rect 324148 323580 324154 323582
rect 384941 323579 385007 323582
rect 327758 322900 327764 322964
rect 327828 322962 327834 322964
rect 329833 322962 329899 322965
rect 330293 322962 330359 322965
rect 327828 322960 330359 322962
rect 327828 322904 329838 322960
rect 329894 322904 330298 322960
rect 330354 322904 330359 322960
rect 327828 322902 330359 322904
rect 327828 322900 327834 322902
rect 329833 322899 329899 322902
rect 330293 322899 330359 322902
rect 326654 322220 326660 322284
rect 326724 322282 326730 322284
rect 330334 322282 330340 322284
rect 326724 322222 330340 322282
rect 326724 322220 326730 322222
rect 330334 322220 330340 322222
rect 330404 322282 330410 322284
rect 385166 322282 385172 322284
rect 330404 322222 385172 322282
rect 330404 322220 330410 322222
rect 385166 322220 385172 322222
rect 385236 322220 385242 322284
rect 324446 322084 324452 322148
rect 324516 322146 324522 322148
rect 385861 322146 385927 322149
rect 324516 322144 385927 322146
rect 324516 322088 385866 322144
rect 385922 322088 385927 322144
rect 324516 322086 385927 322088
rect 324516 322084 324522 322086
rect 385861 322083 385927 322086
rect 320766 321948 320772 322012
rect 320836 322010 320842 322012
rect 349613 322010 349679 322013
rect 320836 322008 349679 322010
rect 320836 321952 349618 322008
rect 349674 321952 349679 322008
rect 320836 321950 349679 321952
rect 320836 321948 320842 321950
rect 349613 321947 349679 321950
rect 308806 321812 308812 321876
rect 308876 321874 308882 321876
rect 339493 321874 339559 321877
rect 339953 321874 340019 321877
rect 308876 321872 340019 321874
rect 308876 321816 339498 321872
rect 339554 321816 339958 321872
rect 340014 321816 340019 321872
rect 308876 321814 340019 321816
rect 308876 321812 308882 321814
rect 339493 321811 339559 321814
rect 339953 321811 340019 321814
rect 202781 321602 202847 321605
rect 327441 321604 327507 321605
rect 283966 321602 283972 321604
rect 202781 321600 283972 321602
rect 202781 321544 202786 321600
rect 202842 321544 283972 321600
rect 202781 321542 283972 321544
rect 202781 321539 202847 321542
rect 283966 321540 283972 321542
rect 284036 321540 284042 321604
rect 327390 321602 327396 321604
rect 327350 321542 327396 321602
rect 327460 321600 327507 321604
rect 327502 321544 327507 321600
rect 327390 321540 327396 321542
rect 327460 321540 327507 321544
rect 327441 321539 327507 321540
rect 327625 321602 327691 321605
rect 336733 321602 336799 321605
rect 386597 321602 386663 321605
rect 387057 321602 387123 321605
rect 327625 321600 387123 321602
rect 327625 321544 327630 321600
rect 327686 321544 336738 321600
rect 336794 321544 386602 321600
rect 386658 321544 387062 321600
rect 387118 321544 387123 321600
rect 327625 321542 387123 321544
rect 327625 321539 327691 321542
rect 336733 321539 336799 321542
rect 386597 321539 386663 321542
rect 387057 321539 387123 321542
rect 272793 321466 272859 321469
rect 272977 321466 273043 321469
rect 278037 321466 278103 321469
rect 272793 321464 278103 321466
rect 272793 321408 272798 321464
rect 272854 321408 272982 321464
rect 273038 321408 278042 321464
rect 278098 321408 278103 321464
rect 272793 321406 278103 321408
rect 272793 321403 272859 321406
rect 272977 321403 273043 321406
rect 278037 321403 278103 321406
rect 320582 321404 320588 321468
rect 320652 321466 320658 321468
rect 328361 321466 328427 321469
rect 320652 321464 328427 321466
rect 320652 321408 328366 321464
rect 328422 321408 328427 321464
rect 320652 321406 328427 321408
rect 320652 321404 320658 321406
rect 328361 321403 328427 321406
rect 282269 321330 282335 321333
rect 294454 321330 294460 321332
rect 282269 321328 294460 321330
rect 282269 321272 282274 321328
rect 282330 321272 294460 321328
rect 282269 321270 294460 321272
rect 282269 321267 282335 321270
rect 294454 321268 294460 321270
rect 294524 321268 294530 321332
rect 320950 321268 320956 321332
rect 321020 321330 321026 321332
rect 321502 321330 321508 321332
rect 321020 321270 321508 321330
rect 321020 321268 321026 321270
rect 321502 321268 321508 321270
rect 321572 321268 321578 321332
rect 322974 321268 322980 321332
rect 323044 321330 323050 321332
rect 330201 321330 330267 321333
rect 330937 321330 331003 321333
rect 323044 321328 331003 321330
rect 323044 321272 330206 321328
rect 330262 321272 330942 321328
rect 330998 321272 331003 321328
rect 323044 321270 331003 321272
rect 323044 321268 323050 321270
rect 330201 321267 330267 321270
rect 330937 321267 331003 321270
rect 225689 321194 225755 321197
rect 279366 321194 279372 321196
rect 225689 321192 279372 321194
rect 225689 321136 225694 321192
rect 225750 321136 279372 321192
rect 225689 321134 279372 321136
rect 225689 321131 225755 321134
rect 279366 321132 279372 321134
rect 279436 321132 279442 321196
rect 294270 321132 294276 321196
rect 294340 321194 294346 321196
rect 295190 321194 295196 321196
rect 294340 321134 295196 321194
rect 294340 321132 294346 321134
rect 295190 321132 295196 321134
rect 295260 321132 295266 321196
rect 301446 321132 301452 321196
rect 301516 321194 301522 321196
rect 306966 321194 306972 321196
rect 301516 321134 306972 321194
rect 301516 321132 301522 321134
rect 306966 321132 306972 321134
rect 307036 321132 307042 321196
rect 318926 321132 318932 321196
rect 318996 321194 319002 321196
rect 327901 321194 327967 321197
rect 318996 321192 327967 321194
rect 318996 321136 327906 321192
rect 327962 321136 327967 321192
rect 318996 321134 327967 321136
rect 318996 321132 319002 321134
rect 327901 321131 327967 321134
rect 328361 321194 328427 321197
rect 340045 321194 340111 321197
rect 328361 321192 340111 321194
rect 328361 321136 328366 321192
rect 328422 321136 340050 321192
rect 340106 321136 340111 321192
rect 328361 321134 340111 321136
rect 328361 321131 328427 321134
rect 340045 321131 340111 321134
rect 217961 321058 218027 321061
rect 272793 321058 272859 321061
rect 217961 321056 272859 321058
rect 217961 321000 217966 321056
rect 218022 321000 272798 321056
rect 272854 321000 272859 321056
rect 217961 320998 272859 321000
rect 217961 320995 218027 320998
rect 272793 320995 272859 320998
rect 273713 321058 273779 321061
rect 278313 321058 278379 321061
rect 303286 321058 303292 321060
rect 273713 321056 303292 321058
rect 273713 321000 273718 321056
rect 273774 321000 278318 321056
rect 278374 321000 303292 321056
rect 273713 320998 303292 321000
rect 273713 320995 273779 320998
rect 278313 320995 278379 320998
rect 303286 320996 303292 320998
rect 303356 320996 303362 321060
rect 321318 320996 321324 321060
rect 321388 321058 321394 321060
rect 327809 321058 327875 321061
rect 321388 321056 327875 321058
rect 321388 321000 327814 321056
rect 327870 321000 327875 321056
rect 321388 320998 327875 321000
rect 321388 320996 321394 320998
rect 327809 320995 327875 320998
rect 338205 321058 338271 321061
rect 378174 321058 378180 321060
rect 338205 321056 378180 321058
rect 338205 321000 338210 321056
rect 338266 321000 378180 321056
rect 338205 320998 378180 321000
rect 338205 320995 338271 320998
rect 378174 320996 378180 320998
rect 378244 320996 378250 321060
rect 206921 320922 206987 320925
rect 271413 320922 271479 320925
rect 206921 320920 285322 320922
rect 206921 320864 206926 320920
rect 206982 320864 271418 320920
rect 271474 320864 285322 320920
rect 206921 320862 285322 320864
rect 206921 320859 206987 320862
rect 271413 320859 271479 320862
rect 210969 320786 211035 320789
rect 275553 320786 275619 320789
rect 282269 320786 282335 320789
rect 210969 320784 275619 320786
rect 210969 320728 210974 320784
rect 211030 320728 275558 320784
rect 275614 320728 275619 320784
rect 210969 320726 275619 320728
rect 210969 320723 211035 320726
rect 275553 320723 275619 320726
rect 277902 320784 282335 320786
rect 277902 320728 282274 320784
rect 282330 320728 282335 320784
rect 277902 320726 282335 320728
rect 275461 320650 275527 320653
rect 277902 320650 277962 320726
rect 282269 320723 282335 320726
rect 283235 320786 283301 320789
rect 283782 320786 283788 320788
rect 283235 320784 283788 320786
rect 283235 320728 283240 320784
rect 283296 320728 283788 320784
rect 283235 320726 283788 320728
rect 283235 320723 283301 320726
rect 283782 320724 283788 320726
rect 283852 320724 283858 320788
rect 283966 320724 283972 320788
rect 284036 320786 284042 320788
rect 284247 320786 284313 320789
rect 284036 320784 284313 320786
rect 284036 320728 284252 320784
rect 284308 320728 284313 320784
rect 284036 320726 284313 320728
rect 285262 320786 285322 320862
rect 287094 320860 287100 320924
rect 287164 320922 287170 320924
rect 346117 320922 346183 320925
rect 287164 320920 346183 320922
rect 287164 320864 346122 320920
rect 346178 320864 346183 320920
rect 287164 320862 346183 320864
rect 287164 320860 287170 320862
rect 346117 320859 346183 320862
rect 287467 320786 287533 320789
rect 288203 320788 288269 320789
rect 288198 320786 288204 320788
rect 285262 320784 287533 320786
rect 285262 320728 287472 320784
rect 287528 320728 287533 320784
rect 285262 320726 287533 320728
rect 288112 320726 288204 320786
rect 284036 320724 284042 320726
rect 284247 320723 284313 320726
rect 287467 320723 287533 320726
rect 288198 320724 288204 320726
rect 288268 320724 288274 320788
rect 290595 320786 290661 320789
rect 290958 320786 290964 320788
rect 290595 320784 290964 320786
rect 290595 320728 290600 320784
rect 290656 320728 290964 320784
rect 290595 320726 290964 320728
rect 288203 320723 288269 320724
rect 290595 320723 290661 320726
rect 290958 320724 290964 320726
rect 291028 320724 291034 320788
rect 291147 320786 291213 320789
rect 291694 320786 291700 320788
rect 291147 320784 291700 320786
rect 291147 320728 291152 320784
rect 291208 320728 291700 320784
rect 291147 320726 291700 320728
rect 291147 320723 291213 320726
rect 291694 320724 291700 320726
rect 291764 320724 291770 320788
rect 291883 320786 291949 320789
rect 292062 320786 292068 320788
rect 291883 320784 292068 320786
rect 291883 320728 291888 320784
rect 291944 320728 292068 320784
rect 291883 320726 292068 320728
rect 291883 320723 291949 320726
rect 292062 320724 292068 320726
rect 292132 320786 292138 320788
rect 292430 320786 292436 320788
rect 292132 320726 292436 320786
rect 292132 320724 292138 320726
rect 292430 320724 292436 320726
rect 292500 320724 292506 320788
rect 292619 320786 292685 320789
rect 295926 320786 295932 320788
rect 292619 320784 295932 320786
rect 292619 320728 292624 320784
rect 292680 320728 295932 320784
rect 292619 320726 295932 320728
rect 292619 320723 292685 320726
rect 295926 320724 295932 320726
rect 295996 320724 296002 320788
rect 296294 320786 296300 320788
rect 296164 320726 296300 320786
rect 275461 320648 277962 320650
rect 275461 320592 275466 320648
rect 275522 320592 277962 320648
rect 275461 320590 277962 320592
rect 278037 320650 278103 320653
rect 283327 320650 283393 320653
rect 283603 320652 283669 320653
rect 283598 320650 283604 320652
rect 278037 320648 283393 320650
rect 278037 320592 278042 320648
rect 278098 320592 283332 320648
rect 283388 320592 283393 320648
rect 278037 320590 283393 320592
rect 283512 320590 283604 320650
rect 275461 320587 275527 320590
rect 278037 320587 278103 320590
rect 283327 320587 283393 320590
rect 283598 320588 283604 320590
rect 283668 320588 283674 320652
rect 283966 320588 283972 320652
rect 284036 320650 284042 320652
rect 286179 320650 286245 320653
rect 284036 320648 286245 320650
rect 284036 320592 286184 320648
rect 286240 320592 286245 320648
rect 284036 320590 286245 320592
rect 284036 320588 284042 320590
rect 283603 320587 283669 320588
rect 286179 320587 286245 320590
rect 286358 320588 286364 320652
rect 286428 320650 286434 320652
rect 286428 320590 295258 320650
rect 286428 320588 286434 320590
rect 275553 320514 275619 320517
rect 281625 320514 281691 320517
rect 275553 320512 281691 320514
rect 275553 320456 275558 320512
rect 275614 320456 281630 320512
rect 281686 320456 281691 320512
rect 275553 320454 281691 320456
rect 275553 320451 275619 320454
rect 281625 320451 281691 320454
rect 282269 320514 282335 320517
rect 282867 320514 282933 320517
rect 282269 320512 282933 320514
rect 282269 320456 282274 320512
rect 282330 320456 282872 320512
rect 282928 320456 282933 320512
rect 282269 320454 282933 320456
rect 282269 320451 282335 320454
rect 282867 320451 282933 320454
rect 283414 320452 283420 320516
rect 283484 320514 283490 320516
rect 283971 320514 284037 320517
rect 285254 320514 285260 320516
rect 283484 320512 284037 320514
rect 283484 320456 283976 320512
rect 284032 320456 284037 320512
rect 283484 320454 284037 320456
rect 283484 320452 283490 320454
rect 283971 320451 284037 320454
rect 284710 320454 285260 320514
rect 270125 320378 270191 320381
rect 284339 320380 284405 320381
rect 283966 320378 283972 320380
rect 270125 320376 283972 320378
rect 270125 320320 270130 320376
rect 270186 320320 283972 320376
rect 270125 320318 283972 320320
rect 270125 320315 270191 320318
rect 283966 320316 283972 320318
rect 284036 320316 284042 320380
rect 284334 320378 284340 320380
rect 284212 320318 284340 320378
rect 284404 320378 284410 320380
rect 284710 320378 284770 320454
rect 285254 320452 285260 320454
rect 285324 320452 285330 320516
rect 285806 320452 285812 320516
rect 285876 320514 285882 320516
rect 286547 320514 286613 320517
rect 286910 320514 286916 320516
rect 285876 320512 286916 320514
rect 285876 320456 286552 320512
rect 286608 320456 286916 320512
rect 285876 320454 286916 320456
rect 285876 320452 285882 320454
rect 286547 320451 286613 320454
rect 286910 320452 286916 320454
rect 286980 320452 286986 320516
rect 288382 320452 288388 320516
rect 288452 320514 288458 320516
rect 288663 320514 288729 320517
rect 288452 320512 288729 320514
rect 288452 320456 288668 320512
rect 288724 320456 288729 320512
rect 288452 320454 288729 320456
rect 288452 320452 288458 320454
rect 288663 320451 288729 320454
rect 292062 320452 292068 320516
rect 292132 320514 292138 320516
rect 292343 320514 292409 320517
rect 292132 320512 292409 320514
rect 292132 320456 292348 320512
rect 292404 320456 292409 320512
rect 292132 320454 292409 320456
rect 292132 320452 292138 320454
rect 292343 320451 292409 320454
rect 292798 320452 292804 320516
rect 292868 320514 292874 320516
rect 293350 320514 293356 320516
rect 292868 320454 293356 320514
rect 292868 320452 292874 320454
rect 293350 320452 293356 320454
rect 293420 320514 293426 320516
rect 293723 320514 293789 320517
rect 293420 320512 293789 320514
rect 293420 320456 293728 320512
rect 293784 320456 293789 320512
rect 293420 320454 293789 320456
rect 293420 320452 293426 320454
rect 293723 320451 293789 320454
rect 293999 320514 294065 320517
rect 294270 320514 294276 320516
rect 293999 320512 294276 320514
rect 293999 320456 294004 320512
rect 294060 320456 294276 320512
rect 293999 320454 294276 320456
rect 293999 320451 294065 320454
rect 294270 320452 294276 320454
rect 294340 320452 294346 320516
rect 294638 320452 294644 320516
rect 294708 320514 294714 320516
rect 294827 320514 294893 320517
rect 294708 320512 294893 320514
rect 294708 320456 294832 320512
rect 294888 320456 294893 320512
rect 294708 320454 294893 320456
rect 295198 320514 295258 320590
rect 295558 320588 295564 320652
rect 295628 320650 295634 320652
rect 296164 320650 296224 320726
rect 296294 320724 296300 320726
rect 296364 320786 296370 320788
rect 296483 320786 296549 320789
rect 296364 320784 296549 320786
rect 296364 320728 296488 320784
rect 296544 320728 296549 320784
rect 296364 320726 296549 320728
rect 296364 320724 296370 320726
rect 296483 320723 296549 320726
rect 296662 320724 296668 320788
rect 296732 320786 296738 320788
rect 297311 320786 297377 320789
rect 297950 320786 297956 320788
rect 296732 320784 297956 320786
rect 296732 320728 297316 320784
rect 297372 320728 297956 320784
rect 296732 320726 297956 320728
rect 296732 320724 296738 320726
rect 297311 320723 297377 320726
rect 297950 320724 297956 320726
rect 298020 320724 298026 320788
rect 298139 320786 298205 320789
rect 299059 320788 299125 320789
rect 298502 320786 298508 320788
rect 298139 320784 298508 320786
rect 298139 320728 298144 320784
rect 298200 320728 298508 320784
rect 298139 320726 298508 320728
rect 298139 320723 298205 320726
rect 298502 320724 298508 320726
rect 298572 320724 298578 320788
rect 299054 320786 299060 320788
rect 298968 320726 299060 320786
rect 299054 320724 299060 320726
rect 299124 320724 299130 320788
rect 302550 320724 302556 320788
rect 302620 320786 302626 320788
rect 303383 320786 303449 320789
rect 302620 320784 303449 320786
rect 302620 320728 303388 320784
rect 303444 320728 303449 320784
rect 302620 320726 303449 320728
rect 302620 320724 302626 320726
rect 299059 320723 299125 320724
rect 303383 320723 303449 320726
rect 306695 320786 306761 320789
rect 308811 320788 308877 320789
rect 323531 320788 323597 320789
rect 324083 320788 324149 320789
rect 306966 320786 306972 320788
rect 306695 320784 306972 320786
rect 306695 320728 306700 320784
rect 306756 320728 306972 320784
rect 306695 320726 306972 320728
rect 306695 320723 306761 320726
rect 306966 320724 306972 320726
rect 307036 320724 307042 320788
rect 308806 320786 308812 320788
rect 308720 320726 308812 320786
rect 308806 320724 308812 320726
rect 308876 320724 308882 320788
rect 323526 320786 323532 320788
rect 311850 320726 323226 320786
rect 323440 320726 323532 320786
rect 308811 320723 308877 320724
rect 311850 320650 311910 320726
rect 295628 320590 296224 320650
rect 296486 320590 311910 320650
rect 295628 320588 295634 320590
rect 296486 320514 296546 320590
rect 312670 320588 312676 320652
rect 312740 320650 312746 320652
rect 313043 320650 313109 320653
rect 315803 320652 315869 320653
rect 312740 320648 313109 320650
rect 312740 320592 313048 320648
rect 313104 320592 313109 320648
rect 312740 320590 313109 320592
rect 312740 320588 312746 320590
rect 313043 320587 313109 320590
rect 314878 320588 314884 320652
rect 314948 320650 314954 320652
rect 315798 320650 315804 320652
rect 314948 320590 315804 320650
rect 314948 320588 314954 320590
rect 315798 320588 315804 320590
rect 315868 320588 315874 320652
rect 316902 320588 316908 320652
rect 316972 320650 316978 320652
rect 317091 320650 317157 320653
rect 316972 320648 317157 320650
rect 316972 320592 317096 320648
rect 317152 320592 317157 320648
rect 316972 320590 317157 320592
rect 316972 320588 316978 320590
rect 315803 320587 315869 320588
rect 317091 320587 317157 320590
rect 317454 320588 317460 320652
rect 317524 320650 317530 320652
rect 317643 320650 317709 320653
rect 318011 320652 318077 320653
rect 318195 320652 318261 320653
rect 318931 320652 318997 320653
rect 318006 320650 318012 320652
rect 317524 320648 317709 320650
rect 317524 320592 317648 320648
rect 317704 320592 317709 320648
rect 317524 320590 317709 320592
rect 317920 320590 318012 320650
rect 317524 320588 317530 320590
rect 317643 320587 317709 320590
rect 318006 320588 318012 320590
rect 318076 320588 318082 320652
rect 318190 320588 318196 320652
rect 318260 320650 318266 320652
rect 318926 320650 318932 320652
rect 318260 320590 318352 320650
rect 318840 320590 318932 320650
rect 318260 320588 318266 320590
rect 318926 320588 318932 320590
rect 318996 320588 319002 320652
rect 319207 320650 319273 320653
rect 321318 320650 321324 320652
rect 319207 320648 321324 320650
rect 319207 320592 319212 320648
rect 319268 320592 321324 320648
rect 319207 320590 321324 320592
rect 318011 320587 318077 320588
rect 318195 320587 318261 320588
rect 318931 320587 318997 320588
rect 319207 320587 319273 320590
rect 321318 320588 321324 320590
rect 321388 320588 321394 320652
rect 322974 320650 322980 320652
rect 321510 320590 322980 320650
rect 295198 320454 296546 320514
rect 294708 320452 294714 320454
rect 294827 320451 294893 320454
rect 296846 320452 296852 320516
rect 296916 320514 296922 320516
rect 297863 320514 297929 320517
rect 296916 320512 297929 320514
rect 296916 320456 297868 320512
rect 297924 320456 297929 320512
rect 296916 320454 297929 320456
rect 296916 320452 296922 320454
rect 297863 320451 297929 320454
rect 298318 320452 298324 320516
rect 298388 320514 298394 320516
rect 298599 320514 298665 320517
rect 298388 320512 298665 320514
rect 298388 320456 298604 320512
rect 298660 320456 298665 320512
rect 298388 320454 298665 320456
rect 298388 320452 298394 320454
rect 298599 320451 298665 320454
rect 298870 320452 298876 320516
rect 298940 320514 298946 320516
rect 302182 320514 302188 320516
rect 298940 320454 302188 320514
rect 298940 320452 298946 320454
rect 302182 320452 302188 320454
rect 302252 320452 302258 320516
rect 305310 320452 305316 320516
rect 305380 320514 305386 320516
rect 305591 320514 305657 320517
rect 306046 320514 306052 320516
rect 305380 320512 306052 320514
rect 305380 320456 305596 320512
rect 305652 320456 306052 320512
rect 305380 320454 306052 320456
rect 305380 320452 305386 320454
rect 305591 320451 305657 320454
rect 306046 320452 306052 320454
rect 306116 320452 306122 320516
rect 307702 320452 307708 320516
rect 307772 320514 307778 320516
rect 308351 320514 308417 320517
rect 307772 320512 308417 320514
rect 307772 320456 308356 320512
rect 308412 320456 308417 320512
rect 307772 320454 308417 320456
rect 307772 320452 307778 320454
rect 308351 320451 308417 320454
rect 310375 320514 310441 320517
rect 310830 320514 310836 320516
rect 310375 320512 310836 320514
rect 310375 320456 310380 320512
rect 310436 320456 310836 320512
rect 310375 320454 310836 320456
rect 310375 320451 310441 320454
rect 310830 320452 310836 320454
rect 310900 320452 310906 320516
rect 321510 320514 321570 320590
rect 322974 320588 322980 320590
rect 323044 320588 323050 320652
rect 323166 320650 323226 320726
rect 323526 320724 323532 320726
rect 323596 320724 323602 320788
rect 324078 320786 324084 320788
rect 323992 320726 324084 320786
rect 324078 320724 324084 320726
rect 324148 320724 324154 320788
rect 324359 320786 324425 320789
rect 324814 320786 324820 320788
rect 324359 320784 324820 320786
rect 324359 320728 324364 320784
rect 324420 320728 324820 320784
rect 324359 320726 324820 320728
rect 323531 320723 323597 320724
rect 324083 320723 324149 320724
rect 324359 320723 324425 320726
rect 324814 320724 324820 320726
rect 324884 320724 324890 320788
rect 325187 320786 325253 320789
rect 325366 320786 325372 320788
rect 325187 320784 325372 320786
rect 325187 320728 325192 320784
rect 325248 320728 325372 320784
rect 325187 320726 325372 320728
rect 325187 320723 325253 320726
rect 325366 320724 325372 320726
rect 325436 320724 325442 320788
rect 325739 320786 325805 320789
rect 326654 320786 326660 320788
rect 325739 320784 326660 320786
rect 325739 320728 325744 320784
rect 325800 320728 326660 320784
rect 325739 320726 326660 320728
rect 325739 320723 325805 320726
rect 326654 320724 326660 320726
rect 326724 320724 326730 320788
rect 327027 320786 327093 320789
rect 327625 320786 327691 320789
rect 345473 320786 345539 320789
rect 327027 320784 327691 320786
rect 327027 320728 327032 320784
rect 327088 320728 327630 320784
rect 327686 320728 327691 320784
rect 327027 320726 327691 320728
rect 327027 320723 327093 320726
rect 327625 320723 327691 320726
rect 331170 320784 345539 320786
rect 331170 320728 345478 320784
rect 345534 320728 345539 320784
rect 331170 320726 345539 320728
rect 331170 320650 331230 320726
rect 345473 320723 345539 320726
rect 323166 320590 331230 320650
rect 334525 320650 334591 320653
rect 338113 320650 338179 320653
rect 334525 320648 338179 320650
rect 334525 320592 334530 320648
rect 334586 320592 338118 320648
rect 338174 320592 338179 320648
rect 334525 320590 338179 320592
rect 334525 320587 334591 320590
rect 338113 320587 338179 320590
rect 322059 320516 322125 320517
rect 322054 320514 322060 320516
rect 311850 320454 321570 320514
rect 321968 320454 322060 320514
rect 284334 320316 284340 320318
rect 284404 320318 284770 320378
rect 284404 320316 284410 320318
rect 285070 320316 285076 320380
rect 285140 320378 285146 320380
rect 285443 320378 285509 320381
rect 285140 320376 285509 320378
rect 285140 320320 285448 320376
rect 285504 320320 285509 320376
rect 285140 320318 285509 320320
rect 285140 320316 285146 320318
rect 284339 320315 284405 320316
rect 285443 320315 285509 320318
rect 285719 320378 285785 320381
rect 286542 320378 286548 320380
rect 285719 320376 286548 320378
rect 285719 320320 285724 320376
rect 285780 320320 286548 320376
rect 285719 320318 286548 320320
rect 285719 320315 285785 320318
rect 286542 320316 286548 320318
rect 286612 320316 286618 320380
rect 287462 320316 287468 320380
rect 287532 320378 287538 320380
rect 287743 320378 287809 320381
rect 289491 320380 289557 320381
rect 287532 320376 287809 320378
rect 287532 320320 287748 320376
rect 287804 320320 287809 320376
rect 287532 320318 287809 320320
rect 287532 320316 287538 320318
rect 287743 320315 287809 320318
rect 288382 320316 288388 320380
rect 288452 320378 288458 320380
rect 289486 320378 289492 320380
rect 288452 320318 289492 320378
rect 288452 320316 288458 320318
rect 289486 320316 289492 320318
rect 289556 320316 289562 320380
rect 290043 320378 290109 320381
rect 290774 320378 290780 320380
rect 290043 320376 290780 320378
rect 290043 320320 290048 320376
rect 290104 320320 290780 320376
rect 290043 320318 290780 320320
rect 289491 320315 289557 320316
rect 290043 320315 290109 320318
rect 290774 320316 290780 320318
rect 290844 320316 290850 320380
rect 291699 320378 291765 320381
rect 292246 320378 292252 320380
rect 291699 320376 292252 320378
rect 291699 320320 291704 320376
rect 291760 320320 292252 320376
rect 291699 320318 292252 320320
rect 291699 320315 291765 320318
rect 292246 320316 292252 320318
rect 292316 320316 292322 320380
rect 292614 320316 292620 320380
rect 292684 320378 292690 320380
rect 294002 320378 294062 320451
rect 292684 320318 294062 320378
rect 292684 320316 292690 320318
rect 294454 320316 294460 320380
rect 294524 320378 294530 320380
rect 307891 320378 307957 320381
rect 309547 320380 309613 320381
rect 309542 320378 309548 320380
rect 294524 320376 307957 320378
rect 294524 320320 307896 320376
rect 307952 320320 307957 320376
rect 294524 320318 307957 320320
rect 309456 320318 309548 320378
rect 294524 320316 294530 320318
rect 307891 320315 307957 320318
rect 309542 320316 309548 320318
rect 309612 320316 309618 320380
rect 309910 320316 309916 320380
rect 309980 320378 309986 320380
rect 310099 320378 310165 320381
rect 310283 320380 310349 320381
rect 310651 320380 310717 320381
rect 311387 320380 311453 320381
rect 309980 320376 310165 320378
rect 309980 320320 310104 320376
rect 310160 320320 310165 320376
rect 309980 320318 310165 320320
rect 309980 320316 309986 320318
rect 309547 320315 309613 320316
rect 310099 320315 310165 320318
rect 310278 320316 310284 320380
rect 310348 320378 310354 320380
rect 310646 320378 310652 320380
rect 310348 320318 310440 320378
rect 310560 320318 310652 320378
rect 310348 320316 310354 320318
rect 310646 320316 310652 320318
rect 310716 320316 310722 320380
rect 311014 320316 311020 320380
rect 311084 320378 311090 320380
rect 311382 320378 311388 320380
rect 311084 320318 311388 320378
rect 311084 320316 311090 320318
rect 311382 320316 311388 320318
rect 311452 320316 311458 320380
rect 310283 320315 310349 320316
rect 310651 320315 310717 320316
rect 311387 320315 311453 320316
rect 275277 320242 275343 320245
rect 275461 320242 275527 320245
rect 275277 320240 275527 320242
rect 275277 320184 275282 320240
rect 275338 320184 275466 320240
rect 275522 320184 275527 320240
rect 275277 320182 275527 320184
rect 275277 320179 275343 320182
rect 275461 320179 275527 320182
rect 281717 320242 281783 320245
rect 282499 320242 282565 320245
rect 292803 320244 292869 320245
rect 292798 320242 292804 320244
rect 281717 320240 282565 320242
rect 281717 320184 281722 320240
rect 281778 320184 282504 320240
rect 282560 320184 282565 320240
rect 281717 320182 282565 320184
rect 281717 320179 281783 320182
rect 282499 320179 282565 320182
rect 284572 320182 292544 320242
rect 292712 320182 292804 320242
rect 279601 320106 279667 320109
rect 283143 320106 283209 320109
rect 279601 320104 283209 320106
rect 279601 320048 279606 320104
rect 279662 320048 283148 320104
rect 283204 320048 283209 320104
rect 279601 320046 283209 320048
rect 279601 320043 279667 320046
rect 283143 320043 283209 320046
rect 283787 320106 283853 320109
rect 283966 320106 283972 320108
rect 283787 320104 283972 320106
rect 283787 320048 283792 320104
rect 283848 320048 283972 320104
rect 283787 320046 283972 320048
rect 283787 320043 283853 320046
rect 283966 320044 283972 320046
rect 284036 320044 284042 320108
rect 215017 319970 215083 319973
rect 284572 319970 284632 320182
rect 284707 320104 284773 320109
rect 284707 320048 284712 320104
rect 284768 320048 284773 320104
rect 284707 320043 284773 320048
rect 284886 320044 284892 320108
rect 284956 320106 284962 320108
rect 285167 320106 285233 320109
rect 285438 320106 285444 320108
rect 284956 320104 285444 320106
rect 284956 320048 285172 320104
rect 285228 320048 285444 320104
rect 284956 320046 285444 320048
rect 284956 320044 284962 320046
rect 285167 320043 285233 320046
rect 285438 320044 285444 320046
rect 285508 320044 285514 320108
rect 285622 320044 285628 320108
rect 285692 320106 285698 320108
rect 286271 320106 286337 320109
rect 287099 320108 287165 320109
rect 287094 320106 287100 320108
rect 285692 320104 286337 320106
rect 285692 320048 286276 320104
rect 286332 320048 286337 320104
rect 285692 320046 286337 320048
rect 286972 320046 287100 320106
rect 285692 320044 285698 320046
rect 286271 320043 286337 320046
rect 287094 320044 287100 320046
rect 287164 320044 287170 320108
rect 288295 320106 288361 320109
rect 288022 320104 288361 320106
rect 288022 320048 288300 320104
rect 288356 320048 288361 320104
rect 288022 320046 288361 320048
rect 287099 320043 287165 320044
rect 215017 319968 284632 319970
rect 215017 319912 215022 319968
rect 215078 319912 284632 319968
rect 215017 319910 284632 319912
rect 215017 319907 215083 319910
rect 272517 319834 272583 319837
rect 280705 319834 280771 319837
rect 281993 319834 282059 319837
rect 272517 319832 282059 319834
rect 272517 319776 272522 319832
rect 272578 319776 280710 319832
rect 280766 319776 281998 319832
rect 282054 319776 282059 319832
rect 272517 319774 282059 319776
rect 272517 319771 272583 319774
rect 280705 319771 280771 319774
rect 281993 319771 282059 319774
rect 284293 319834 284359 319837
rect 284710 319834 284770 320043
rect 284293 319832 284770 319834
rect 284293 319776 284298 319832
rect 284354 319776 284770 319832
rect 284293 319774 284770 319776
rect 284293 319771 284359 319774
rect 213085 319698 213151 319701
rect 273989 319698 274055 319701
rect 274541 319698 274607 319701
rect 213085 319696 274607 319698
rect 213085 319640 213090 319696
rect 213146 319640 273994 319696
rect 274050 319640 274546 319696
rect 274602 319640 274607 319696
rect 213085 319638 274607 319640
rect 213085 319635 213151 319638
rect 273989 319635 274055 319638
rect 274541 319635 274607 319638
rect 285581 319698 285647 319701
rect 286358 319698 286364 319700
rect 285581 319696 286364 319698
rect 285581 319640 285586 319696
rect 285642 319640 286364 319696
rect 285581 319638 286364 319640
rect 285581 319635 285647 319638
rect 286358 319636 286364 319638
rect 286428 319636 286434 319700
rect 287102 319698 287162 320043
rect 288022 319834 288082 320046
rect 288295 320043 288361 320046
rect 288571 320104 288637 320109
rect 288571 320048 288576 320104
rect 288632 320048 288637 320104
rect 288571 320043 288637 320048
rect 288750 320044 288756 320108
rect 288820 320106 288826 320108
rect 288939 320106 289005 320109
rect 288820 320104 289005 320106
rect 288820 320048 288944 320104
rect 289000 320048 289005 320104
rect 288820 320046 289005 320048
rect 288820 320044 288826 320046
rect 288939 320043 289005 320046
rect 289118 320044 289124 320108
rect 289188 320106 289194 320108
rect 289307 320106 289373 320109
rect 289188 320104 289373 320106
rect 289188 320048 289312 320104
rect 289368 320048 289373 320104
rect 289188 320046 289373 320048
rect 289188 320044 289194 320046
rect 289307 320043 289373 320046
rect 289675 320104 289741 320109
rect 289675 320048 289680 320104
rect 289736 320048 289741 320104
rect 289675 320043 289741 320048
rect 289859 320104 289925 320109
rect 289859 320048 289864 320104
rect 289920 320048 289925 320104
rect 289859 320043 289925 320048
rect 290411 320104 290477 320109
rect 290411 320048 290416 320104
rect 290472 320048 290477 320104
rect 290411 320043 290477 320048
rect 290590 320044 290596 320108
rect 290660 320106 290666 320108
rect 290871 320106 290937 320109
rect 290660 320104 290937 320106
rect 290660 320048 290876 320104
rect 290932 320048 290937 320104
rect 290660 320046 290937 320048
rect 290660 320044 290666 320046
rect 290871 320043 290937 320046
rect 291423 320106 291489 320109
rect 291878 320106 291884 320108
rect 291423 320104 291884 320106
rect 291423 320048 291428 320104
rect 291484 320048 291884 320104
rect 291423 320046 291884 320048
rect 291423 320043 291489 320046
rect 291878 320044 291884 320046
rect 291948 320044 291954 320108
rect 292159 320106 292225 320109
rect 292159 320104 292406 320106
rect 292159 320048 292164 320104
rect 292220 320048 292406 320104
rect 292159 320046 292406 320048
rect 292159 320043 292225 320046
rect 288249 319834 288315 319837
rect 288022 319832 288315 319834
rect 288022 319776 288254 319832
rect 288310 319776 288315 319832
rect 288022 319774 288315 319776
rect 288249 319771 288315 319774
rect 287329 319698 287395 319701
rect 287102 319696 287395 319698
rect 287102 319640 287334 319696
rect 287390 319640 287395 319696
rect 287102 319638 287395 319640
rect 287329 319635 287395 319638
rect 287789 319698 287855 319701
rect 287973 319698 288039 319701
rect 287789 319696 288039 319698
rect 287789 319640 287794 319696
rect 287850 319640 287978 319696
rect 288034 319640 288039 319696
rect 287789 319638 288039 319640
rect 288574 319698 288634 320043
rect 289678 319837 289738 320043
rect 289678 319832 289787 319837
rect 289678 319776 289726 319832
rect 289782 319776 289787 319832
rect 289678 319774 289787 319776
rect 289721 319771 289787 319774
rect 289445 319698 289511 319701
rect 288574 319696 289511 319698
rect 288574 319640 289450 319696
rect 289506 319640 289511 319696
rect 288574 319638 289511 319640
rect 289862 319698 289922 320043
rect 290414 319837 290474 320043
rect 292346 319970 292406 320046
rect 292070 319910 292406 319970
rect 292484 319970 292544 320182
rect 292798 320180 292804 320182
rect 292868 320180 292874 320244
rect 292982 320180 292988 320244
rect 293052 320242 293058 320244
rect 293171 320242 293237 320245
rect 294183 320242 294249 320245
rect 293052 320240 293237 320242
rect 293052 320184 293176 320240
rect 293232 320184 293237 320240
rect 293052 320182 293237 320184
rect 293052 320180 293058 320182
rect 292803 320179 292869 320180
rect 293171 320179 293237 320182
rect 294140 320240 294249 320242
rect 294140 320184 294188 320240
rect 294244 320184 294249 320240
rect 294140 320179 294249 320184
rect 294551 320242 294617 320245
rect 294822 320242 294828 320244
rect 294551 320240 294828 320242
rect 294551 320184 294556 320240
rect 294612 320184 294828 320240
rect 294551 320182 294828 320184
rect 294551 320179 294617 320182
rect 294822 320180 294828 320182
rect 294892 320180 294898 320244
rect 295742 320180 295748 320244
rect 295812 320242 295818 320244
rect 295931 320242 295997 320245
rect 297035 320244 297101 320245
rect 296478 320242 296484 320244
rect 295812 320240 296484 320242
rect 295812 320184 295936 320240
rect 295992 320184 296484 320240
rect 295812 320182 296484 320184
rect 295812 320180 295818 320182
rect 295931 320179 295997 320182
rect 296478 320180 296484 320182
rect 296548 320180 296554 320244
rect 297030 320242 297036 320244
rect 296944 320182 297036 320242
rect 297030 320180 297036 320182
rect 297100 320180 297106 320244
rect 297403 320242 297469 320245
rect 298415 320242 298481 320245
rect 302003 320244 302069 320245
rect 299422 320242 299428 320244
rect 297403 320240 297834 320242
rect 297403 320184 297408 320240
rect 297464 320184 297834 320240
rect 297403 320182 297834 320184
rect 297035 320179 297101 320180
rect 297403 320179 297469 320182
rect 293166 320044 293172 320108
rect 293236 320106 293242 320108
rect 293447 320106 293513 320109
rect 293236 320104 293513 320106
rect 293236 320048 293452 320104
rect 293508 320048 293513 320104
rect 293236 320046 293513 320048
rect 293236 320044 293242 320046
rect 293447 320043 293513 320046
rect 292484 319939 293280 319970
rect 292484 319934 293329 319939
rect 292484 319910 293268 319934
rect 290414 319832 290523 319837
rect 290414 319776 290462 319832
rect 290518 319776 290523 319832
rect 290414 319774 290523 319776
rect 290457 319771 290523 319774
rect 292070 319701 292130 319910
rect 293220 319878 293268 319910
rect 293324 319878 293329 319934
rect 293220 319873 293329 319878
rect 290273 319698 290339 319701
rect 289862 319696 290339 319698
rect 289862 319640 290278 319696
rect 290334 319640 290339 319696
rect 289862 319638 290339 319640
rect 287789 319635 287855 319638
rect 287973 319635 288039 319638
rect 289445 319635 289511 319638
rect 290273 319635 290339 319638
rect 291101 319700 291167 319701
rect 291101 319696 291148 319700
rect 291212 319698 291218 319700
rect 291101 319640 291106 319696
rect 291101 319636 291148 319640
rect 291212 319638 291258 319698
rect 292070 319696 292179 319701
rect 292070 319640 292118 319696
rect 292174 319640 292179 319696
rect 292070 319638 292179 319640
rect 291212 319636 291218 319638
rect 291101 319635 291167 319636
rect 292113 319635 292179 319638
rect 292481 319698 292547 319701
rect 293033 319698 293099 319701
rect 292481 319696 293099 319698
rect 292481 319640 292486 319696
rect 292542 319640 293038 319696
rect 293094 319640 293099 319696
rect 292481 319638 293099 319640
rect 293220 319698 293280 319873
rect 294140 319837 294200 320179
rect 294275 320104 294341 320109
rect 294459 320108 294525 320109
rect 294275 320048 294280 320104
rect 294336 320048 294341 320104
rect 294275 320043 294341 320048
rect 294454 320044 294460 320108
rect 294524 320106 294530 320108
rect 294735 320106 294801 320109
rect 295190 320106 295196 320108
rect 294524 320046 294616 320106
rect 294735 320104 295196 320106
rect 294735 320048 294740 320104
rect 294796 320048 295196 320104
rect 294735 320046 295196 320048
rect 294524 320044 294530 320046
rect 294459 320043 294525 320044
rect 294735 320043 294801 320046
rect 295190 320044 295196 320046
rect 295260 320044 295266 320108
rect 296115 320106 296181 320109
rect 295750 320104 296181 320106
rect 295750 320048 296120 320104
rect 296176 320048 296181 320104
rect 295750 320046 296181 320048
rect 294278 319970 294338 320043
rect 295006 319970 295012 319972
rect 294278 319910 295012 319970
rect 295006 319908 295012 319910
rect 295076 319908 295082 319972
rect 295290 319939 295534 319970
rect 295290 319934 295537 319939
rect 295290 319910 295476 319934
rect 294137 319832 294203 319837
rect 294137 319776 294142 319832
rect 294198 319776 294203 319832
rect 294137 319771 294203 319776
rect 294413 319834 294479 319837
rect 295290 319834 295350 319910
rect 295471 319878 295476 319910
rect 295532 319878 295537 319934
rect 295471 319873 295537 319878
rect 294413 319832 295350 319834
rect 294413 319776 294418 319832
rect 294474 319776 295350 319832
rect 294413 319774 295350 319776
rect 294413 319771 294479 319774
rect 295609 319698 295675 319701
rect 295750 319698 295810 320046
rect 296115 320043 296181 320046
rect 296299 320104 296365 320109
rect 296299 320048 296304 320104
rect 296360 320048 296365 320104
rect 296299 320043 296365 320048
rect 297219 320104 297285 320109
rect 297587 320108 297653 320109
rect 297582 320106 297588 320108
rect 297219 320048 297224 320104
rect 297280 320048 297285 320104
rect 297219 320043 297285 320048
rect 297460 320046 297588 320106
rect 297582 320044 297588 320046
rect 297652 320044 297658 320108
rect 297587 320043 297653 320044
rect 296161 319836 296227 319837
rect 296110 319834 296116 319836
rect 296070 319774 296116 319834
rect 296180 319832 296227 319836
rect 296222 319776 296227 319832
rect 296110 319772 296116 319774
rect 296180 319772 296227 319776
rect 296161 319771 296227 319772
rect 293220 319638 293786 319698
rect 292481 319635 292547 319638
rect 293033 319635 293099 319638
rect 207933 319562 207999 319565
rect 281809 319562 281875 319565
rect 282545 319562 282611 319565
rect 292665 319562 292731 319565
rect 207933 319560 282611 319562
rect 207933 319504 207938 319560
rect 207994 319504 281814 319560
rect 281870 319504 282550 319560
rect 282606 319504 282611 319560
rect 207933 319502 282611 319504
rect 207933 319499 207999 319502
rect 281809 319499 281875 319502
rect 282545 319499 282611 319502
rect 282686 319560 292731 319562
rect 282686 319504 292670 319560
rect 292726 319504 292731 319560
rect 282686 319502 292731 319504
rect 208025 319426 208091 319429
rect 281717 319426 281783 319429
rect 208025 319424 281783 319426
rect -960 319290 480 319380
rect 208025 319368 208030 319424
rect 208086 319368 281722 319424
rect 281778 319368 281783 319424
rect 208025 319366 281783 319368
rect 208025 319363 208091 319366
rect 281717 319363 281783 319366
rect 281901 319426 281967 319429
rect 282686 319426 282746 319502
rect 292665 319499 292731 319502
rect 292798 319500 292804 319564
rect 292868 319562 292874 319564
rect 293585 319562 293651 319565
rect 292868 319560 293651 319562
rect 292868 319504 293590 319560
rect 293646 319504 293651 319560
rect 292868 319502 293651 319504
rect 293726 319562 293786 319638
rect 295609 319696 295810 319698
rect 295609 319640 295614 319696
rect 295670 319640 295810 319696
rect 295609 319638 295810 319640
rect 296161 319698 296227 319701
rect 296302 319698 296362 320043
rect 296161 319696 296362 319698
rect 296161 319640 296166 319696
rect 296222 319640 296362 319696
rect 296161 319638 296362 319640
rect 297222 319701 297282 320043
rect 297590 319836 297650 320043
rect 297582 319772 297588 319836
rect 297652 319772 297658 319836
rect 297774 319834 297834 320182
rect 298415 320240 299428 320242
rect 298415 320184 298420 320240
rect 298476 320184 299428 320240
rect 298415 320182 299428 320184
rect 298415 320179 298481 320182
rect 299422 320180 299428 320182
rect 299492 320180 299498 320244
rect 300894 320180 300900 320244
rect 300964 320242 300970 320244
rect 301998 320242 302004 320244
rect 300964 320182 302004 320242
rect 300964 320180 300970 320182
rect 301998 320180 302004 320182
rect 302068 320180 302074 320244
rect 302182 320180 302188 320244
rect 302252 320242 302258 320244
rect 307702 320242 307708 320244
rect 302252 320182 307708 320242
rect 302252 320180 302258 320182
rect 307702 320180 307708 320182
rect 307772 320180 307778 320244
rect 307983 320242 308049 320245
rect 311850 320242 311910 320454
rect 322054 320452 322060 320454
rect 322124 320452 322130 320516
rect 322243 320514 322309 320517
rect 323347 320516 323413 320517
rect 322606 320514 322612 320516
rect 322243 320512 322612 320514
rect 322243 320456 322248 320512
rect 322304 320456 322612 320512
rect 322243 320454 322612 320456
rect 322059 320451 322125 320452
rect 322243 320451 322309 320454
rect 322606 320452 322612 320454
rect 322676 320452 322682 320516
rect 323342 320514 323348 320516
rect 323256 320454 323348 320514
rect 323342 320452 323348 320454
rect 323412 320452 323418 320516
rect 323526 320452 323532 320516
rect 323596 320514 323602 320516
rect 323807 320514 323873 320517
rect 323596 320512 323873 320514
rect 323596 320456 323812 320512
rect 323868 320456 323873 320512
rect 323596 320454 323873 320456
rect 323596 320452 323602 320454
rect 323347 320451 323413 320452
rect 323807 320451 323873 320454
rect 324635 320514 324701 320517
rect 324998 320514 325004 320516
rect 324635 320512 325004 320514
rect 324635 320456 324640 320512
rect 324696 320456 325004 320512
rect 324635 320454 325004 320456
rect 324635 320451 324701 320454
rect 324998 320452 325004 320454
rect 325068 320452 325074 320516
rect 326107 320514 326173 320517
rect 327625 320514 327691 320517
rect 326107 320512 327691 320514
rect 326107 320456 326112 320512
rect 326168 320456 327630 320512
rect 327686 320456 327691 320512
rect 326107 320454 327691 320456
rect 326107 320451 326173 320454
rect 327625 320451 327691 320454
rect 327809 320514 327875 320517
rect 327809 320512 335370 320514
rect 327809 320456 327814 320512
rect 327870 320456 335370 320512
rect 327809 320454 335370 320456
rect 327809 320451 327875 320454
rect 316447 320378 316513 320381
rect 316447 320376 318994 320378
rect 316447 320320 316452 320376
rect 316508 320320 318994 320376
rect 316447 320318 318994 320320
rect 316447 320315 316513 320318
rect 307983 320240 311910 320242
rect 307983 320184 307988 320240
rect 308044 320184 311910 320240
rect 307983 320182 311910 320184
rect 312031 320242 312097 320245
rect 312675 320242 312741 320245
rect 313595 320242 313661 320245
rect 313958 320242 313964 320244
rect 312031 320240 312370 320242
rect 312031 320184 312036 320240
rect 312092 320184 312370 320240
rect 312031 320182 312370 320184
rect 302003 320179 302069 320180
rect 307983 320179 308049 320182
rect 312031 320179 312097 320182
rect 298047 320106 298113 320109
rect 299243 320108 299309 320109
rect 299238 320106 299244 320108
rect 298004 320104 298113 320106
rect 298004 320048 298052 320104
rect 298108 320048 298113 320104
rect 298004 320043 298113 320048
rect 299152 320046 299244 320106
rect 299238 320044 299244 320046
rect 299308 320044 299314 320108
rect 299611 320106 299677 320109
rect 299790 320106 299796 320108
rect 299611 320104 299796 320106
rect 299611 320048 299616 320104
rect 299672 320048 299796 320104
rect 299611 320046 299796 320048
rect 299243 320043 299309 320044
rect 299611 320043 299677 320046
rect 299790 320044 299796 320046
rect 299860 320044 299866 320108
rect 300715 320104 300781 320109
rect 300715 320048 300720 320104
rect 300776 320048 300781 320104
rect 300715 320043 300781 320048
rect 300899 320104 300965 320109
rect 300899 320048 300904 320104
rect 300960 320048 300965 320104
rect 300899 320043 300965 320048
rect 301262 320044 301268 320108
rect 301332 320106 301338 320108
rect 301727 320106 301793 320109
rect 301332 320104 301793 320106
rect 301332 320048 301732 320104
rect 301788 320048 301793 320104
rect 301332 320046 301793 320048
rect 301332 320044 301338 320046
rect 301727 320043 301793 320046
rect 302187 320104 302253 320109
rect 302187 320048 302192 320104
rect 302248 320048 302253 320104
rect 302187 320043 302253 320048
rect 302366 320044 302372 320108
rect 302436 320106 302442 320108
rect 302831 320106 302897 320109
rect 303935 320106 304001 320109
rect 302436 320104 302897 320106
rect 302436 320048 302836 320104
rect 302892 320048 302897 320104
rect 302436 320046 302897 320048
rect 302436 320044 302442 320046
rect 302831 320043 302897 320046
rect 303662 320104 304001 320106
rect 303662 320048 303940 320104
rect 303996 320048 304001 320104
rect 303662 320046 304001 320048
rect 298004 319972 298064 320043
rect 297950 319908 297956 319972
rect 298020 319910 298064 319972
rect 298878 319939 299352 319970
rect 298875 319934 299352 319939
rect 298020 319908 298026 319910
rect 298875 319878 298880 319934
rect 298936 319910 299352 319934
rect 298936 319878 298941 319910
rect 298875 319873 298941 319878
rect 298001 319834 298067 319837
rect 297774 319832 298067 319834
rect 297774 319776 298006 319832
rect 298062 319776 298067 319832
rect 297774 319774 298067 319776
rect 298001 319771 298067 319774
rect 299292 319701 299352 319910
rect 297222 319696 297331 319701
rect 297222 319640 297270 319696
rect 297326 319640 297331 319696
rect 297222 319638 297331 319640
rect 295609 319635 295675 319638
rect 296161 319635 296227 319638
rect 297265 319635 297331 319638
rect 298185 319698 298251 319701
rect 298502 319698 298508 319700
rect 298185 319696 298508 319698
rect 298185 319640 298190 319696
rect 298246 319640 298508 319696
rect 298185 319638 298508 319640
rect 298185 319635 298251 319638
rect 298502 319636 298508 319638
rect 298572 319636 298578 319700
rect 298737 319698 298803 319701
rect 299054 319698 299060 319700
rect 298737 319696 299060 319698
rect 298737 319640 298742 319696
rect 298798 319640 299060 319696
rect 298737 319638 299060 319640
rect 298737 319635 298803 319638
rect 299054 319636 299060 319638
rect 299124 319636 299130 319700
rect 299289 319696 299355 319701
rect 299289 319640 299294 319696
rect 299350 319640 299355 319696
rect 299289 319635 299355 319640
rect 299565 319698 299631 319701
rect 300718 319698 300778 320043
rect 299565 319696 300778 319698
rect 299565 319640 299570 319696
rect 299626 319640 300778 319696
rect 299565 319638 300778 319640
rect 300902 319698 300962 320043
rect 301630 319970 301636 319972
rect 301270 319939 301636 319970
rect 301267 319934 301636 319939
rect 301267 319878 301272 319934
rect 301328 319910 301636 319934
rect 301328 319878 301333 319910
rect 301630 319908 301636 319910
rect 301700 319908 301706 319972
rect 301267 319873 301333 319878
rect 301313 319698 301379 319701
rect 300902 319696 301379 319698
rect 300902 319640 301318 319696
rect 301374 319640 301379 319696
rect 300902 319638 301379 319640
rect 299565 319635 299631 319638
rect 301313 319635 301379 319638
rect 301865 319698 301931 319701
rect 302190 319698 302250 320043
rect 302555 319934 302621 319939
rect 302555 319878 302560 319934
rect 302616 319878 302621 319934
rect 302555 319873 302621 319878
rect 301865 319696 302250 319698
rect 301865 319640 301870 319696
rect 301926 319640 302250 319696
rect 301865 319638 302250 319640
rect 302558 319698 302618 319873
rect 302693 319698 302759 319701
rect 303337 319700 303403 319701
rect 302558 319696 302759 319698
rect 302558 319640 302698 319696
rect 302754 319640 302759 319696
rect 302558 319638 302759 319640
rect 301865 319635 301931 319638
rect 302693 319635 302759 319638
rect 303286 319636 303292 319700
rect 303356 319698 303403 319700
rect 303662 319698 303722 320046
rect 303935 320043 304001 320046
rect 304211 320104 304277 320109
rect 304211 320048 304216 320104
rect 304272 320048 304277 320104
rect 304211 320043 304277 320048
rect 304579 320104 304645 320109
rect 304579 320048 304584 320104
rect 304640 320048 304645 320104
rect 304579 320043 304645 320048
rect 305494 320044 305500 320108
rect 305564 320106 305570 320108
rect 305867 320106 305933 320109
rect 306327 320106 306393 320109
rect 305564 320104 305933 320106
rect 305564 320048 305872 320104
rect 305928 320048 305933 320104
rect 305564 320046 305933 320048
rect 305564 320044 305570 320046
rect 305867 320043 305933 320046
rect 306054 320104 306393 320106
rect 306054 320048 306332 320104
rect 306388 320048 306393 320104
rect 306054 320046 306393 320048
rect 304214 319701 304274 320043
rect 304582 319701 304642 320043
rect 305131 319934 305197 319939
rect 305131 319878 305136 319934
rect 305192 319878 305197 319934
rect 305678 319908 305684 319972
rect 305748 319970 305754 319972
rect 306054 319970 306114 320046
rect 306327 320043 306393 320046
rect 306971 320104 307037 320109
rect 307523 320108 307589 320109
rect 307518 320106 307524 320108
rect 306971 320048 306976 320104
rect 307032 320048 307037 320104
rect 306971 320043 307037 320048
rect 307432 320046 307524 320106
rect 307518 320044 307524 320046
rect 307588 320044 307594 320108
rect 307702 320044 307708 320108
rect 307772 320106 307778 320108
rect 308627 320106 308693 320109
rect 308990 320106 308996 320108
rect 307772 320104 308996 320106
rect 307772 320048 308632 320104
rect 308688 320048 308996 320104
rect 307772 320046 308996 320048
rect 307772 320044 307778 320046
rect 307523 320043 307589 320044
rect 308627 320043 308693 320046
rect 308990 320044 308996 320046
rect 309060 320044 309066 320108
rect 309731 320106 309797 320109
rect 309596 320104 309797 320106
rect 309596 320048 309736 320104
rect 309792 320048 309797 320104
rect 309596 320046 309797 320048
rect 305748 319910 306114 319970
rect 305748 319908 305754 319910
rect 305131 319873 305197 319878
rect 303356 319696 303448 319698
rect 303398 319640 303448 319696
rect 303356 319638 303448 319640
rect 303662 319638 304090 319698
rect 304214 319696 304323 319701
rect 304214 319640 304262 319696
rect 304318 319640 304323 319696
rect 304214 319638 304323 319640
rect 303356 319636 303403 319638
rect 303337 319635 303403 319636
rect 304030 319565 304090 319638
rect 304257 319635 304323 319638
rect 304533 319696 304642 319701
rect 304533 319640 304538 319696
rect 304594 319640 304642 319696
rect 304533 319638 304642 319640
rect 304533 319635 304599 319638
rect 293726 319502 302618 319562
rect 304030 319560 304139 319565
rect 304030 319504 304078 319560
rect 304134 319504 304139 319560
rect 304030 319502 304139 319504
rect 292868 319500 292874 319502
rect 293585 319499 293651 319502
rect 281901 319424 282746 319426
rect 281901 319368 281906 319424
rect 281962 319368 282746 319424
rect 281901 319366 282746 319368
rect 283281 319426 283347 319429
rect 283598 319426 283604 319428
rect 283281 319424 283604 319426
rect 283281 319368 283286 319424
rect 283342 319368 283604 319424
rect 283281 319366 283604 319368
rect 281901 319363 281967 319366
rect 283281 319363 283347 319366
rect 283598 319364 283604 319366
rect 283668 319364 283674 319428
rect 283741 319426 283807 319429
rect 302366 319426 302372 319428
rect 283741 319424 302372 319426
rect 283741 319368 283746 319424
rect 283802 319368 302372 319424
rect 283741 319366 302372 319368
rect 283741 319363 283807 319366
rect 302366 319364 302372 319366
rect 302436 319364 302442 319428
rect 302558 319426 302618 319502
rect 304073 319499 304139 319502
rect 304993 319562 305059 319565
rect 305134 319562 305194 319873
rect 306741 319834 306807 319837
rect 306974 319834 307034 320043
rect 309596 319837 309656 320046
rect 309731 320043 309797 320046
rect 309915 320104 309981 320109
rect 310927 320106 310993 320109
rect 309915 320048 309920 320104
rect 309976 320048 309981 320104
rect 309915 320043 309981 320048
rect 310470 320104 310993 320106
rect 310470 320048 310932 320104
rect 310988 320048 310993 320104
rect 310470 320046 310993 320048
rect 309918 319837 309978 320043
rect 306741 319832 307034 319834
rect 306741 319776 306746 319832
rect 306802 319776 307034 319832
rect 306741 319774 307034 319776
rect 309593 319832 309659 319837
rect 309593 319776 309598 319832
rect 309654 319776 309659 319832
rect 306741 319771 306807 319774
rect 309593 319771 309659 319776
rect 309869 319832 309978 319837
rect 309869 319776 309874 319832
rect 309930 319776 309978 319832
rect 309869 319774 309978 319776
rect 310145 319834 310211 319837
rect 310470 319834 310530 320046
rect 310927 320043 310993 320046
rect 311198 320044 311204 320108
rect 311268 320106 311274 320108
rect 311663 320106 311729 320109
rect 311939 320108 312005 320109
rect 311268 320104 311729 320106
rect 311268 320048 311668 320104
rect 311724 320048 311729 320104
rect 311268 320046 311729 320048
rect 311268 320044 311274 320046
rect 311663 320043 311729 320046
rect 311934 320044 311940 320108
rect 312004 320106 312010 320108
rect 312004 320046 312096 320106
rect 312004 320044 312010 320046
rect 311939 320043 312005 320044
rect 310145 319832 310530 319834
rect 310145 319776 310150 319832
rect 310206 319776 310530 319832
rect 310145 319774 310530 319776
rect 312310 319834 312370 320182
rect 312675 320240 313290 320242
rect 312675 320184 312680 320240
rect 312736 320184 313290 320240
rect 312675 320182 313290 320184
rect 312675 320179 312741 320182
rect 312486 320044 312492 320108
rect 312556 320106 312562 320108
rect 312767 320106 312833 320109
rect 313038 320106 313044 320108
rect 312556 320104 313044 320106
rect 312556 320048 312772 320104
rect 312828 320048 313044 320104
rect 312556 320046 313044 320048
rect 312556 320044 312562 320046
rect 312767 320043 312833 320046
rect 313038 320044 313044 320046
rect 313108 320044 313114 320108
rect 312813 319834 312879 319837
rect 312310 319832 312879 319834
rect 312310 319776 312818 319832
rect 312874 319776 312879 319832
rect 312310 319774 312879 319776
rect 309869 319771 309935 319774
rect 310145 319771 310211 319774
rect 312813 319771 312879 319774
rect 313089 319834 313155 319837
rect 313230 319834 313290 320182
rect 313595 320240 313964 320242
rect 313595 320184 313600 320240
rect 313656 320184 313964 320240
rect 313595 320182 313964 320184
rect 313595 320179 313661 320182
rect 313958 320180 313964 320182
rect 314028 320180 314034 320244
rect 314147 320242 314213 320245
rect 314326 320242 314332 320244
rect 314147 320240 314332 320242
rect 314147 320184 314152 320240
rect 314208 320184 314332 320240
rect 314147 320182 314332 320184
rect 314147 320179 314213 320182
rect 314326 320180 314332 320182
rect 314396 320180 314402 320244
rect 316631 320242 316697 320245
rect 316036 320240 316697 320242
rect 316036 320184 316636 320240
rect 316692 320184 316697 320240
rect 316036 320182 316697 320184
rect 313411 320104 313477 320109
rect 313411 320048 313416 320104
rect 313472 320048 313477 320104
rect 313411 320043 313477 320048
rect 313590 320044 313596 320108
rect 313660 320106 313666 320108
rect 314142 320106 314148 320108
rect 313660 320046 314148 320106
rect 313660 320044 313666 320046
rect 314142 320044 314148 320046
rect 314212 320106 314218 320108
rect 314423 320106 314489 320109
rect 314883 320106 314949 320109
rect 314212 320104 314489 320106
rect 314212 320048 314428 320104
rect 314484 320048 314489 320104
rect 314212 320046 314489 320048
rect 314212 320044 314218 320046
rect 314423 320043 314489 320046
rect 314702 320104 314949 320106
rect 314702 320048 314888 320104
rect 314944 320048 314949 320104
rect 314702 320046 314949 320048
rect 313089 319832 313290 319834
rect 313089 319776 313094 319832
rect 313150 319776 313290 319832
rect 313089 319774 313290 319776
rect 313089 319771 313155 319774
rect 309542 319636 309548 319700
rect 309612 319698 309618 319700
rect 311893 319698 311959 319701
rect 309612 319696 311959 319698
rect 309612 319640 311898 319696
rect 311954 319640 311959 319696
rect 309612 319638 311959 319640
rect 309612 319636 309618 319638
rect 311893 319635 311959 319638
rect 313273 319698 313339 319701
rect 313414 319698 313474 320043
rect 314702 319837 314762 320046
rect 314883 320043 314949 320046
rect 315062 320044 315068 320108
rect 315132 320106 315138 320108
rect 315251 320106 315317 320109
rect 315614 320106 315620 320108
rect 315132 320104 315620 320106
rect 315132 320048 315256 320104
rect 315312 320048 315620 320104
rect 315132 320046 315620 320048
rect 315132 320044 315138 320046
rect 315251 320043 315317 320046
rect 315614 320044 315620 320046
rect 315684 320044 315690 320108
rect 313687 319834 313753 319837
rect 313273 319696 313474 319698
rect 313273 319640 313278 319696
rect 313334 319640 313474 319696
rect 313273 319638 313474 319640
rect 313644 319832 313753 319834
rect 313644 319776 313692 319832
rect 313748 319776 313753 319832
rect 313644 319771 313753 319776
rect 314653 319832 314762 319837
rect 314653 319776 314658 319832
rect 314714 319776 314762 319832
rect 314653 319774 314762 319776
rect 314653 319771 314719 319774
rect 313273 319635 313339 319638
rect 313644 319565 313704 319771
rect 316036 319701 316096 320182
rect 316631 320179 316697 320182
rect 317735 320242 317801 320245
rect 318558 320242 318564 320244
rect 317735 320240 318564 320242
rect 317735 320184 317740 320240
rect 317796 320184 318564 320240
rect 317735 320182 318564 320184
rect 317735 320179 317801 320182
rect 318558 320180 318564 320182
rect 318628 320180 318634 320244
rect 318934 320242 318994 320318
rect 319294 320316 319300 320380
rect 319364 320378 319370 320380
rect 320127 320378 320193 320381
rect 319364 320376 320193 320378
rect 319364 320320 320132 320376
rect 320188 320320 320193 320376
rect 319364 320318 320193 320320
rect 319364 320316 319370 320318
rect 320127 320315 320193 320318
rect 320311 320378 320377 320381
rect 320582 320378 320588 320380
rect 320311 320376 320588 320378
rect 320311 320320 320316 320376
rect 320372 320320 320588 320376
rect 320311 320318 320588 320320
rect 320311 320315 320377 320318
rect 320582 320316 320588 320318
rect 320652 320316 320658 320380
rect 320771 320378 320837 320381
rect 321318 320378 321324 320380
rect 320771 320376 321324 320378
rect 320771 320320 320776 320376
rect 320832 320320 321324 320376
rect 320771 320318 321324 320320
rect 320771 320315 320837 320318
rect 321318 320316 321324 320318
rect 321388 320316 321394 320380
rect 321599 320378 321665 320381
rect 322422 320378 322428 320380
rect 321599 320376 322428 320378
rect 321599 320320 321604 320376
rect 321660 320320 322428 320376
rect 321599 320318 322428 320320
rect 321599 320315 321665 320318
rect 322422 320316 322428 320318
rect 322492 320316 322498 320380
rect 323255 320378 323321 320381
rect 324267 320380 324333 320381
rect 323894 320378 323900 320380
rect 323255 320376 323900 320378
rect 323255 320320 323260 320376
rect 323316 320320 323900 320376
rect 323255 320318 323900 320320
rect 323255 320315 323321 320318
rect 323894 320316 323900 320318
rect 323964 320316 323970 320380
rect 324262 320378 324268 320380
rect 324176 320318 324268 320378
rect 324262 320316 324268 320318
rect 324332 320316 324338 320380
rect 324446 320316 324452 320380
rect 324516 320378 324522 320380
rect 325463 320378 325529 320381
rect 324516 320376 325529 320378
rect 324516 320320 325468 320376
rect 325524 320320 325529 320376
rect 324516 320318 325529 320320
rect 324516 320316 324522 320318
rect 324267 320315 324333 320316
rect 325463 320315 325529 320318
rect 326383 320378 326449 320381
rect 327395 320380 327461 320381
rect 326654 320378 326660 320380
rect 326383 320376 326660 320378
rect 326383 320320 326388 320376
rect 326444 320320 326660 320376
rect 326383 320318 326660 320320
rect 326383 320315 326449 320318
rect 326654 320316 326660 320318
rect 326724 320316 326730 320380
rect 327390 320378 327396 320380
rect 327304 320318 327396 320378
rect 327390 320316 327396 320318
rect 327460 320316 327466 320380
rect 327625 320378 327691 320381
rect 327758 320378 327764 320380
rect 327625 320376 327764 320378
rect 327625 320320 327630 320376
rect 327686 320320 327764 320376
rect 327625 320318 327764 320320
rect 327395 320315 327461 320316
rect 327625 320315 327691 320318
rect 327758 320316 327764 320318
rect 327828 320316 327834 320380
rect 327901 320378 327967 320381
rect 334525 320378 334591 320381
rect 327901 320376 334591 320378
rect 327901 320320 327906 320376
rect 327962 320320 334530 320376
rect 334586 320320 334591 320376
rect 327901 320318 334591 320320
rect 335310 320378 335370 320454
rect 336825 320378 336891 320381
rect 337929 320378 337995 320381
rect 335310 320376 337995 320378
rect 335310 320320 336830 320376
rect 336886 320320 337934 320376
rect 337990 320320 337995 320376
rect 335310 320318 337995 320320
rect 327901 320315 327967 320318
rect 334525 320315 334591 320318
rect 336825 320315 336891 320318
rect 337929 320315 337995 320318
rect 336917 320242 336983 320245
rect 318934 320240 336983 320242
rect 318934 320184 336922 320240
rect 336978 320184 336983 320240
rect 318934 320182 336983 320184
rect 336917 320179 336983 320182
rect 338113 320242 338179 320245
rect 339309 320242 339375 320245
rect 338113 320240 339375 320242
rect 338113 320184 338118 320240
rect 338174 320184 339314 320240
rect 339370 320184 339375 320240
rect 338113 320182 339375 320184
rect 338113 320179 338179 320182
rect 339309 320179 339375 320182
rect 316171 320104 316237 320109
rect 316171 320048 316176 320104
rect 316232 320048 316237 320104
rect 316171 320043 316237 320048
rect 316718 320044 316724 320108
rect 316788 320106 316794 320108
rect 316907 320106 316973 320109
rect 317270 320106 317276 320108
rect 316788 320104 317276 320106
rect 316788 320048 316912 320104
rect 316968 320048 317276 320104
rect 316788 320046 317276 320048
rect 316788 320044 316794 320046
rect 316907 320043 316973 320046
rect 317270 320044 317276 320046
rect 317340 320044 317346 320108
rect 317638 320044 317644 320108
rect 317708 320106 317714 320108
rect 318287 320106 318353 320109
rect 317708 320104 318353 320106
rect 317708 320048 318292 320104
rect 318348 320048 318353 320104
rect 317708 320046 318353 320048
rect 317708 320044 317714 320046
rect 318287 320043 318353 320046
rect 318563 320106 318629 320109
rect 319115 320108 319181 320109
rect 319110 320106 319116 320108
rect 318563 320104 318810 320106
rect 318563 320048 318568 320104
rect 318624 320048 318810 320104
rect 318563 320046 318810 320048
rect 319024 320046 319116 320106
rect 318563 320043 318629 320046
rect 313958 319636 313964 319700
rect 314028 319698 314034 319700
rect 314101 319698 314167 319701
rect 314028 319696 314167 319698
rect 314028 319640 314106 319696
rect 314162 319640 314167 319696
rect 314028 319638 314167 319640
rect 314028 319636 314034 319638
rect 314101 319635 314167 319638
rect 315430 319636 315436 319700
rect 315500 319698 315506 319700
rect 315573 319698 315639 319701
rect 315500 319696 315639 319698
rect 315500 319640 315578 319696
rect 315634 319640 315639 319696
rect 315500 319638 315639 319640
rect 315500 319636 315506 319638
rect 315573 319635 315639 319638
rect 316033 319696 316099 319701
rect 316033 319640 316038 319696
rect 316094 319640 316099 319696
rect 316033 319635 316099 319640
rect 316174 319698 316234 320043
rect 318750 319970 318810 320046
rect 319110 320044 319116 320046
rect 319180 320044 319186 320108
rect 319478 320044 319484 320108
rect 319548 320106 319554 320108
rect 319667 320106 319733 320109
rect 320030 320106 320036 320108
rect 319548 320104 320036 320106
rect 319548 320048 319672 320104
rect 319728 320048 320036 320104
rect 319548 320046 320036 320048
rect 319548 320044 319554 320046
rect 319115 320043 319181 320044
rect 319667 320043 319733 320046
rect 320030 320044 320036 320046
rect 320100 320044 320106 320108
rect 320398 320044 320404 320108
rect 320468 320106 320474 320108
rect 320679 320106 320745 320109
rect 320468 320104 320745 320106
rect 320468 320048 320684 320104
rect 320740 320048 320745 320104
rect 320468 320046 320745 320048
rect 320468 320044 320474 320046
rect 320679 320043 320745 320046
rect 321323 320106 321389 320109
rect 321502 320106 321508 320108
rect 321323 320104 321508 320106
rect 321323 320048 321328 320104
rect 321384 320048 321508 320104
rect 321323 320046 321508 320048
rect 321323 320043 321389 320046
rect 321502 320044 321508 320046
rect 321572 320044 321578 320108
rect 322519 320104 322585 320109
rect 322519 320048 322524 320104
rect 322580 320048 322585 320104
rect 322519 320043 322585 320048
rect 324630 320044 324636 320108
rect 324700 320106 324706 320108
rect 324911 320106 324977 320109
rect 326843 320108 326909 320109
rect 326838 320106 326844 320108
rect 324700 320104 324977 320106
rect 324700 320048 324916 320104
rect 324972 320048 324977 320104
rect 324700 320046 324977 320048
rect 326752 320046 326844 320106
rect 324700 320044 324706 320046
rect 324911 320043 324977 320046
rect 326838 320044 326844 320046
rect 326908 320044 326914 320108
rect 327211 320106 327277 320109
rect 328913 320106 328979 320109
rect 331673 320106 331739 320109
rect 327211 320104 328979 320106
rect 327211 320048 327216 320104
rect 327272 320048 328918 320104
rect 328974 320048 328979 320104
rect 327211 320046 328979 320048
rect 326843 320043 326909 320044
rect 327211 320043 327277 320046
rect 328913 320043 328979 320046
rect 329054 320104 331739 320106
rect 329054 320048 331678 320104
rect 331734 320048 331739 320104
rect 329054 320046 331739 320048
rect 322522 319970 322582 320043
rect 329054 319970 329114 320046
rect 331673 320043 331739 320046
rect 318750 319910 319546 319970
rect 319253 319834 319319 319837
rect 317232 319832 319319 319834
rect 317232 319776 319258 319832
rect 319314 319776 319319 319832
rect 317232 319774 319319 319776
rect 317045 319698 317111 319701
rect 316174 319696 317111 319698
rect 316174 319640 317050 319696
rect 317106 319640 317111 319696
rect 316174 319638 317111 319640
rect 317045 319635 317111 319638
rect 304993 319560 305194 319562
rect 304993 319504 304998 319560
rect 305054 319504 305194 319560
rect 304993 319502 305194 319504
rect 304993 319499 305059 319502
rect 309910 319500 309916 319564
rect 309980 319562 309986 319564
rect 310145 319562 310211 319565
rect 310697 319564 310763 319565
rect 309980 319560 310211 319562
rect 309980 319504 310150 319560
rect 310206 319504 310211 319560
rect 309980 319502 310211 319504
rect 309980 319500 309986 319502
rect 310145 319499 310211 319502
rect 310646 319500 310652 319564
rect 310716 319562 310763 319564
rect 310716 319560 310808 319562
rect 310758 319504 310808 319560
rect 310716 319502 310808 319504
rect 313641 319560 313707 319565
rect 313641 319504 313646 319560
rect 313702 319504 313707 319560
rect 310716 319500 310763 319502
rect 310697 319499 310763 319500
rect 313641 319499 313707 319504
rect 317232 319426 317292 319774
rect 319253 319771 319319 319774
rect 317873 319698 317939 319701
rect 319486 319698 319546 319910
rect 321231 319936 321297 319939
rect 321231 319934 321570 319936
rect 321231 319878 321236 319934
rect 321292 319878 321570 319934
rect 322522 319910 329114 319970
rect 329189 319970 329255 319973
rect 333973 319970 334039 319973
rect 329189 319968 334039 319970
rect 329189 319912 329194 319968
rect 329250 319912 333978 319968
rect 334034 319912 334039 319968
rect 329189 319910 334039 319912
rect 329189 319907 329255 319910
rect 333973 319907 334039 319910
rect 321231 319876 321570 319878
rect 321231 319873 321297 319876
rect 320173 319698 320239 319701
rect 317873 319696 318074 319698
rect 317873 319640 317878 319696
rect 317934 319640 318074 319696
rect 317873 319638 318074 319640
rect 319486 319696 320239 319698
rect 319486 319640 320178 319696
rect 320234 319640 320239 319696
rect 319486 319638 320239 319640
rect 317873 319635 317939 319638
rect 317454 319500 317460 319564
rect 317524 319562 317530 319564
rect 317873 319562 317939 319565
rect 317524 319560 317939 319562
rect 317524 319504 317878 319560
rect 317934 319504 317939 319560
rect 317524 319502 317939 319504
rect 318014 319562 318074 319638
rect 320173 319635 320239 319638
rect 321369 319698 321435 319701
rect 321510 319698 321570 319876
rect 322105 319834 322171 319837
rect 352414 319834 352420 319836
rect 322105 319832 352420 319834
rect 322105 319776 322110 319832
rect 322166 319776 352420 319832
rect 322105 319774 352420 319776
rect 322105 319771 322171 319774
rect 352414 319772 352420 319774
rect 352484 319772 352490 319836
rect 321369 319696 321570 319698
rect 321369 319640 321374 319696
rect 321430 319640 321570 319696
rect 321369 319638 321570 319640
rect 321737 319698 321803 319701
rect 322289 319698 322355 319701
rect 321737 319696 322355 319698
rect 321737 319640 321742 319696
rect 321798 319640 322294 319696
rect 322350 319640 322355 319696
rect 321737 319638 322355 319640
rect 321369 319635 321435 319638
rect 321737 319635 321803 319638
rect 322289 319635 322355 319638
rect 322422 319636 322428 319700
rect 322492 319698 322498 319700
rect 322657 319698 322723 319701
rect 322492 319696 322723 319698
rect 322492 319640 322662 319696
rect 322718 319640 322723 319696
rect 322492 319638 322723 319640
rect 322492 319636 322498 319638
rect 322657 319635 322723 319638
rect 323209 319698 323275 319701
rect 324037 319700 324103 319701
rect 323894 319698 323900 319700
rect 323209 319696 323900 319698
rect 323209 319640 323214 319696
rect 323270 319640 323900 319696
rect 323209 319638 323900 319640
rect 323209 319635 323275 319638
rect 323894 319636 323900 319638
rect 323964 319636 323970 319700
rect 324037 319696 324084 319700
rect 324148 319698 324154 319700
rect 324037 319640 324042 319696
rect 324037 319636 324084 319640
rect 324148 319638 324194 319698
rect 324148 319636 324154 319638
rect 324814 319636 324820 319700
rect 324884 319698 324890 319700
rect 324957 319698 325023 319701
rect 330518 319698 330524 319700
rect 324884 319696 330524 319698
rect 324884 319640 324962 319696
rect 325018 319640 330524 319696
rect 324884 319638 330524 319640
rect 324884 319636 324890 319638
rect 324037 319635 324103 319636
rect 324957 319635 325023 319638
rect 330518 319636 330524 319638
rect 330588 319636 330594 319700
rect 333881 319698 333947 319701
rect 362718 319698 362724 319700
rect 333881 319696 362724 319698
rect 333881 319640 333886 319696
rect 333942 319640 362724 319696
rect 333881 319638 362724 319640
rect 333881 319635 333947 319638
rect 362718 319636 362724 319638
rect 362788 319636 362794 319700
rect 318149 319562 318215 319565
rect 318014 319560 318215 319562
rect 318014 319504 318154 319560
rect 318210 319504 318215 319560
rect 318014 319502 318215 319504
rect 317524 319500 317530 319502
rect 317873 319499 317939 319502
rect 318149 319499 318215 319502
rect 321737 319562 321803 319565
rect 322054 319562 322060 319564
rect 321737 319560 322060 319562
rect 321737 319504 321742 319560
rect 321798 319504 322060 319560
rect 321737 319502 322060 319504
rect 321737 319499 321803 319502
rect 322054 319500 322060 319502
rect 322124 319500 322130 319564
rect 322473 319562 322539 319565
rect 326337 319562 326403 319565
rect 322473 319560 326403 319562
rect 322473 319504 322478 319560
rect 322534 319504 326342 319560
rect 326398 319504 326403 319560
rect 322473 319502 326403 319504
rect 322473 319499 322539 319502
rect 326337 319499 326403 319502
rect 326797 319564 326863 319565
rect 326797 319560 326844 319564
rect 326908 319562 326914 319564
rect 327073 319562 327139 319565
rect 367134 319562 367140 319564
rect 326797 319504 326802 319560
rect 326797 319500 326844 319504
rect 326908 319502 326954 319562
rect 327073 319560 367140 319562
rect 327073 319504 327078 319560
rect 327134 319504 367140 319560
rect 327073 319502 367140 319504
rect 326908 319500 326914 319502
rect 326797 319499 326863 319500
rect 327073 319499 327139 319502
rect 367134 319500 367140 319502
rect 367204 319500 367210 319564
rect 318241 319428 318307 319429
rect 302558 319366 317292 319426
rect 318190 319364 318196 319428
rect 318260 319426 318307 319428
rect 318977 319426 319043 319429
rect 320449 319428 320515 319429
rect 319294 319426 319300 319428
rect 318260 319424 318352 319426
rect 318302 319368 318352 319424
rect 318260 319366 318352 319368
rect 318977 319424 319300 319426
rect 318977 319368 318982 319424
rect 319038 319368 319300 319424
rect 318977 319366 319300 319368
rect 318260 319364 318307 319366
rect 318241 319363 318307 319364
rect 318977 319363 319043 319366
rect 319294 319364 319300 319366
rect 319364 319364 319370 319428
rect 320398 319364 320404 319428
rect 320468 319426 320515 319428
rect 320817 319426 320883 319429
rect 321318 319426 321324 319428
rect 320468 319424 320560 319426
rect 320510 319368 320560 319424
rect 320468 319366 320560 319368
rect 320817 319424 321324 319426
rect 320817 319368 320822 319424
rect 320878 319368 321324 319424
rect 320817 319366 321324 319368
rect 320468 319364 320515 319366
rect 320449 319363 320515 319364
rect 320817 319363 320883 319366
rect 321318 319364 321324 319366
rect 321388 319364 321394 319428
rect 321829 319426 321895 319429
rect 329189 319426 329255 319429
rect 321829 319424 329255 319426
rect 321829 319368 321834 319424
rect 321890 319368 329194 319424
rect 329250 319368 329255 319424
rect 321829 319366 329255 319368
rect 321829 319363 321895 319366
rect 329189 319363 329255 319366
rect 3417 319290 3483 319293
rect -960 319288 3483 319290
rect -960 319232 3422 319288
rect 3478 319232 3483 319288
rect -960 319230 3483 319232
rect -960 319140 480 319230
rect 3417 319227 3483 319230
rect 273161 319290 273227 319293
rect 285857 319290 285923 319293
rect 273161 319288 285923 319290
rect 273161 319232 273166 319288
rect 273222 319232 285862 319288
rect 285918 319232 285923 319288
rect 273161 319230 285923 319232
rect 273161 319227 273227 319230
rect 285857 319227 285923 319230
rect 287462 319228 287468 319292
rect 287532 319290 287538 319292
rect 287697 319290 287763 319293
rect 288617 319292 288683 319293
rect 287532 319288 287763 319290
rect 287532 319232 287702 319288
rect 287758 319232 287763 319288
rect 287532 319230 287763 319232
rect 287532 319228 287538 319230
rect 287697 319227 287763 319230
rect 288566 319228 288572 319292
rect 288636 319290 288683 319292
rect 291837 319290 291903 319293
rect 292430 319290 292436 319292
rect 288636 319288 288728 319290
rect 288678 319232 288728 319288
rect 288636 319230 288728 319232
rect 291837 319288 292436 319290
rect 291837 319232 291842 319288
rect 291898 319232 292436 319288
rect 291837 319230 292436 319232
rect 288636 319228 288683 319230
rect 288617 319227 288683 319228
rect 291837 319227 291903 319230
rect 292430 319228 292436 319230
rect 292500 319228 292506 319292
rect 294137 319290 294203 319293
rect 297081 319290 297147 319293
rect 298369 319292 298435 319293
rect 294137 319288 297147 319290
rect 294137 319232 294142 319288
rect 294198 319232 297086 319288
rect 297142 319232 297147 319288
rect 294137 319230 297147 319232
rect 294137 319227 294203 319230
rect 297081 319227 297147 319230
rect 298318 319228 298324 319292
rect 298388 319290 298435 319292
rect 298388 319288 298480 319290
rect 298430 319232 298480 319288
rect 298388 319230 298480 319232
rect 298388 319228 298435 319230
rect 298686 319228 298692 319292
rect 298756 319290 298762 319292
rect 305177 319290 305243 319293
rect 298756 319288 305243 319290
rect 298756 319232 305182 319288
rect 305238 319232 305243 319288
rect 298756 319230 305243 319232
rect 298756 319228 298762 319230
rect 298369 319227 298435 319228
rect 305177 319227 305243 319230
rect 310237 319290 310303 319293
rect 310830 319290 310836 319292
rect 310237 319288 310836 319290
rect 310237 319232 310242 319288
rect 310298 319232 310836 319288
rect 310237 319230 310836 319232
rect 310237 319227 310303 319230
rect 310830 319228 310836 319230
rect 310900 319228 310906 319292
rect 314193 319290 314259 319293
rect 332869 319290 332935 319293
rect 333881 319290 333947 319293
rect 314193 319288 333947 319290
rect 314193 319232 314198 319288
rect 314254 319232 332874 319288
rect 332930 319232 333886 319288
rect 333942 319232 333947 319288
rect 314193 319230 333947 319232
rect 314193 319227 314259 319230
rect 332869 319227 332935 319230
rect 333881 319227 333947 319230
rect 274541 319154 274607 319157
rect 283005 319154 283071 319157
rect 288709 319156 288775 319157
rect 288709 319154 288756 319156
rect 274541 319152 283071 319154
rect 274541 319096 274546 319152
rect 274602 319096 283010 319152
rect 283066 319096 283071 319152
rect 274541 319094 283071 319096
rect 288664 319152 288756 319154
rect 288664 319096 288714 319152
rect 288664 319094 288756 319096
rect 274541 319091 274607 319094
rect 283005 319091 283071 319094
rect 288709 319092 288756 319094
rect 288820 319092 288826 319156
rect 290733 319154 290799 319157
rect 291694 319154 291700 319156
rect 290733 319152 291700 319154
rect 290733 319096 290738 319152
rect 290794 319096 291700 319152
rect 290733 319094 291700 319096
rect 288709 319091 288775 319092
rect 290733 319091 290799 319094
rect 291694 319092 291700 319094
rect 291764 319092 291770 319156
rect 294505 319154 294571 319157
rect 302141 319154 302207 319157
rect 294505 319152 302207 319154
rect 294505 319096 294510 319152
rect 294566 319096 302146 319152
rect 302202 319096 302207 319152
rect 294505 319094 302207 319096
rect 294505 319091 294571 319094
rect 302141 319091 302207 319094
rect 317505 319154 317571 319157
rect 318333 319154 318399 319157
rect 317505 319152 318399 319154
rect 317505 319096 317510 319152
rect 317566 319096 318338 319152
rect 318394 319096 318399 319152
rect 317505 319094 318399 319096
rect 317505 319091 317571 319094
rect 318333 319091 318399 319094
rect 319253 319154 319319 319157
rect 322105 319154 322171 319157
rect 319253 319152 322171 319154
rect 319253 319096 319258 319152
rect 319314 319096 322110 319152
rect 322166 319096 322171 319152
rect 319253 319094 322171 319096
rect 319253 319091 319319 319094
rect 322105 319091 322171 319094
rect 322933 319154 322999 319157
rect 338205 319154 338271 319157
rect 322933 319152 338271 319154
rect 322933 319096 322938 319152
rect 322994 319096 338210 319152
rect 338266 319096 338271 319152
rect 322933 319094 338271 319096
rect 322933 319091 322999 319094
rect 338205 319091 338271 319094
rect 281993 319018 282059 319021
rect 313641 319018 313707 319021
rect 281993 319016 313707 319018
rect 281993 318960 281998 319016
rect 282054 318960 313646 319016
rect 313702 318960 313707 319016
rect 281993 318958 313707 318960
rect 281993 318955 282059 318958
rect 313641 318955 313707 318958
rect 317413 319018 317479 319021
rect 318006 319018 318012 319020
rect 317413 319016 318012 319018
rect 317413 318960 317418 319016
rect 317474 318960 318012 319016
rect 317413 318958 318012 318960
rect 317413 318955 317479 318958
rect 318006 318956 318012 318958
rect 318076 318956 318082 319020
rect 321001 319018 321067 319021
rect 321134 319018 321140 319020
rect 321001 319016 321140 319018
rect 321001 318960 321006 319016
rect 321062 318960 321140 319016
rect 321001 318958 321140 318960
rect 321001 318955 321067 318958
rect 321134 318956 321140 318958
rect 321204 318956 321210 319020
rect 322105 319018 322171 319021
rect 322606 319018 322612 319020
rect 322105 319016 322612 319018
rect 322105 318960 322110 319016
rect 322166 318960 322612 319016
rect 322105 318958 322612 318960
rect 322105 318955 322171 318958
rect 322606 318956 322612 318958
rect 322676 318956 322682 319020
rect 323342 318956 323348 319020
rect 323412 319018 323418 319020
rect 323485 319018 323551 319021
rect 324221 319020 324287 319021
rect 325049 319020 325115 319021
rect 324221 319018 324268 319020
rect 323412 319016 323551 319018
rect 323412 318960 323490 319016
rect 323546 318960 323551 319016
rect 323412 318958 323551 318960
rect 324176 319016 324268 319018
rect 324176 318960 324226 319016
rect 324176 318958 324268 318960
rect 323412 318956 323418 318958
rect 323485 318955 323551 318958
rect 324221 318956 324268 318958
rect 324332 318956 324338 319020
rect 324998 319018 325004 319020
rect 324958 318958 325004 319018
rect 325068 319016 325115 319020
rect 325110 318960 325115 319016
rect 324998 318956 325004 318958
rect 325068 318956 325115 318960
rect 324221 318955 324287 318956
rect 325049 318955 325115 318956
rect 325233 319018 325299 319021
rect 325417 319018 325483 319021
rect 326705 319020 326771 319021
rect 327441 319020 327507 319021
rect 325233 319016 325483 319018
rect 325233 318960 325238 319016
rect 325294 318960 325422 319016
rect 325478 318960 325483 319016
rect 325233 318958 325483 318960
rect 325233 318955 325299 318958
rect 325417 318955 325483 318958
rect 326654 318956 326660 319020
rect 326724 319018 326771 319020
rect 326724 319016 326816 319018
rect 326766 318960 326816 319016
rect 326724 318958 326816 318960
rect 326724 318956 326771 318958
rect 327390 318956 327396 319020
rect 327460 319018 327507 319020
rect 377305 319018 377371 319021
rect 327460 319016 327552 319018
rect 327502 318960 327552 319016
rect 327460 318958 327552 318960
rect 328410 319016 377371 319018
rect 328410 318960 377310 319016
rect 377366 318960 377371 319016
rect 328410 318958 377371 318960
rect 327460 318956 327507 318958
rect 326705 318955 326771 318956
rect 327441 318955 327507 318956
rect 283097 318882 283163 318885
rect 283966 318882 283972 318884
rect 283097 318880 283972 318882
rect 283097 318824 283102 318880
rect 283158 318824 283972 318880
rect 283097 318822 283972 318824
rect 283097 318819 283163 318822
rect 283966 318820 283972 318822
rect 284036 318820 284042 318884
rect 290590 318820 290596 318884
rect 290660 318882 290666 318884
rect 290825 318882 290891 318885
rect 290660 318880 290891 318882
rect 290660 318824 290830 318880
rect 290886 318824 290891 318880
rect 290660 318822 290891 318824
rect 290660 318820 290666 318822
rect 290825 318819 290891 318822
rect 291009 318882 291075 318885
rect 291142 318882 291148 318884
rect 291009 318880 291148 318882
rect 291009 318824 291014 318880
rect 291070 318824 291148 318880
rect 291009 318822 291148 318824
rect 291009 318819 291075 318822
rect 291142 318820 291148 318822
rect 291212 318820 291218 318884
rect 304206 318820 304212 318884
rect 304276 318882 304282 318884
rect 305494 318882 305500 318884
rect 304276 318822 305500 318882
rect 304276 318820 304282 318822
rect 305494 318820 305500 318822
rect 305564 318820 305570 318884
rect 319805 318882 319871 318885
rect 328410 318882 328470 318958
rect 377305 318955 377371 318958
rect 319805 318880 328470 318882
rect 319805 318824 319810 318880
rect 319866 318824 328470 318880
rect 319805 318822 328470 318824
rect 319805 318819 319871 318822
rect 282821 318746 282887 318749
rect 283782 318746 283788 318748
rect 282821 318744 283788 318746
rect 282821 318688 282826 318744
rect 282882 318688 283788 318744
rect 282821 318686 283788 318688
rect 282821 318683 282887 318686
rect 283782 318684 283788 318686
rect 283852 318684 283858 318748
rect 284569 318746 284635 318749
rect 287646 318746 287652 318748
rect 284569 318744 287652 318746
rect 284569 318688 284574 318744
rect 284630 318688 287652 318744
rect 284569 318686 287652 318688
rect 284569 318683 284635 318686
rect 287646 318684 287652 318686
rect 287716 318684 287722 318748
rect 302366 318684 302372 318748
rect 302436 318746 302442 318748
rect 302693 318746 302759 318749
rect 317137 318748 317203 318749
rect 302436 318744 302759 318746
rect 302436 318688 302698 318744
rect 302754 318688 302759 318744
rect 302436 318686 302759 318688
rect 302436 318684 302442 318686
rect 302693 318683 302759 318686
rect 316350 318684 316356 318748
rect 316420 318746 316426 318748
rect 317086 318746 317092 318748
rect 316420 318686 317092 318746
rect 317156 318744 317203 318748
rect 317198 318688 317203 318744
rect 316420 318684 316426 318686
rect 317086 318684 317092 318686
rect 317156 318684 317203 318688
rect 317137 318683 317203 318684
rect 318885 318746 318951 318749
rect 319662 318746 319668 318748
rect 318885 318744 319668 318746
rect 318885 318688 318890 318744
rect 318946 318688 319668 318744
rect 318885 318686 319668 318688
rect 318885 318683 318951 318686
rect 319662 318684 319668 318686
rect 319732 318684 319738 318748
rect 324497 318746 324563 318749
rect 329741 318746 329807 318749
rect 324497 318744 329807 318746
rect 324497 318688 324502 318744
rect 324558 318688 329746 318744
rect 329802 318688 329807 318744
rect 324497 318686 329807 318688
rect 324497 318683 324563 318686
rect 329741 318683 329807 318686
rect 227161 318610 227227 318613
rect 283414 318610 283420 318612
rect 227161 318608 283420 318610
rect 227161 318552 227166 318608
rect 227222 318552 283420 318608
rect 227161 318550 283420 318552
rect 227161 318547 227227 318550
rect 283414 318548 283420 318550
rect 283484 318548 283490 318612
rect 285397 318610 285463 318613
rect 288934 318610 288940 318612
rect 285397 318608 288940 318610
rect 285397 318552 285402 318608
rect 285458 318552 288940 318608
rect 285397 318550 288940 318552
rect 285397 318547 285463 318550
rect 288934 318548 288940 318550
rect 289004 318548 289010 318612
rect 297081 318610 297147 318613
rect 302550 318610 302556 318612
rect 297081 318608 302556 318610
rect 297081 318552 297086 318608
rect 297142 318552 302556 318608
rect 297081 318550 302556 318552
rect 297081 318547 297147 318550
rect 302550 318548 302556 318550
rect 302620 318548 302626 318612
rect 309358 318548 309364 318612
rect 309428 318610 309434 318612
rect 309501 318610 309567 318613
rect 310094 318610 310100 318612
rect 309428 318608 310100 318610
rect 309428 318552 309506 318608
rect 309562 318552 310100 318608
rect 309428 318550 310100 318552
rect 309428 318548 309434 318550
rect 309501 318547 309567 318550
rect 310094 318548 310100 318550
rect 310164 318548 310170 318612
rect 316861 318610 316927 318613
rect 317137 318610 317203 318613
rect 316861 318608 317203 318610
rect 316861 318552 316866 318608
rect 316922 318552 317142 318608
rect 317198 318552 317203 318608
rect 316861 318550 317203 318552
rect 316861 318547 316927 318550
rect 317137 318547 317203 318550
rect 319897 318610 319963 318613
rect 328494 318610 328500 318612
rect 319897 318608 328500 318610
rect 319897 318552 319902 318608
rect 319958 318552 328500 318608
rect 319897 318550 328500 318552
rect 319897 318547 319963 318550
rect 328494 318548 328500 318550
rect 328564 318548 328570 318612
rect 329649 318610 329715 318613
rect 331305 318610 331371 318613
rect 329649 318608 331371 318610
rect 329649 318552 329654 318608
rect 329710 318552 331310 318608
rect 331366 318552 331371 318608
rect 329649 318550 331371 318552
rect 329649 318547 329715 318550
rect 331305 318547 331371 318550
rect 233325 318474 233391 318477
rect 284334 318474 284340 318476
rect 233325 318472 284340 318474
rect 233325 318416 233330 318472
rect 233386 318416 284340 318472
rect 233325 318414 284340 318416
rect 233325 318411 233391 318414
rect 284334 318412 284340 318414
rect 284404 318412 284410 318476
rect 294229 318474 294295 318477
rect 316861 318476 316927 318477
rect 294454 318474 294460 318476
rect 294229 318472 294460 318474
rect 294229 318416 294234 318472
rect 294290 318416 294460 318472
rect 294229 318414 294460 318416
rect 294229 318411 294295 318414
rect 294454 318412 294460 318414
rect 294524 318412 294530 318476
rect 316861 318474 316908 318476
rect 316816 318472 316908 318474
rect 316816 318416 316866 318472
rect 316816 318414 316908 318416
rect 316861 318412 316908 318414
rect 316972 318412 316978 318476
rect 323342 318412 323348 318476
rect 323412 318474 323418 318476
rect 324037 318474 324103 318477
rect 323412 318472 324103 318474
rect 323412 318416 324042 318472
rect 324098 318416 324103 318472
rect 323412 318414 324103 318416
rect 323412 318412 323418 318414
rect 316861 318411 316927 318412
rect 324037 318411 324103 318414
rect 247534 318276 247540 318340
rect 247604 318338 247610 318340
rect 285438 318338 285444 318340
rect 247604 318278 285444 318338
rect 247604 318276 247610 318278
rect 285438 318276 285444 318278
rect 285508 318276 285514 318340
rect 289302 318338 289308 318340
rect 288022 318278 289308 318338
rect 269849 318202 269915 318205
rect 288022 318202 288082 318278
rect 289302 318276 289308 318278
rect 289372 318338 289378 318340
rect 289629 318338 289695 318341
rect 289372 318336 289695 318338
rect 289372 318280 289634 318336
rect 289690 318280 289695 318336
rect 289372 318278 289695 318280
rect 289372 318276 289378 318278
rect 289629 318275 289695 318278
rect 290089 318338 290155 318341
rect 297173 318338 297239 318341
rect 290089 318336 297239 318338
rect 290089 318280 290094 318336
rect 290150 318280 297178 318336
rect 297234 318280 297239 318336
rect 290089 318278 297239 318280
rect 290089 318275 290155 318278
rect 297173 318275 297239 318278
rect 306414 318276 306420 318340
rect 306484 318338 306490 318340
rect 307477 318338 307543 318341
rect 306484 318336 307543 318338
rect 306484 318280 307482 318336
rect 307538 318280 307543 318336
rect 306484 318278 307543 318280
rect 306484 318276 306490 318278
rect 307477 318275 307543 318278
rect 321553 318338 321619 318341
rect 329189 318338 329255 318341
rect 321553 318336 329255 318338
rect 321553 318280 321558 318336
rect 321614 318280 329194 318336
rect 329250 318280 329255 318336
rect 321553 318278 329255 318280
rect 321553 318275 321619 318278
rect 329189 318275 329255 318278
rect 292021 318204 292087 318205
rect 292021 318202 292068 318204
rect 269849 318200 288082 318202
rect 269849 318144 269854 318200
rect 269910 318144 288082 318200
rect 269849 318142 288082 318144
rect 291976 318200 292068 318202
rect 291976 318144 292026 318200
rect 291976 318142 292068 318144
rect 269849 318139 269915 318142
rect 292021 318140 292068 318142
rect 292132 318140 292138 318204
rect 302325 318202 302391 318205
rect 292530 318200 302391 318202
rect 292530 318144 302330 318200
rect 302386 318144 302391 318200
rect 292530 318142 302391 318144
rect 292021 318139 292087 318140
rect 237966 318004 237972 318068
rect 238036 318066 238042 318068
rect 259177 318066 259243 318069
rect 238036 318064 259243 318066
rect 238036 318008 259182 318064
rect 259238 318008 259243 318064
rect 238036 318006 259243 318008
rect 238036 318004 238042 318006
rect 259177 318003 259243 318006
rect 291326 318004 291332 318068
rect 291396 318066 291402 318068
rect 292530 318066 292590 318142
rect 302325 318139 302391 318142
rect 323485 318202 323551 318205
rect 331489 318202 331555 318205
rect 332317 318202 332383 318205
rect 323485 318200 332383 318202
rect 323485 318144 323490 318200
rect 323546 318144 331494 318200
rect 331550 318144 332322 318200
rect 332378 318144 332383 318200
rect 323485 318142 332383 318144
rect 323485 318139 323551 318142
rect 331489 318139 331555 318142
rect 332317 318139 332383 318142
rect 291396 318006 292590 318066
rect 299289 318066 299355 318069
rect 299422 318066 299428 318068
rect 299289 318064 299428 318066
rect 299289 318008 299294 318064
rect 299350 318008 299428 318064
rect 299289 318006 299428 318008
rect 291396 318004 291402 318006
rect 299289 318003 299355 318006
rect 299422 318004 299428 318006
rect 299492 318004 299498 318068
rect 303470 318004 303476 318068
rect 303540 318066 303546 318068
rect 304533 318066 304599 318069
rect 303540 318064 304599 318066
rect 303540 318008 304538 318064
rect 304594 318008 304599 318064
rect 303540 318006 304599 318008
rect 303540 318004 303546 318006
rect 304533 318003 304599 318006
rect 318742 318004 318748 318068
rect 318812 318066 318818 318068
rect 318885 318066 318951 318069
rect 318812 318064 318951 318066
rect 318812 318008 318890 318064
rect 318946 318008 318951 318064
rect 318812 318006 318951 318008
rect 318812 318004 318818 318006
rect 318885 318003 318951 318006
rect 324037 318066 324103 318069
rect 329373 318066 329439 318069
rect 324037 318064 329439 318066
rect 324037 318008 324042 318064
rect 324098 318008 329378 318064
rect 329434 318008 329439 318064
rect 324037 318006 329439 318008
rect 324037 318003 324103 318006
rect 329373 318003 329439 318006
rect 329925 318066 329991 318069
rect 369894 318066 369900 318068
rect 329925 318064 369900 318066
rect 329925 318008 329930 318064
rect 329986 318008 369900 318064
rect 329925 318006 369900 318008
rect 329925 318003 329991 318006
rect 369894 318004 369900 318006
rect 369964 318004 369970 318068
rect 279601 317930 279667 317933
rect 280705 317930 280771 317933
rect 298185 317932 298251 317933
rect 279601 317928 292590 317930
rect 279601 317872 279606 317928
rect 279662 317872 280710 317928
rect 280766 317872 292590 317928
rect 279601 317870 292590 317872
rect 279601 317867 279667 317870
rect 280705 317867 280771 317870
rect 283230 317732 283236 317796
rect 283300 317794 283306 317796
rect 284017 317794 284083 317797
rect 283300 317792 284083 317794
rect 283300 317736 284022 317792
rect 284078 317736 284083 317792
rect 283300 317734 284083 317736
rect 283300 317732 283306 317734
rect 284017 317731 284083 317734
rect 284385 317794 284451 317797
rect 285397 317794 285463 317797
rect 284385 317792 285463 317794
rect 284385 317736 284390 317792
rect 284446 317736 285402 317792
rect 285458 317736 285463 317792
rect 284385 317734 285463 317736
rect 284385 317731 284451 317734
rect 285397 317731 285463 317734
rect 291142 317732 291148 317796
rect 291212 317794 291218 317796
rect 291837 317794 291903 317797
rect 291212 317792 291903 317794
rect 291212 317736 291842 317792
rect 291898 317736 291903 317792
rect 291212 317734 291903 317736
rect 292530 317794 292590 317870
rect 298134 317868 298140 317932
rect 298204 317930 298251 317932
rect 298204 317928 298296 317930
rect 298246 317872 298296 317928
rect 298204 317870 298296 317872
rect 298204 317868 298251 317870
rect 299606 317868 299612 317932
rect 299676 317930 299682 317932
rect 300301 317930 300367 317933
rect 299676 317928 300367 317930
rect 299676 317872 300306 317928
rect 300362 317872 300367 317928
rect 299676 317870 300367 317872
rect 299676 317868 299682 317870
rect 298185 317867 298251 317868
rect 300301 317867 300367 317870
rect 302734 317868 302740 317932
rect 302804 317930 302810 317932
rect 303061 317930 303127 317933
rect 302804 317928 303127 317930
rect 302804 317872 303066 317928
rect 303122 317872 303127 317928
rect 302804 317870 303127 317872
rect 302804 317868 302810 317870
rect 303061 317867 303127 317870
rect 304257 317930 304323 317933
rect 304574 317930 304580 317932
rect 304257 317928 304580 317930
rect 304257 317872 304262 317928
rect 304318 317872 304580 317928
rect 304257 317870 304580 317872
rect 304257 317867 304323 317870
rect 304574 317868 304580 317870
rect 304644 317868 304650 317932
rect 306966 317868 306972 317932
rect 307036 317930 307042 317932
rect 307201 317930 307267 317933
rect 307036 317928 307267 317930
rect 307036 317872 307206 317928
rect 307262 317872 307267 317928
rect 307036 317870 307267 317872
rect 307036 317868 307042 317870
rect 307201 317867 307267 317870
rect 311750 317868 311756 317932
rect 311820 317930 311826 317932
rect 313365 317930 313431 317933
rect 313825 317932 313891 317933
rect 311820 317928 313431 317930
rect 311820 317872 313370 317928
rect 313426 317872 313431 317928
rect 311820 317870 313431 317872
rect 311820 317868 311826 317870
rect 313365 317867 313431 317870
rect 313774 317868 313780 317932
rect 313844 317930 313891 317932
rect 314009 317930 314075 317933
rect 315573 317930 315639 317933
rect 320766 317930 320772 317932
rect 313844 317928 313936 317930
rect 313886 317872 313936 317928
rect 313844 317870 313936 317872
rect 314009 317928 315639 317930
rect 314009 317872 314014 317928
rect 314070 317872 315578 317928
rect 315634 317872 315639 317928
rect 314009 317870 315639 317872
rect 313844 317868 313891 317870
rect 313825 317867 313891 317868
rect 314009 317867 314075 317870
rect 315573 317867 315639 317870
rect 320038 317870 320772 317930
rect 313273 317794 313339 317797
rect 320038 317794 320098 317870
rect 320766 317868 320772 317870
rect 320836 317868 320842 317932
rect 320909 317930 320975 317933
rect 323209 317932 323275 317933
rect 320909 317928 321570 317930
rect 320909 317872 320914 317928
rect 320970 317872 321570 317928
rect 320909 317870 321570 317872
rect 320909 317867 320975 317870
rect 292530 317792 313339 317794
rect 292530 317736 313278 317792
rect 313334 317736 313339 317792
rect 292530 317734 313339 317736
rect 291212 317732 291218 317734
rect 291837 317731 291903 317734
rect 313273 317731 313339 317734
rect 315990 317734 320098 317794
rect 283281 317658 283347 317661
rect 273210 317656 283347 317658
rect 273210 317600 283286 317656
rect 283342 317600 283347 317656
rect 273210 317598 283347 317600
rect 225781 317522 225847 317525
rect 273210 317522 273270 317598
rect 283281 317595 283347 317598
rect 297173 317658 297239 317661
rect 315990 317658 316050 317734
rect 320214 317732 320220 317796
rect 320284 317794 320290 317796
rect 321001 317794 321067 317797
rect 320284 317792 321067 317794
rect 320284 317736 321006 317792
rect 321062 317736 321067 317792
rect 320284 317734 321067 317736
rect 321510 317794 321570 317870
rect 323158 317868 323164 317932
rect 323228 317930 323275 317932
rect 328913 317930 328979 317933
rect 329046 317930 329052 317932
rect 323228 317928 323320 317930
rect 323270 317872 323320 317928
rect 323228 317870 323320 317872
rect 328913 317928 329052 317930
rect 328913 317872 328918 317928
rect 328974 317872 329052 317928
rect 328913 317870 329052 317872
rect 323228 317868 323275 317870
rect 323209 317867 323275 317868
rect 328913 317867 328979 317870
rect 329046 317868 329052 317870
rect 329116 317868 329122 317932
rect 326654 317794 326660 317796
rect 321510 317734 326660 317794
rect 320284 317732 320290 317734
rect 321001 317731 321067 317734
rect 326654 317732 326660 317734
rect 326724 317732 326730 317796
rect 327257 317794 327323 317797
rect 327993 317794 328059 317797
rect 328310 317794 328316 317796
rect 327257 317792 328316 317794
rect 327257 317736 327262 317792
rect 327318 317736 327998 317792
rect 328054 317736 328316 317792
rect 327257 317734 328316 317736
rect 327257 317731 327323 317734
rect 327993 317731 328059 317734
rect 328310 317732 328316 317734
rect 328380 317732 328386 317796
rect 297173 317656 316050 317658
rect 297173 317600 297178 317656
rect 297234 317600 316050 317656
rect 297173 317598 316050 317600
rect 316125 317658 316191 317661
rect 317270 317658 317276 317660
rect 316125 317656 317276 317658
rect 316125 317600 316130 317656
rect 316186 317600 317276 317656
rect 316125 317598 317276 317600
rect 297173 317595 297239 317598
rect 316125 317595 316191 317598
rect 317270 317596 317276 317598
rect 317340 317596 317346 317660
rect 326613 317658 326679 317661
rect 327022 317658 327028 317660
rect 326613 317656 327028 317658
rect 326613 317600 326618 317656
rect 326674 317600 327028 317656
rect 326613 317598 327028 317600
rect 326613 317595 326679 317598
rect 327022 317596 327028 317598
rect 327092 317596 327098 317660
rect 329741 317658 329807 317661
rect 332685 317658 332751 317661
rect 329741 317656 332751 317658
rect 329741 317600 329746 317656
rect 329802 317600 332690 317656
rect 332746 317600 332751 317656
rect 329741 317598 332751 317600
rect 329741 317595 329807 317598
rect 332685 317595 332751 317598
rect 225781 317520 273270 317522
rect 225781 317464 225786 317520
rect 225842 317464 273270 317520
rect 225781 317462 273270 317464
rect 225781 317459 225847 317462
rect 283046 317460 283052 317524
rect 283116 317522 283122 317524
rect 283649 317522 283715 317525
rect 283116 317520 283715 317522
rect 283116 317464 283654 317520
rect 283710 317464 283715 317520
rect 283116 317462 283715 317464
rect 283116 317460 283122 317462
rect 283649 317459 283715 317462
rect 289169 317522 289235 317525
rect 290089 317522 290155 317525
rect 289169 317520 290155 317522
rect 289169 317464 289174 317520
rect 289230 317464 290094 317520
rect 290150 317464 290155 317520
rect 289169 317462 290155 317464
rect 289169 317459 289235 317462
rect 290089 317459 290155 317462
rect 293677 317522 293743 317525
rect 295926 317522 295932 317524
rect 293677 317520 295932 317522
rect 293677 317464 293682 317520
rect 293738 317464 295932 317520
rect 293677 317462 295932 317464
rect 293677 317459 293743 317462
rect 295926 317460 295932 317462
rect 295996 317460 296002 317524
rect 297081 317522 297147 317525
rect 297725 317522 297791 317525
rect 297081 317520 297791 317522
rect 297081 317464 297086 317520
rect 297142 317464 297730 317520
rect 297786 317464 297791 317520
rect 297081 317462 297791 317464
rect 297081 317459 297147 317462
rect 297725 317459 297791 317462
rect 299422 317460 299428 317524
rect 299492 317522 299498 317524
rect 300025 317522 300091 317525
rect 299492 317520 300091 317522
rect 299492 317464 300030 317520
rect 300086 317464 300091 317520
rect 299492 317462 300091 317464
rect 299492 317460 299498 317462
rect 300025 317459 300091 317462
rect 301078 317460 301084 317524
rect 301148 317522 301154 317524
rect 301957 317522 302023 317525
rect 301148 317520 302023 317522
rect 301148 317464 301962 317520
rect 302018 317464 302023 317520
rect 301148 317462 302023 317464
rect 301148 317460 301154 317462
rect 301957 317459 302023 317462
rect 302918 317460 302924 317524
rect 302988 317522 302994 317524
rect 303245 317522 303311 317525
rect 304441 317524 304507 317525
rect 304390 317522 304396 317524
rect 302988 317520 303311 317522
rect 302988 317464 303250 317520
rect 303306 317464 303311 317520
rect 302988 317462 303311 317464
rect 304350 317462 304396 317522
rect 304460 317520 304507 317524
rect 304502 317464 304507 317520
rect 302988 317460 302994 317462
rect 303245 317459 303311 317462
rect 304390 317460 304396 317462
rect 304460 317460 304507 317464
rect 304441 317459 304507 317460
rect 306741 317522 306807 317525
rect 307518 317522 307524 317524
rect 306741 317520 307524 317522
rect 306741 317464 306746 317520
rect 306802 317464 307524 317520
rect 306741 317462 307524 317464
rect 306741 317459 306807 317462
rect 307518 317460 307524 317462
rect 307588 317460 307594 317524
rect 312537 317522 312603 317525
rect 312670 317522 312676 317524
rect 312537 317520 312676 317522
rect 312537 317464 312542 317520
rect 312598 317464 312676 317520
rect 312537 317462 312676 317464
rect 312537 317459 312603 317462
rect 312670 317460 312676 317462
rect 312740 317460 312746 317524
rect 315614 317460 315620 317524
rect 315684 317522 315690 317524
rect 315757 317522 315823 317525
rect 315684 317520 315823 317522
rect 315684 317464 315762 317520
rect 315818 317464 315823 317520
rect 315684 317462 315823 317464
rect 315684 317460 315690 317462
rect 315757 317459 315823 317462
rect 316534 317460 316540 317524
rect 316604 317522 316610 317524
rect 317229 317522 317295 317525
rect 318425 317524 318491 317525
rect 318374 317522 318380 317524
rect 316604 317520 317295 317522
rect 316604 317464 317234 317520
rect 317290 317464 317295 317520
rect 316604 317462 317295 317464
rect 318334 317462 318380 317522
rect 318444 317520 318491 317524
rect 318486 317464 318491 317520
rect 316604 317460 316610 317462
rect 317229 317459 317295 317462
rect 318374 317460 318380 317462
rect 318444 317460 318491 317464
rect 318425 317459 318491 317460
rect 320265 317522 320331 317525
rect 321318 317522 321324 317524
rect 320265 317520 321324 317522
rect 320265 317464 320270 317520
rect 320326 317464 321324 317520
rect 320265 317462 321324 317464
rect 320265 317459 320331 317462
rect 321318 317460 321324 317462
rect 321388 317460 321394 317524
rect 321686 317460 321692 317524
rect 321756 317522 321762 317524
rect 322197 317522 322263 317525
rect 321756 317520 322263 317522
rect 321756 317464 322202 317520
rect 322258 317464 322263 317520
rect 321756 317462 322263 317464
rect 321756 317460 321762 317462
rect 322197 317459 322263 317462
rect 326981 317522 327047 317525
rect 334985 317522 335051 317525
rect 326981 317520 335051 317522
rect 326981 317464 326986 317520
rect 327042 317464 334990 317520
rect 335046 317464 335051 317520
rect 326981 317462 335051 317464
rect 326981 317459 327047 317462
rect 334985 317459 335051 317462
rect 266353 317386 266419 317389
rect 267549 317386 267615 317389
rect 289353 317386 289419 317389
rect 266353 317384 289419 317386
rect 266353 317328 266358 317384
rect 266414 317328 267554 317384
rect 267610 317328 289358 317384
rect 289414 317328 289419 317384
rect 266353 317326 289419 317328
rect 266353 317323 266419 317326
rect 267549 317323 267615 317326
rect 289353 317323 289419 317326
rect 324865 317386 324931 317389
rect 390921 317386 390987 317389
rect 324865 317384 390987 317386
rect 324865 317328 324870 317384
rect 324926 317328 390926 317384
rect 390982 317328 390987 317384
rect 324865 317326 390987 317328
rect 324865 317323 324931 317326
rect 390921 317323 390987 317326
rect 272977 317250 273043 317253
rect 284201 317250 284267 317253
rect 272977 317248 284267 317250
rect 272977 317192 272982 317248
rect 273038 317192 284206 317248
rect 284262 317192 284267 317248
rect 272977 317190 284267 317192
rect 272977 317187 273043 317190
rect 284201 317187 284267 317190
rect 325233 317250 325299 317253
rect 385677 317250 385743 317253
rect 325233 317248 385743 317250
rect 325233 317192 325238 317248
rect 325294 317192 385682 317248
rect 385738 317192 385743 317248
rect 325233 317190 385743 317192
rect 325233 317187 325299 317190
rect 385677 317187 385743 317190
rect 272793 317114 272859 317117
rect 317045 317114 317111 317117
rect 272793 317112 317111 317114
rect 272793 317056 272798 317112
rect 272854 317056 317050 317112
rect 317106 317056 317111 317112
rect 272793 317054 317111 317056
rect 272793 317051 272859 317054
rect 317045 317051 317111 317054
rect 326797 317114 326863 317117
rect 386505 317114 386571 317117
rect 326797 317112 386571 317114
rect 326797 317056 326802 317112
rect 326858 317056 386510 317112
rect 386566 317056 386571 317112
rect 326797 317054 386571 317056
rect 326797 317051 326863 317054
rect 386505 317051 386571 317054
rect 223430 316916 223436 316980
rect 223500 316978 223506 316980
rect 242525 316978 242591 316981
rect 223500 316976 242591 316978
rect 223500 316920 242530 316976
rect 242586 316920 242591 316976
rect 223500 316918 242591 316920
rect 223500 316916 223506 316918
rect 242525 316915 242591 316918
rect 306966 316916 306972 316980
rect 307036 316978 307042 316980
rect 366398 316978 366404 316980
rect 307036 316918 366404 316978
rect 307036 316916 307042 316918
rect 366398 316916 366404 316918
rect 366468 316916 366474 316980
rect 231710 316780 231716 316844
rect 231780 316842 231786 316844
rect 290733 316842 290799 316845
rect 231780 316840 290799 316842
rect 231780 316784 290738 316840
rect 290794 316784 290799 316840
rect 231780 316782 290799 316784
rect 231780 316780 231786 316782
rect 290733 316779 290799 316782
rect 322381 316842 322447 316845
rect 322381 316840 331230 316842
rect 322381 316784 322386 316840
rect 322442 316784 331230 316840
rect 322381 316782 331230 316784
rect 322381 316779 322447 316782
rect 206829 316706 206895 316709
rect 272241 316706 272307 316709
rect 272977 316706 273043 316709
rect 206829 316704 273043 316706
rect 206829 316648 206834 316704
rect 206890 316648 272246 316704
rect 272302 316648 272982 316704
rect 273038 316648 273043 316704
rect 206829 316646 273043 316648
rect 206829 316643 206895 316646
rect 272241 316643 272307 316646
rect 272977 316643 273043 316646
rect 296897 316706 296963 316709
rect 297950 316706 297956 316708
rect 296897 316704 297956 316706
rect 296897 316648 296902 316704
rect 296958 316648 297956 316704
rect 296897 316646 297956 316648
rect 296897 316643 296963 316646
rect 297950 316644 297956 316646
rect 298020 316644 298026 316708
rect 303061 316706 303127 316709
rect 319110 316706 319116 316708
rect 303061 316704 319116 316706
rect 303061 316648 303066 316704
rect 303122 316648 319116 316704
rect 303061 316646 319116 316648
rect 303061 316643 303127 316646
rect 319110 316644 319116 316646
rect 319180 316644 319186 316708
rect 326889 316706 326955 316709
rect 328453 316706 328519 316709
rect 326889 316704 328519 316706
rect 326889 316648 326894 316704
rect 326950 316648 328458 316704
rect 328514 316648 328519 316704
rect 326889 316646 328519 316648
rect 331170 316706 331230 316782
rect 339585 316706 339651 316709
rect 340505 316706 340571 316709
rect 331170 316704 340571 316706
rect 331170 316648 339590 316704
rect 339646 316648 340510 316704
rect 340566 316648 340571 316704
rect 331170 316646 340571 316648
rect 326889 316643 326955 316646
rect 328453 316643 328519 316646
rect 339585 316643 339651 316646
rect 340505 316643 340571 316646
rect 338205 316570 338271 316573
rect 338614 316570 338620 316572
rect 331170 316568 338620 316570
rect 331170 316512 338210 316568
rect 338266 316512 338620 316568
rect 331170 316510 338620 316512
rect 276933 316434 276999 316437
rect 303245 316434 303311 316437
rect 276933 316432 303311 316434
rect 276933 316376 276938 316432
rect 276994 316376 303250 316432
rect 303306 316376 303311 316432
rect 276933 316374 303311 316376
rect 276933 316371 276999 316374
rect 303245 316371 303311 316374
rect 326654 316372 326660 316436
rect 326724 316434 326730 316436
rect 331170 316434 331230 316510
rect 338205 316507 338271 316510
rect 338614 316508 338620 316510
rect 338684 316508 338690 316572
rect 326724 316374 331230 316434
rect 326724 316372 326730 316374
rect 272977 316298 273043 316301
rect 304901 316298 304967 316301
rect 272977 316296 304967 316298
rect 272977 316240 272982 316296
rect 273038 316240 304906 316296
rect 304962 316240 304967 316296
rect 272977 316238 304967 316240
rect 272977 316235 273043 316238
rect 304901 316235 304967 316238
rect 326613 316298 326679 316301
rect 326797 316298 326863 316301
rect 326613 316296 326863 316298
rect 326613 316240 326618 316296
rect 326674 316240 326802 316296
rect 326858 316240 326863 316296
rect 326613 316238 326863 316240
rect 326613 316235 326679 316238
rect 326797 316235 326863 316238
rect 328862 316236 328868 316300
rect 328932 316298 328938 316300
rect 329189 316298 329255 316301
rect 328932 316296 329255 316298
rect 328932 316240 329194 316296
rect 329250 316240 329255 316296
rect 328932 316238 329255 316240
rect 328932 316236 328938 316238
rect 329189 316235 329255 316238
rect 273805 316162 273871 316165
rect 320173 316162 320239 316165
rect 273805 316160 320239 316162
rect 273805 316104 273810 316160
rect 273866 316104 320178 316160
rect 320234 316104 320239 316160
rect 273805 316102 320239 316104
rect 273805 316099 273871 316102
rect 320173 316099 320239 316102
rect 328678 316100 328684 316164
rect 328748 316162 328754 316164
rect 329373 316162 329439 316165
rect 328748 316160 329439 316162
rect 328748 316104 329378 316160
rect 329434 316104 329439 316160
rect 328748 316102 329439 316104
rect 328748 316100 328754 316102
rect 329373 316099 329439 316102
rect 238569 316026 238635 316029
rect 271781 316026 271847 316029
rect 238569 316024 271847 316026
rect 238569 315968 238574 316024
rect 238630 315968 271786 316024
rect 271842 315968 271847 316024
rect 238569 315966 271847 315968
rect 238569 315963 238635 315966
rect 271781 315963 271847 315966
rect 294413 316026 294479 316029
rect 295190 316026 295196 316028
rect 294413 316024 295196 316026
rect 294413 315968 294418 316024
rect 294474 315968 295196 316024
rect 294413 315966 295196 315968
rect 294413 315963 294479 315966
rect 295190 315964 295196 315966
rect 295260 315964 295266 316028
rect 314101 316026 314167 316029
rect 333605 316026 333671 316029
rect 314101 316024 333671 316026
rect 314101 315968 314106 316024
rect 314162 315968 333610 316024
rect 333666 315968 333671 316024
rect 314101 315966 333671 315968
rect 314101 315963 314167 315966
rect 333605 315963 333671 315966
rect 237230 315828 237236 315892
rect 237300 315890 237306 315892
rect 296478 315890 296484 315892
rect 237300 315830 296484 315890
rect 237300 315828 237306 315830
rect 296478 315828 296484 315830
rect 296548 315828 296554 315892
rect 301497 315890 301563 315893
rect 360142 315890 360148 315892
rect 301497 315888 360148 315890
rect 301497 315832 301502 315888
rect 301558 315832 360148 315888
rect 301497 315830 360148 315832
rect 301497 315827 301563 315830
rect 360142 315828 360148 315830
rect 360212 315828 360218 315892
rect 235206 315692 235212 315756
rect 235276 315754 235282 315756
rect 288157 315754 288223 315757
rect 235276 315752 288223 315754
rect 235276 315696 288162 315752
rect 288218 315696 288223 315752
rect 235276 315694 288223 315696
rect 235276 315692 235282 315694
rect 288157 315691 288223 315694
rect 291193 315754 291259 315757
rect 291326 315754 291332 315756
rect 291193 315752 291332 315754
rect 291193 315696 291198 315752
rect 291254 315696 291332 315752
rect 291193 315694 291332 315696
rect 291193 315691 291259 315694
rect 291326 315692 291332 315694
rect 291396 315692 291402 315756
rect 294689 315754 294755 315757
rect 296846 315754 296852 315756
rect 294689 315752 296852 315754
rect 294689 315696 294694 315752
rect 294750 315696 296852 315752
rect 294689 315694 296852 315696
rect 294689 315691 294755 315694
rect 296846 315692 296852 315694
rect 296916 315692 296922 315756
rect 301630 315692 301636 315756
rect 301700 315754 301706 315756
rect 301773 315754 301839 315757
rect 301700 315752 301839 315754
rect 301700 315696 301778 315752
rect 301834 315696 301839 315752
rect 301700 315694 301839 315696
rect 301700 315692 301706 315694
rect 301773 315691 301839 315694
rect 320817 315754 320883 315757
rect 321001 315754 321067 315757
rect 379605 315754 379671 315757
rect 320817 315752 379671 315754
rect 320817 315696 320822 315752
rect 320878 315696 321006 315752
rect 321062 315696 379610 315752
rect 379666 315696 379671 315752
rect 320817 315694 379671 315696
rect 320817 315691 320883 315694
rect 321001 315691 321067 315694
rect 379605 315691 379671 315694
rect 224718 315556 224724 315620
rect 224788 315618 224794 315620
rect 233325 315618 233391 315621
rect 224788 315616 233391 315618
rect 224788 315560 233330 315616
rect 233386 315560 233391 315616
rect 224788 315558 233391 315560
rect 224788 315556 224794 315558
rect 233325 315555 233391 315558
rect 237046 315556 237052 315620
rect 237116 315618 237122 315620
rect 297030 315618 297036 315620
rect 237116 315558 297036 315618
rect 237116 315556 237122 315558
rect 297030 315556 297036 315558
rect 297100 315556 297106 315620
rect 301405 315618 301471 315621
rect 314142 315618 314148 315620
rect 301405 315616 314148 315618
rect 301405 315560 301410 315616
rect 301466 315560 314148 315616
rect 301405 315558 314148 315560
rect 301405 315555 301471 315558
rect 314142 315556 314148 315558
rect 314212 315556 314218 315620
rect 326153 315618 326219 315621
rect 382774 315618 382780 315620
rect 326153 315616 382780 315618
rect 326153 315560 326158 315616
rect 326214 315560 382780 315616
rect 326153 315558 382780 315560
rect 326153 315555 326219 315558
rect 382774 315556 382780 315558
rect 382844 315556 382850 315620
rect 217777 315482 217843 315485
rect 294689 315482 294755 315485
rect 296110 315482 296116 315484
rect 217777 315480 294755 315482
rect 217777 315424 217782 315480
rect 217838 315424 294694 315480
rect 294750 315424 294755 315480
rect 217777 315422 294755 315424
rect 217777 315419 217843 315422
rect 294689 315419 294755 315422
rect 295290 315422 296116 315482
rect 212349 315346 212415 315349
rect 295290 315346 295350 315422
rect 296110 315420 296116 315422
rect 296180 315420 296186 315484
rect 312353 315482 312419 315485
rect 334065 315482 334131 315485
rect 335169 315482 335235 315485
rect 312353 315480 335235 315482
rect 312353 315424 312358 315480
rect 312414 315424 334070 315480
rect 334126 315424 335174 315480
rect 335230 315424 335235 315480
rect 312353 315422 335235 315424
rect 312353 315419 312419 315422
rect 334065 315419 334131 315422
rect 335169 315419 335235 315422
rect 212349 315344 295350 315346
rect 212349 315288 212354 315344
rect 212410 315288 295350 315344
rect 212349 315286 295350 315288
rect 212349 315283 212415 315286
rect 295926 315284 295932 315348
rect 295996 315346 296002 315348
rect 316718 315346 316724 315348
rect 295996 315286 316724 315346
rect 295996 315284 296002 315286
rect 316718 315284 316724 315286
rect 316788 315284 316794 315348
rect 327349 315346 327415 315349
rect 339217 315346 339283 315349
rect 327349 315344 339283 315346
rect 327349 315288 327354 315344
rect 327410 315288 339222 315344
rect 339278 315288 339283 315344
rect 327349 315286 339283 315288
rect 327349 315283 327415 315286
rect 339217 315283 339283 315286
rect 278037 315210 278103 315213
rect 301497 315210 301563 315213
rect 278037 315208 301563 315210
rect 278037 315152 278042 315208
rect 278098 315152 301502 315208
rect 301558 315152 301563 315208
rect 278037 315150 301563 315152
rect 278037 315147 278103 315150
rect 301497 315147 301563 315150
rect 319437 315210 319503 315213
rect 319989 315210 320055 315213
rect 390829 315210 390895 315213
rect 319437 315208 390895 315210
rect 319437 315152 319442 315208
rect 319498 315152 319994 315208
rect 320050 315152 390834 315208
rect 390890 315152 390895 315208
rect 319437 315150 390895 315152
rect 319437 315147 319503 315150
rect 319989 315147 320055 315150
rect 390829 315147 390895 315150
rect 271781 315074 271847 315077
rect 299238 315074 299244 315076
rect 271781 315072 299244 315074
rect 271781 315016 271786 315072
rect 271842 315016 299244 315072
rect 271781 315014 299244 315016
rect 271781 315011 271847 315014
rect 299238 315012 299244 315014
rect 299308 315012 299314 315076
rect 288157 314938 288223 314941
rect 295742 314938 295748 314940
rect 288157 314936 295748 314938
rect 288157 314880 288162 314936
rect 288218 314880 295748 314936
rect 288157 314878 295748 314880
rect 288157 314875 288223 314878
rect 295742 314876 295748 314878
rect 295812 314876 295818 314940
rect 307569 314668 307635 314669
rect 307518 314604 307524 314668
rect 307588 314666 307635 314668
rect 323393 314666 323459 314669
rect 332409 314666 332475 314669
rect 307588 314664 307680 314666
rect 307630 314608 307680 314664
rect 307588 314606 307680 314608
rect 311850 314664 332475 314666
rect 311850 314608 323398 314664
rect 323454 314608 332414 314664
rect 332470 314608 332475 314664
rect 311850 314606 332475 314608
rect 307588 314604 307635 314606
rect 307569 314603 307635 314604
rect 232262 314468 232268 314532
rect 232332 314530 232338 314532
rect 268837 314530 268903 314533
rect 292665 314530 292731 314533
rect 232332 314528 292731 314530
rect 232332 314472 268842 314528
rect 268898 314472 292670 314528
rect 292726 314472 292731 314528
rect 232332 314470 292731 314472
rect 232332 314468 232338 314470
rect 268837 314467 268903 314470
rect 292665 314467 292731 314470
rect 299841 314530 299907 314533
rect 311850 314530 311910 314606
rect 323393 314603 323459 314606
rect 332409 314603 332475 314606
rect 299841 314528 311910 314530
rect 299841 314472 299846 314528
rect 299902 314472 311910 314528
rect 299841 314470 311910 314472
rect 314101 314530 314167 314533
rect 318742 314530 318748 314532
rect 314101 314528 318748 314530
rect 314101 314472 314106 314528
rect 314162 314472 318748 314528
rect 314101 314470 318748 314472
rect 299841 314467 299907 314470
rect 314101 314467 314167 314470
rect 318742 314468 318748 314470
rect 318812 314468 318818 314532
rect 325141 314530 325207 314533
rect 325325 314530 325391 314533
rect 390737 314530 390803 314533
rect 325141 314528 390803 314530
rect 325141 314472 325146 314528
rect 325202 314472 325330 314528
rect 325386 314472 390742 314528
rect 390798 314472 390803 314528
rect 325141 314470 390803 314472
rect 325141 314467 325207 314470
rect 325325 314467 325391 314470
rect 390737 314467 390803 314470
rect 241094 314332 241100 314396
rect 241164 314394 241170 314396
rect 277761 314394 277827 314397
rect 301221 314394 301287 314397
rect 323577 314394 323643 314397
rect 388161 314394 388227 314397
rect 241164 314392 301287 314394
rect 241164 314336 277766 314392
rect 277822 314336 301226 314392
rect 301282 314336 301287 314392
rect 241164 314334 301287 314336
rect 241164 314332 241170 314334
rect 277761 314331 277827 314334
rect 301221 314331 301287 314334
rect 311850 314392 388227 314394
rect 311850 314336 323582 314392
rect 323638 314336 388166 314392
rect 388222 314336 388227 314392
rect 311850 314334 388227 314336
rect 223982 314196 223988 314260
rect 224052 314258 224058 314260
rect 263317 314258 263383 314261
rect 224052 314256 263383 314258
rect 224052 314200 263322 314256
rect 263378 314200 263383 314256
rect 224052 314198 263383 314200
rect 224052 314196 224058 314198
rect 263317 314195 263383 314198
rect 298093 314258 298159 314261
rect 298870 314258 298876 314260
rect 298093 314256 298876 314258
rect 298093 314200 298098 314256
rect 298154 314200 298876 314256
rect 298093 314198 298876 314200
rect 298093 314195 298159 314198
rect 298870 314196 298876 314198
rect 298940 314196 298946 314260
rect 301681 314258 301747 314261
rect 311850 314258 311910 314334
rect 323577 314331 323643 314334
rect 388161 314331 388227 314334
rect 301681 314256 311910 314258
rect 301681 314200 301686 314256
rect 301742 314200 311910 314256
rect 301681 314198 311910 314200
rect 326521 314258 326587 314261
rect 387333 314258 387399 314261
rect 326521 314256 387399 314258
rect 326521 314200 326526 314256
rect 326582 314200 387338 314256
rect 387394 314200 387399 314256
rect 326521 314198 387399 314200
rect 301681 314195 301747 314198
rect 326521 314195 326587 314198
rect 387333 314195 387399 314198
rect 223246 314060 223252 314124
rect 223316 314122 223322 314124
rect 238753 314122 238819 314125
rect 223316 314120 238819 314122
rect 223316 314064 238758 314120
rect 238814 314064 238819 314120
rect 223316 314062 238819 314064
rect 223316 314060 223322 314062
rect 238753 314059 238819 314062
rect 244590 314060 244596 314124
rect 244660 314122 244666 314124
rect 305310 314122 305316 314124
rect 244660 314062 305316 314122
rect 244660 314060 244666 314062
rect 305310 314060 305316 314062
rect 305380 314060 305386 314124
rect 232814 313924 232820 313988
rect 232884 313986 232890 313988
rect 292982 313986 292988 313988
rect 232884 313926 292988 313986
rect 232884 313924 232890 313926
rect 292982 313924 292988 313926
rect 293052 313924 293058 313988
rect 296253 313986 296319 313989
rect 325325 313986 325391 313989
rect 393405 313986 393471 313989
rect 477493 313986 477559 313989
rect 296253 313984 325391 313986
rect 296253 313928 296258 313984
rect 296314 313928 325330 313984
rect 325386 313928 325391 313984
rect 296253 313926 325391 313928
rect 296253 313923 296319 313926
rect 325325 313923 325391 313926
rect 393270 313984 477559 313986
rect 393270 313928 393410 313984
rect 393466 313928 477498 313984
rect 477554 313928 477559 313984
rect 393270 313926 477559 313928
rect 239438 313788 239444 313852
rect 239508 313850 239514 313852
rect 269665 313850 269731 313853
rect 299422 313850 299428 313852
rect 239508 313848 299428 313850
rect 239508 313792 269670 313848
rect 269726 313792 299428 313848
rect 239508 313790 299428 313792
rect 239508 313788 239514 313790
rect 269665 313787 269731 313790
rect 299422 313788 299428 313790
rect 299492 313788 299498 313852
rect 319529 313850 319595 313853
rect 393270 313850 393330 313926
rect 393405 313923 393471 313926
rect 477493 313923 477559 313926
rect 319529 313848 393330 313850
rect 319529 313792 319534 313848
rect 319590 313792 393330 313848
rect 319529 313790 393330 313792
rect 319529 313787 319595 313790
rect 241278 313652 241284 313716
rect 241348 313714 241354 313716
rect 271689 313714 271755 313717
rect 241348 313712 271755 313714
rect 241348 313656 271694 313712
rect 271750 313656 271755 313712
rect 241348 313654 271755 313656
rect 241348 313652 241354 313654
rect 271689 313651 271755 313654
rect 293861 313714 293927 313717
rect 324681 313714 324747 313717
rect 327349 313714 327415 313717
rect 293861 313712 327415 313714
rect 293861 313656 293866 313712
rect 293922 313656 324686 313712
rect 324742 313656 327354 313712
rect 327410 313656 327415 313712
rect 293861 313654 327415 313656
rect 293861 313651 293927 313654
rect 324681 313651 324747 313654
rect 327349 313651 327415 313654
rect 267365 313578 267431 313581
rect 299606 313578 299612 313580
rect 267365 313576 299612 313578
rect 267365 313520 267370 313576
rect 267426 313520 299612 313576
rect 267365 313518 299612 313520
rect 267365 313515 267431 313518
rect 299606 313516 299612 313518
rect 299676 313516 299682 313580
rect 300853 313578 300919 313581
rect 301446 313578 301452 313580
rect 300853 313576 301452 313578
rect 300853 313520 300858 313576
rect 300914 313520 301452 313576
rect 300853 313518 301452 313520
rect 300853 313515 300919 313518
rect 301446 313516 301452 313518
rect 301516 313516 301522 313580
rect 271689 313442 271755 313445
rect 301221 313442 301287 313445
rect 271689 313440 301287 313442
rect 271689 313384 271694 313440
rect 271750 313384 301226 313440
rect 301282 313384 301287 313440
rect 271689 313382 301287 313384
rect 271689 313379 271755 313382
rect 301221 313379 301287 313382
rect 247902 313108 247908 313172
rect 247972 313170 247978 313172
rect 307753 313170 307819 313173
rect 247972 313168 307819 313170
rect 247972 313112 307758 313168
rect 307814 313112 307819 313168
rect 247972 313110 307819 313112
rect 247972 313108 247978 313110
rect 307753 313107 307819 313110
rect 323853 313170 323919 313173
rect 384389 313170 384455 313173
rect 323853 313168 384455 313170
rect 323853 313112 323858 313168
rect 323914 313112 384394 313168
rect 384450 313112 384455 313168
rect 323853 313110 384455 313112
rect 323853 313107 323919 313110
rect 384389 313107 384455 313110
rect 249558 312972 249564 313036
rect 249628 313034 249634 313036
rect 309358 313034 309364 313036
rect 249628 312974 309364 313034
rect 249628 312972 249634 312974
rect 309358 312972 309364 312974
rect 309428 312972 309434 313036
rect 320909 313034 320975 313037
rect 321461 313034 321527 313037
rect 381169 313034 381235 313037
rect 320909 313032 383670 313034
rect 320909 312976 320914 313032
rect 320970 312976 321466 313032
rect 321522 312976 381174 313032
rect 381230 312976 383670 313032
rect 320909 312974 383670 312976
rect 320909 312971 320975 312974
rect 321461 312971 321527 312974
rect 381169 312971 381235 312974
rect 252318 312836 252324 312900
rect 252388 312898 252394 312900
rect 311893 312898 311959 312901
rect 252388 312896 311959 312898
rect 252388 312840 311898 312896
rect 311954 312840 311959 312896
rect 252388 312838 311959 312840
rect 252388 312836 252394 312838
rect 311893 312835 311959 312838
rect 323209 312898 323275 312901
rect 324129 312898 324195 312901
rect 344093 312898 344159 312901
rect 323209 312896 344159 312898
rect 323209 312840 323214 312896
rect 323270 312840 324134 312896
rect 324190 312840 344098 312896
rect 344154 312840 344159 312896
rect 323209 312838 344159 312840
rect 323209 312835 323275 312838
rect 324129 312835 324195 312838
rect 344093 312835 344159 312838
rect 226190 312700 226196 312764
rect 226260 312762 226266 312764
rect 249793 312762 249859 312765
rect 226260 312760 249859 312762
rect 226260 312704 249798 312760
rect 249854 312704 249859 312760
rect 226260 312702 249859 312704
rect 226260 312700 226266 312702
rect 249793 312699 249859 312702
rect 251766 312700 251772 312764
rect 251836 312762 251842 312764
rect 326061 312762 326127 312765
rect 326981 312762 327047 312765
rect 333697 312762 333763 312765
rect 251836 312702 302250 312762
rect 251836 312700 251842 312702
rect 299841 312628 299907 312629
rect 234286 312564 234292 312628
rect 234356 312626 234362 312628
rect 292614 312626 292620 312628
rect 234356 312566 292620 312626
rect 234356 312564 234362 312566
rect 292614 312564 292620 312566
rect 292684 312564 292690 312628
rect 299790 312626 299796 312628
rect 299750 312566 299796 312626
rect 299860 312624 299907 312628
rect 299902 312568 299907 312624
rect 299790 312564 299796 312566
rect 299860 312564 299907 312568
rect 302190 312626 302250 312702
rect 326061 312760 333763 312762
rect 326061 312704 326066 312760
rect 326122 312704 326986 312760
rect 327042 312704 333702 312760
rect 333758 312704 333763 312760
rect 326061 312702 333763 312704
rect 326061 312699 326127 312702
rect 326981 312699 327047 312702
rect 333697 312699 333763 312702
rect 311934 312626 311940 312628
rect 302190 312566 311940 312626
rect 311934 312564 311940 312566
rect 312004 312626 312010 312628
rect 313181 312626 313247 312629
rect 312004 312624 313247 312626
rect 312004 312568 313186 312624
rect 313242 312568 313247 312624
rect 312004 312566 313247 312568
rect 312004 312564 312010 312566
rect 299841 312563 299907 312564
rect 313181 312563 313247 312566
rect 327022 312564 327028 312628
rect 327092 312626 327098 312628
rect 334249 312626 334315 312629
rect 327092 312624 334315 312626
rect 327092 312568 334254 312624
rect 334310 312568 334315 312624
rect 327092 312566 334315 312568
rect 327092 312564 327098 312566
rect 334249 312563 334315 312566
rect 222009 312490 222075 312493
rect 311382 312490 311388 312492
rect 222009 312488 311388 312490
rect 222009 312432 222014 312488
rect 222070 312432 311388 312488
rect 222009 312430 311388 312432
rect 222009 312427 222075 312430
rect 311382 312428 311388 312430
rect 311452 312428 311458 312492
rect 383610 312490 383670 312974
rect 502333 312490 502399 312493
rect 383610 312488 502399 312490
rect 383610 312432 502338 312488
rect 502394 312432 502399 312488
rect 383610 312430 502399 312432
rect 502333 312427 502399 312430
rect 234470 312292 234476 312356
rect 234540 312354 234546 312356
rect 293350 312354 293356 312356
rect 234540 312294 293356 312354
rect 234540 312292 234546 312294
rect 293350 312292 293356 312294
rect 293420 312292 293426 312356
rect 309133 312218 309199 312221
rect 310278 312218 310284 312220
rect 309133 312216 310284 312218
rect 309133 312160 309138 312216
rect 309194 312160 310284 312216
rect 309133 312158 310284 312160
rect 309133 312155 309199 312158
rect 310278 312156 310284 312158
rect 310348 312156 310354 312220
rect 579613 312082 579679 312085
rect 583520 312082 584960 312172
rect 579613 312080 584960 312082
rect 579613 312024 579618 312080
rect 579674 312024 584960 312080
rect 579613 312022 584960 312024
rect 579613 312019 579679 312022
rect 282862 311884 282868 311948
rect 282932 311946 282938 311948
rect 283230 311946 283236 311948
rect 282932 311886 283236 311946
rect 282932 311884 282938 311886
rect 283230 311884 283236 311886
rect 283300 311884 283306 311948
rect 583520 311932 584960 312022
rect 316585 311810 316651 311813
rect 317229 311810 317295 311813
rect 381445 311810 381511 311813
rect 316585 311808 381511 311810
rect 316585 311752 316590 311808
rect 316646 311752 317234 311808
rect 317290 311752 381450 311808
rect 381506 311752 381511 311808
rect 316585 311750 381511 311752
rect 316585 311747 316651 311750
rect 317229 311747 317295 311750
rect 381445 311747 381511 311750
rect 232630 311612 232636 311676
rect 232700 311674 232706 311676
rect 291142 311674 291148 311676
rect 232700 311614 291148 311674
rect 232700 311612 232706 311614
rect 291142 311612 291148 311614
rect 291212 311612 291218 311676
rect 318374 311612 318380 311676
rect 318444 311674 318450 311676
rect 318742 311674 318748 311676
rect 318444 311614 318748 311674
rect 318444 311612 318450 311614
rect 318742 311612 318748 311614
rect 318812 311674 318818 311676
rect 330845 311674 330911 311677
rect 318812 311672 330911 311674
rect 318812 311616 330850 311672
rect 330906 311616 330911 311672
rect 318812 311614 330911 311616
rect 318812 311612 318818 311614
rect 330845 311611 330911 311614
rect 230054 311476 230060 311540
rect 230124 311538 230130 311540
rect 289997 311538 290063 311541
rect 379145 311538 379211 311541
rect 230124 311536 290063 311538
rect 230124 311480 290002 311536
rect 290058 311480 290063 311536
rect 230124 311478 290063 311480
rect 230124 311476 230130 311478
rect 289997 311475 290063 311478
rect 322430 311536 379211 311538
rect 322430 311480 379150 311536
rect 379206 311480 379211 311536
rect 322430 311478 379211 311480
rect 231342 311340 231348 311404
rect 231412 311402 231418 311404
rect 291878 311402 291884 311404
rect 231412 311342 291884 311402
rect 231412 311340 231418 311342
rect 291878 311340 291884 311342
rect 291948 311340 291954 311404
rect 231158 311204 231164 311268
rect 231228 311266 231234 311268
rect 292246 311266 292252 311268
rect 231228 311206 292252 311266
rect 231228 311204 231234 311206
rect 292246 311204 292252 311206
rect 292316 311204 292322 311268
rect 317873 311266 317939 311269
rect 318517 311266 318583 311269
rect 322430 311266 322490 311478
rect 379145 311475 379211 311478
rect 329005 311402 329071 311405
rect 380934 311402 380940 311404
rect 329005 311400 380940 311402
rect 329005 311344 329010 311400
rect 329066 311344 380940 311400
rect 329005 311342 380940 311344
rect 329005 311339 329071 311342
rect 380934 311340 380940 311342
rect 381004 311340 381010 311404
rect 317873 311264 322490 311266
rect 317873 311208 317878 311264
rect 317934 311208 318522 311264
rect 318578 311208 322490 311264
rect 317873 311206 322490 311208
rect 324405 311266 324471 311269
rect 324957 311266 325023 311269
rect 324405 311264 374010 311266
rect 324405 311208 324410 311264
rect 324466 311208 324962 311264
rect 325018 311208 374010 311264
rect 324405 311206 374010 311208
rect 317873 311203 317939 311206
rect 318517 311203 318583 311206
rect 324405 311203 324471 311206
rect 324957 311203 325023 311206
rect 229318 311068 229324 311132
rect 229388 311130 229394 311132
rect 290774 311130 290780 311132
rect 229388 311070 290780 311130
rect 229388 311068 229394 311070
rect 290774 311068 290780 311070
rect 290844 311068 290850 311132
rect 322013 311130 322079 311133
rect 322197 311130 322263 311133
rect 329005 311130 329071 311133
rect 322013 311128 329071 311130
rect 322013 311072 322018 311128
rect 322074 311072 322202 311128
rect 322258 311072 329010 311128
rect 329066 311072 329071 311128
rect 322013 311070 329071 311072
rect 373950 311130 374010 311206
rect 387977 311130 388043 311133
rect 552657 311130 552723 311133
rect 373950 311128 552723 311130
rect 373950 311072 387982 311128
rect 388038 311072 552662 311128
rect 552718 311072 552723 311128
rect 373950 311070 552723 311072
rect 322013 311067 322079 311070
rect 322197 311067 322263 311070
rect 329005 311067 329071 311070
rect 387977 311067 388043 311070
rect 552657 311067 552723 311070
rect 287646 310932 287652 310996
rect 287716 310994 287722 310996
rect 322105 310994 322171 310997
rect 287716 310992 322171 310994
rect 287716 310936 322110 310992
rect 322166 310936 322171 310992
rect 287716 310934 322171 310936
rect 287716 310932 287722 310934
rect 322105 310931 322171 310934
rect 289169 310858 289235 310861
rect 318742 310858 318748 310860
rect 289169 310856 318748 310858
rect 289169 310800 289174 310856
rect 289230 310800 318748 310856
rect 289169 310798 318748 310800
rect 289169 310795 289235 310798
rect 318742 310796 318748 310798
rect 318812 310796 318818 310860
rect 261937 310450 262003 310453
rect 288433 310450 288499 310453
rect 258030 310448 288499 310450
rect 258030 310392 261942 310448
rect 261998 310392 288438 310448
rect 288494 310392 288499 310448
rect 258030 310390 288499 310392
rect 228950 310252 228956 310316
rect 229020 310314 229026 310316
rect 258030 310314 258090 310390
rect 261937 310387 262003 310390
rect 288433 310387 288499 310390
rect 291101 310450 291167 310453
rect 298686 310450 298692 310452
rect 291101 310448 298692 310450
rect 291101 310392 291106 310448
rect 291162 310392 298692 310448
rect 291101 310390 298692 310392
rect 291101 310387 291167 310390
rect 298686 310388 298692 310390
rect 298756 310388 298762 310452
rect 330385 310450 330451 310453
rect 393313 310450 393379 310453
rect 330385 310448 393379 310450
rect 330385 310392 330390 310448
rect 330446 310392 393318 310448
rect 393374 310392 393379 310448
rect 330385 310390 393379 310392
rect 330385 310387 330451 310390
rect 393313 310387 393379 310390
rect 286041 310314 286107 310317
rect 229020 310254 258090 310314
rect 267690 310312 286107 310314
rect 267690 310256 286046 310312
rect 286102 310256 286107 310312
rect 267690 310254 286107 310256
rect 229020 310252 229026 310254
rect 227478 310116 227484 310180
rect 227548 310178 227554 310180
rect 264881 310178 264947 310181
rect 267690 310178 267750 310254
rect 286041 310251 286107 310254
rect 323301 310314 323367 310317
rect 324221 310314 324287 310317
rect 392117 310314 392183 310317
rect 323301 310312 392183 310314
rect 323301 310256 323306 310312
rect 323362 310256 324226 310312
rect 324282 310256 392122 310312
rect 392178 310256 392183 310312
rect 323301 310254 392183 310256
rect 323301 310251 323367 310254
rect 324221 310251 324287 310254
rect 392117 310251 392183 310254
rect 227548 310176 267750 310178
rect 227548 310120 264886 310176
rect 264942 310120 267750 310176
rect 227548 310118 267750 310120
rect 321921 310178 321987 310181
rect 322565 310178 322631 310181
rect 330385 310178 330451 310181
rect 387885 310178 387951 310181
rect 321921 310176 330451 310178
rect 321921 310120 321926 310176
rect 321982 310120 322570 310176
rect 322626 310120 330390 310176
rect 330446 310120 330451 310176
rect 321921 310118 330451 310120
rect 227548 310116 227554 310118
rect 264881 310115 264947 310118
rect 321921 310115 321987 310118
rect 322565 310115 322631 310118
rect 330385 310115 330451 310118
rect 330526 310176 387951 310178
rect 330526 310120 387890 310176
rect 387946 310120 387951 310176
rect 330526 310118 387951 310120
rect 228214 309980 228220 310044
rect 228284 310042 228290 310044
rect 288198 310042 288204 310044
rect 228284 309982 288204 310042
rect 228284 309980 228290 309982
rect 288198 309980 288204 309982
rect 288268 309980 288274 310044
rect 322933 310042 322999 310045
rect 330526 310042 330586 310118
rect 387885 310115 387951 310118
rect 322933 310040 330586 310042
rect 322933 309984 322938 310040
rect 322994 309984 330586 310040
rect 322933 309982 330586 309984
rect 330753 310042 330819 310045
rect 390553 310042 390619 310045
rect 330753 310040 390619 310042
rect 330753 309984 330758 310040
rect 330814 309984 390558 310040
rect 390614 309984 390619 310040
rect 330753 309982 390619 309984
rect 322933 309979 322999 309982
rect 330753 309979 330819 309982
rect 390553 309979 390619 309982
rect 244774 309844 244780 309908
rect 244844 309906 244850 309908
rect 304993 309906 305059 309909
rect 244844 309904 305059 309906
rect 244844 309848 304998 309904
rect 305054 309848 305059 309904
rect 244844 309846 305059 309848
rect 244844 309844 244850 309846
rect 304993 309843 305059 309846
rect 308254 309844 308260 309908
rect 308324 309906 308330 309908
rect 315614 309906 315620 309908
rect 308324 309846 315620 309906
rect 308324 309844 308330 309846
rect 315614 309844 315620 309846
rect 315684 309906 315690 309908
rect 375966 309906 375972 309908
rect 315684 309846 375972 309906
rect 315684 309844 315690 309846
rect 375966 309844 375972 309846
rect 376036 309844 376042 309908
rect 225454 309708 225460 309772
rect 225524 309770 225530 309772
rect 286358 309770 286364 309772
rect 225524 309710 286364 309770
rect 225524 309708 225530 309710
rect 286358 309708 286364 309710
rect 286428 309708 286434 309772
rect 286501 309770 286567 309773
rect 322933 309770 322999 309773
rect 286501 309768 322999 309770
rect 286501 309712 286506 309768
rect 286562 309712 322938 309768
rect 322994 309712 322999 309768
rect 286501 309710 322999 309712
rect 286501 309707 286567 309710
rect 322933 309707 322999 309710
rect 326705 309770 326771 309773
rect 330753 309770 330819 309773
rect 326705 309768 330819 309770
rect 326705 309712 326710 309768
rect 326766 309712 330758 309768
rect 330814 309712 330819 309768
rect 326705 309710 330819 309712
rect 326705 309707 326771 309710
rect 330753 309707 330819 309710
rect 271597 309634 271663 309637
rect 328453 309634 328519 309637
rect 271597 309632 328519 309634
rect 271597 309576 271602 309632
rect 271658 309576 328458 309632
rect 328514 309576 328519 309632
rect 271597 309574 328519 309576
rect 271597 309571 271663 309574
rect 328453 309571 328519 309574
rect 318977 309090 319043 309093
rect 319897 309090 319963 309093
rect 318977 309088 319963 309090
rect 318977 309032 318982 309088
rect 319038 309032 319902 309088
rect 319958 309032 319963 309088
rect 318977 309030 319963 309032
rect 318977 309027 319043 309030
rect 319897 309027 319963 309030
rect 321829 309090 321895 309093
rect 322289 309090 322355 309093
rect 323025 309090 323091 309093
rect 324037 309090 324103 309093
rect 392025 309090 392091 309093
rect 321829 309088 322858 309090
rect 321829 309032 321834 309088
rect 321890 309032 322294 309088
rect 322350 309032 322858 309088
rect 321829 309030 322858 309032
rect 321829 309027 321895 309030
rect 322289 309027 322355 309030
rect 322798 308954 322858 309030
rect 323025 309088 392091 309090
rect 323025 309032 323030 309088
rect 323086 309032 324042 309088
rect 324098 309032 392030 309088
rect 392086 309032 392091 309088
rect 323025 309030 392091 309032
rect 323025 309027 323091 309030
rect 324037 309027 324103 309030
rect 392025 309027 392091 309030
rect 381077 308954 381143 308957
rect 322798 308952 381143 308954
rect 322798 308896 381082 308952
rect 381138 308896 381143 308952
rect 322798 308894 381143 308896
rect 381077 308891 381143 308894
rect 269665 308818 269731 308821
rect 312670 308818 312676 308820
rect 269665 308816 312676 308818
rect 269665 308760 269670 308816
rect 269726 308760 312676 308816
rect 269665 308758 312676 308760
rect 269665 308755 269731 308758
rect 312670 308756 312676 308758
rect 312740 308818 312746 308820
rect 370681 308818 370747 308821
rect 312740 308816 370747 308818
rect 312740 308760 370686 308816
rect 370742 308760 370747 308816
rect 312740 308758 370747 308760
rect 312740 308756 312746 308758
rect 370681 308755 370747 308758
rect 298829 308682 298895 308685
rect 303470 308682 303476 308684
rect 298829 308680 303476 308682
rect 298829 308624 298834 308680
rect 298890 308624 303476 308680
rect 298829 308622 303476 308624
rect 298829 308619 298895 308622
rect 303470 308620 303476 308622
rect 303540 308682 303546 308684
rect 355174 308682 355180 308684
rect 303540 308622 355180 308682
rect 303540 308620 303546 308622
rect 355174 308620 355180 308622
rect 355244 308620 355250 308684
rect 238518 308484 238524 308548
rect 238588 308546 238594 308548
rect 298093 308546 298159 308549
rect 238588 308544 298159 308546
rect 238588 308488 298098 308544
rect 298154 308488 298159 308544
rect 238588 308486 298159 308488
rect 238588 308484 238594 308486
rect 298093 308483 298159 308486
rect 319897 308546 319963 308549
rect 342846 308546 342852 308548
rect 319897 308544 342852 308546
rect 319897 308488 319902 308544
rect 319958 308488 342852 308544
rect 319897 308486 342852 308488
rect 319897 308483 319963 308486
rect 342846 308484 342852 308486
rect 342916 308484 342922 308548
rect 234102 308348 234108 308412
rect 234172 308410 234178 308412
rect 294822 308410 294828 308412
rect 234172 308350 294828 308410
rect 234172 308348 234178 308350
rect 294822 308348 294828 308350
rect 294892 308348 294898 308412
rect 299974 308348 299980 308412
rect 300044 308410 300050 308412
rect 309777 308410 309843 308413
rect 300044 308408 309843 308410
rect 300044 308352 309782 308408
rect 309838 308352 309843 308408
rect 300044 308350 309843 308352
rect 300044 308348 300050 308350
rect 309777 308347 309843 308350
rect 236862 307668 236868 307732
rect 236932 307730 236938 307732
rect 296478 307730 296484 307732
rect 236932 307670 296484 307730
rect 236932 307668 236938 307670
rect 296478 307668 296484 307670
rect 296548 307668 296554 307732
rect 321093 307730 321159 307733
rect 380433 307730 380499 307733
rect 321093 307728 380499 307730
rect 321093 307672 321098 307728
rect 321154 307672 380438 307728
rect 380494 307672 380499 307728
rect 321093 307670 380499 307672
rect 321093 307667 321159 307670
rect 380433 307667 380499 307670
rect 204897 307594 204963 307597
rect 266169 307594 266235 307597
rect 283046 307594 283052 307596
rect 204897 307592 283052 307594
rect 204897 307536 204902 307592
rect 204958 307536 266174 307592
rect 266230 307536 283052 307592
rect 204897 307534 283052 307536
rect 204897 307531 204963 307534
rect 266169 307531 266235 307534
rect 283046 307532 283052 307534
rect 283116 307532 283122 307596
rect 325969 307594 326035 307597
rect 326429 307594 326495 307597
rect 384982 307594 384988 307596
rect 325969 307592 384988 307594
rect 325969 307536 325974 307592
rect 326030 307536 326434 307592
rect 326490 307536 384988 307592
rect 325969 307534 384988 307536
rect 325969 307531 326035 307534
rect 326429 307531 326495 307534
rect 384982 307532 384988 307534
rect 385052 307532 385058 307596
rect 212073 307458 212139 307461
rect 289118 307458 289124 307460
rect 212073 307456 289124 307458
rect 212073 307400 212078 307456
rect 212134 307400 289124 307456
rect 212073 307398 289124 307400
rect 212073 307395 212139 307398
rect 289118 307396 289124 307398
rect 289188 307396 289194 307460
rect 357934 307458 357940 307460
rect 306330 307398 357940 307458
rect 216121 307322 216187 307325
rect 297582 307322 297588 307324
rect 216121 307320 297588 307322
rect 216121 307264 216126 307320
rect 216182 307264 297588 307320
rect 216121 307262 297588 307264
rect 216121 307259 216187 307262
rect 297582 307260 297588 307262
rect 297652 307260 297658 307324
rect 218973 307186 219039 307189
rect 302693 307186 302759 307189
rect 306330 307186 306390 307398
rect 357934 307396 357940 307398
rect 358004 307396 358010 307460
rect 308949 307322 309015 307325
rect 356646 307322 356652 307324
rect 308949 307320 356652 307322
rect 308949 307264 308954 307320
rect 309010 307264 356652 307320
rect 308949 307262 356652 307264
rect 308949 307259 309015 307262
rect 356646 307260 356652 307262
rect 356716 307260 356722 307324
rect 218973 307184 306390 307186
rect 218973 307128 218978 307184
rect 219034 307128 302698 307184
rect 302754 307128 306390 307184
rect 218973 307126 306390 307128
rect 218973 307123 219039 307126
rect 302693 307123 302759 307126
rect 210141 307050 210207 307053
rect 301262 307050 301268 307052
rect 210141 307048 301268 307050
rect 210141 306992 210146 307048
rect 210202 306992 301268 307048
rect 210141 306990 301268 306992
rect 210141 306987 210207 306990
rect 301262 306988 301268 306990
rect 301332 306988 301338 307052
rect 222694 306852 222700 306916
rect 222764 306914 222770 306916
rect 260741 306914 260807 306917
rect 222764 306912 260807 306914
rect 222764 306856 260746 306912
rect 260802 306856 260807 306912
rect 222764 306854 260807 306856
rect 222764 306852 222770 306854
rect 260741 306851 260807 306854
rect 282085 306914 282151 306917
rect 329046 306914 329052 306916
rect 282085 306912 329052 306914
rect 282085 306856 282090 306912
rect 282146 306856 329052 306912
rect 282085 306854 329052 306856
rect 282085 306851 282151 306854
rect 329046 306852 329052 306854
rect 329116 306852 329122 306916
rect 238569 306506 238635 306509
rect 238702 306506 238708 306508
rect 238569 306504 238708 306506
rect 238569 306448 238574 306504
rect 238630 306448 238708 306504
rect 238569 306446 238708 306448
rect 238569 306443 238635 306446
rect 238702 306444 238708 306446
rect 238772 306444 238778 306508
rect 317689 306370 317755 306373
rect 389173 306370 389239 306373
rect 317689 306368 389239 306370
rect -960 306234 480 306324
rect 317689 306312 317694 306368
rect 317750 306312 389178 306368
rect 389234 306312 389239 306368
rect 317689 306310 389239 306312
rect 317689 306307 317755 306310
rect 389173 306307 389239 306310
rect 4061 306234 4127 306237
rect 238661 306236 238727 306237
rect 238661 306234 238708 306236
rect -960 306232 4127 306234
rect -960 306176 4066 306232
rect 4122 306176 4127 306232
rect -960 306174 4127 306176
rect 238616 306232 238708 306234
rect 238772 306234 238778 306236
rect 321737 306234 321803 306237
rect 389265 306234 389331 306237
rect 238616 306176 238666 306232
rect 238616 306174 238708 306176
rect -960 306084 480 306174
rect 4061 306171 4127 306174
rect 238661 306172 238708 306174
rect 238772 306174 238854 306234
rect 321737 306232 389331 306234
rect 321737 306176 321742 306232
rect 321798 306176 389270 306232
rect 389326 306176 389331 306232
rect 321737 306174 389331 306176
rect 238772 306172 238778 306174
rect 238661 306171 238727 306172
rect 321737 306171 321803 306174
rect 389265 306171 389331 306174
rect 325877 306098 325943 306101
rect 326797 306098 326863 306101
rect 391933 306098 391999 306101
rect 325877 306096 391999 306098
rect 325877 306040 325882 306096
rect 325938 306040 326802 306096
rect 326858 306040 391938 306096
rect 391994 306040 391999 306096
rect 325877 306038 391999 306040
rect 325877 306035 325943 306038
rect 326797 306035 326863 306038
rect 391933 306035 391999 306038
rect 319713 305962 319779 305965
rect 377254 305962 377260 305964
rect 319713 305960 377260 305962
rect 319713 305904 319718 305960
rect 319774 305904 377260 305960
rect 319713 305902 377260 305904
rect 319713 305899 319779 305902
rect 377254 305900 377260 305902
rect 377324 305900 377330 305964
rect 316534 305826 316540 305828
rect 315990 305766 316540 305826
rect 306005 305690 306071 305693
rect 315990 305690 316050 305766
rect 316534 305764 316540 305766
rect 316604 305826 316610 305828
rect 355317 305826 355383 305829
rect 316604 305824 355383 305826
rect 316604 305768 355322 305824
rect 355378 305768 355383 305824
rect 316604 305766 355383 305768
rect 316604 305764 316610 305766
rect 355317 305763 355383 305766
rect 306005 305688 316050 305690
rect 306005 305632 306010 305688
rect 306066 305632 316050 305688
rect 306005 305630 316050 305632
rect 306005 305627 306071 305630
rect 317689 305010 317755 305013
rect 318333 305010 318399 305013
rect 317689 305008 318399 305010
rect 317689 304952 317694 305008
rect 317750 304952 318338 305008
rect 318394 304952 318399 305008
rect 317689 304950 318399 304952
rect 317689 304947 317755 304950
rect 318333 304947 318399 304950
rect 321737 305010 321803 305013
rect 322841 305010 322907 305013
rect 321737 305008 322907 305010
rect 321737 304952 321742 305008
rect 321798 304952 322846 305008
rect 322902 304952 322907 305008
rect 321737 304950 322907 304952
rect 321737 304947 321803 304950
rect 322841 304947 322907 304950
rect 327574 304948 327580 305012
rect 327644 305010 327650 305012
rect 570597 305010 570663 305013
rect 327644 305008 570663 305010
rect 327644 304952 570602 305008
rect 570658 304952 570663 305008
rect 327644 304950 570663 304952
rect 327644 304948 327650 304950
rect 570597 304947 570663 304950
rect 269021 304874 269087 304877
rect 282862 304874 282868 304876
rect 269021 304872 282868 304874
rect 269021 304816 269026 304872
rect 269082 304816 282868 304872
rect 269021 304814 282868 304816
rect 269021 304811 269087 304814
rect 282862 304812 282868 304814
rect 282932 304812 282938 304876
rect 320766 304812 320772 304876
rect 320836 304874 320842 304876
rect 379462 304874 379468 304876
rect 320836 304814 379468 304874
rect 320836 304812 320842 304814
rect 379462 304812 379468 304814
rect 379532 304812 379538 304876
rect 209313 304738 209379 304741
rect 304574 304738 304580 304740
rect 209313 304736 304580 304738
rect 209313 304680 209318 304736
rect 209374 304680 304580 304736
rect 209313 304678 304580 304680
rect 209313 304675 209379 304678
rect 304574 304676 304580 304678
rect 304644 304738 304650 304740
rect 362902 304738 362908 304740
rect 304644 304678 362908 304738
rect 304644 304676 304650 304678
rect 362902 304676 362908 304678
rect 362972 304676 362978 304740
rect 296345 304602 296411 304605
rect 312077 304602 312143 304605
rect 367686 304602 367692 304604
rect 296345 304600 367692 304602
rect 296345 304544 296350 304600
rect 296406 304544 312082 304600
rect 312138 304544 367692 304600
rect 296345 304542 367692 304544
rect 296345 304539 296411 304542
rect 312077 304539 312143 304542
rect 367686 304540 367692 304542
rect 367756 304540 367762 304604
rect 235574 304404 235580 304468
rect 235644 304466 235650 304468
rect 295333 304466 295399 304469
rect 235644 304464 295399 304466
rect 235644 304408 295338 304464
rect 295394 304408 295399 304464
rect 235644 304406 295399 304408
rect 235644 304404 235650 304406
rect 295333 304403 295399 304406
rect 310697 304466 310763 304469
rect 320725 304466 320791 304469
rect 363454 304466 363460 304468
rect 310697 304464 320791 304466
rect 310697 304408 310702 304464
rect 310758 304408 320730 304464
rect 320786 304408 320791 304464
rect 310697 304406 320791 304408
rect 310697 304403 310763 304406
rect 320725 304403 320791 304406
rect 320958 304406 363460 304466
rect 206461 304330 206527 304333
rect 269021 304330 269087 304333
rect 206461 304328 269087 304330
rect 206461 304272 206466 304328
rect 206522 304272 269026 304328
rect 269082 304272 269087 304328
rect 206461 304270 269087 304272
rect 206461 304267 206527 304270
rect 269021 304267 269087 304270
rect 310881 304330 310947 304333
rect 320958 304330 321018 304406
rect 363454 304404 363460 304406
rect 363524 304404 363530 304468
rect 310881 304328 321018 304330
rect 310881 304272 310886 304328
rect 310942 304272 321018 304328
rect 310881 304270 321018 304272
rect 321277 304330 321343 304333
rect 357566 304330 357572 304332
rect 321277 304328 357572 304330
rect 321277 304272 321282 304328
rect 321338 304272 357572 304328
rect 321277 304270 357572 304272
rect 310881 304267 310947 304270
rect 321277 304267 321343 304270
rect 357566 304268 357572 304270
rect 357636 304268 357642 304332
rect 297817 304194 297883 304197
rect 314377 304194 314443 304197
rect 350758 304194 350764 304196
rect 297817 304192 350764 304194
rect 297817 304136 297822 304192
rect 297878 304136 314382 304192
rect 314438 304136 350764 304192
rect 297817 304134 350764 304136
rect 297817 304131 297883 304134
rect 314377 304131 314443 304134
rect 350758 304132 350764 304134
rect 350828 304132 350834 304196
rect 310697 303786 310763 303789
rect 311249 303786 311315 303789
rect 310697 303784 311315 303786
rect 310697 303728 310702 303784
rect 310758 303728 311254 303784
rect 311310 303728 311315 303784
rect 310697 303726 311315 303728
rect 310697 303723 310763 303726
rect 311249 303723 311315 303726
rect 310881 303650 310947 303653
rect 311433 303650 311499 303653
rect 310881 303648 311499 303650
rect 310881 303592 310886 303648
rect 310942 303592 311438 303648
rect 311494 303592 311499 303648
rect 310881 303590 311499 303592
rect 310881 303587 310947 303590
rect 311433 303587 311499 303590
rect 314837 303650 314903 303653
rect 314837 303648 314946 303650
rect 314837 303592 314842 303648
rect 314898 303592 314946 303648
rect 314837 303587 314946 303592
rect 301129 303516 301195 303517
rect 301078 303514 301084 303516
rect 301038 303454 301084 303514
rect 301148 303512 301195 303516
rect 301190 303456 301195 303512
rect 301078 303452 301084 303454
rect 301148 303452 301195 303456
rect 302918 303452 302924 303516
rect 302988 303514 302994 303516
rect 303429 303514 303495 303517
rect 302988 303512 303495 303514
rect 302988 303456 303434 303512
rect 303490 303456 303495 303512
rect 302988 303454 303495 303456
rect 302988 303452 302994 303454
rect 301129 303451 301195 303452
rect 303429 303451 303495 303454
rect 313273 303378 313339 303381
rect 314886 303378 314946 303587
rect 326889 303514 326955 303517
rect 394877 303514 394943 303517
rect 395981 303514 396047 303517
rect 326889 303512 396047 303514
rect 326889 303456 326894 303512
rect 326950 303456 394882 303512
rect 394938 303456 395986 303512
rect 396042 303456 396047 303512
rect 326889 303454 396047 303456
rect 326889 303451 326955 303454
rect 394877 303451 394943 303454
rect 395981 303451 396047 303454
rect 373206 303378 373212 303380
rect 313273 303376 373212 303378
rect 313273 303320 313278 303376
rect 313334 303320 373212 303376
rect 313273 303318 373212 303320
rect 313273 303315 313339 303318
rect 373206 303316 373212 303318
rect 373276 303316 373282 303380
rect 303521 303242 303587 303245
rect 360694 303242 360700 303244
rect 303521 303240 360700 303242
rect 303521 303184 303526 303240
rect 303582 303184 360700 303240
rect 303521 303182 360700 303184
rect 303521 303179 303587 303182
rect 360694 303180 360700 303182
rect 360764 303180 360770 303244
rect 285305 302970 285371 302973
rect 301129 302970 301195 302973
rect 285305 302968 301195 302970
rect 285305 302912 285310 302968
rect 285366 302912 301134 302968
rect 301190 302912 301195 302968
rect 285305 302910 301195 302912
rect 285305 302907 285371 302910
rect 301129 302907 301195 302910
rect 267549 302834 267615 302837
rect 325785 302834 325851 302837
rect 326889 302834 326955 302837
rect 267549 302832 326955 302834
rect 267549 302776 267554 302832
rect 267610 302776 325790 302832
rect 325846 302776 326894 302832
rect 326950 302776 326955 302832
rect 267549 302774 326955 302776
rect 267549 302771 267615 302774
rect 325785 302771 325851 302774
rect 326889 302771 326955 302774
rect 239254 302228 239260 302292
rect 239324 302290 239330 302292
rect 300577 302290 300643 302293
rect 239324 302288 300643 302290
rect 239324 302232 300582 302288
rect 300638 302232 300643 302288
rect 239324 302230 300643 302232
rect 239324 302228 239330 302230
rect 300577 302227 300643 302230
rect 302550 302228 302556 302292
rect 302620 302290 302626 302292
rect 302918 302290 302924 302292
rect 302620 302230 302924 302290
rect 302620 302228 302626 302230
rect 302918 302228 302924 302230
rect 302988 302228 302994 302292
rect 299013 302154 299079 302157
rect 358854 302154 358860 302156
rect 296670 302152 358860 302154
rect 296670 302096 299018 302152
rect 299074 302096 358860 302152
rect 296670 302094 358860 302096
rect 285213 302018 285279 302021
rect 296670 302018 296730 302094
rect 299013 302091 299079 302094
rect 358854 302092 358860 302094
rect 358924 302092 358930 302156
rect 285213 302016 296730 302018
rect 285213 301960 285218 302016
rect 285274 301960 296730 302016
rect 285213 301958 296730 301960
rect 285213 301955 285279 301958
rect 304942 301956 304948 302020
rect 305012 302018 305018 302020
rect 305494 302018 305500 302020
rect 305012 301958 305500 302018
rect 305012 301956 305018 301958
rect 305494 301956 305500 301958
rect 305564 302018 305570 302020
rect 307753 302018 307819 302021
rect 305564 302016 307819 302018
rect 305564 301960 307758 302016
rect 307814 301960 307819 302016
rect 305564 301958 307819 301960
rect 305564 301956 305570 301958
rect 307753 301955 307819 301958
rect 325141 302018 325207 302021
rect 325417 302018 325483 302021
rect 383694 302018 383700 302020
rect 325141 302016 383700 302018
rect 325141 301960 325146 302016
rect 325202 301960 325422 302016
rect 325478 301960 383700 302016
rect 325141 301958 383700 301960
rect 325141 301955 325207 301958
rect 325417 301955 325483 301958
rect 383694 301956 383700 301958
rect 383764 301956 383770 302020
rect 291377 301882 291443 301885
rect 292113 301882 292179 301885
rect 350574 301882 350580 301884
rect 291377 301880 350580 301882
rect 291377 301824 291382 301880
rect 291438 301824 292118 301880
rect 292174 301824 350580 301880
rect 291377 301822 350580 301824
rect 291377 301819 291443 301822
rect 292113 301819 292179 301822
rect 350574 301820 350580 301822
rect 350644 301820 350650 301884
rect 240910 301684 240916 301748
rect 240980 301746 240986 301748
rect 300669 301746 300735 301749
rect 240980 301744 300735 301746
rect 240980 301688 300674 301744
rect 300730 301688 300735 301744
rect 240980 301686 300735 301688
rect 240980 301684 240986 301686
rect 300669 301683 300735 301686
rect 223798 301548 223804 301612
rect 223868 301610 223874 301612
rect 227161 301610 227227 301613
rect 223868 301608 227227 301610
rect 223868 301552 227166 301608
rect 227222 301552 227227 301608
rect 223868 301550 227227 301552
rect 223868 301548 223874 301550
rect 227161 301547 227227 301550
rect 246430 301548 246436 301612
rect 246500 301610 246506 301612
rect 304942 301610 304948 301612
rect 246500 301550 304948 301610
rect 246500 301548 246506 301550
rect 304942 301548 304948 301550
rect 305012 301548 305018 301612
rect 235390 301412 235396 301476
rect 235460 301474 235466 301476
rect 295333 301474 295399 301477
rect 235460 301472 295399 301474
rect 235460 301416 295338 301472
rect 295394 301416 295399 301472
rect 235460 301414 295399 301416
rect 235460 301412 235466 301414
rect 295333 301411 295399 301414
rect 305821 301474 305887 301477
rect 321502 301474 321508 301476
rect 305821 301472 321508 301474
rect 305821 301416 305826 301472
rect 305882 301416 321508 301472
rect 305821 301414 321508 301416
rect 305821 301411 305887 301414
rect 321502 301412 321508 301414
rect 321572 301474 321578 301476
rect 321645 301474 321711 301477
rect 321572 301472 321711 301474
rect 321572 301416 321650 301472
rect 321706 301416 321711 301472
rect 321572 301414 321711 301416
rect 321572 301412 321578 301414
rect 321645 301411 321711 301414
rect 274582 301276 274588 301340
rect 274652 301338 274658 301340
rect 275829 301338 275895 301341
rect 274652 301336 275895 301338
rect 274652 301280 275834 301336
rect 275890 301280 275895 301336
rect 274652 301278 275895 301280
rect 274652 301276 274658 301278
rect 275829 301275 275895 301278
rect 318241 300794 318307 300797
rect 384757 300794 384823 300797
rect 318241 300792 384823 300794
rect 318241 300736 318246 300792
rect 318302 300736 384762 300792
rect 384818 300736 384823 300792
rect 318241 300734 384823 300736
rect 318241 300731 318307 300734
rect 384757 300731 384823 300734
rect 323485 300658 323551 300661
rect 381486 300658 381492 300660
rect 323485 300656 381492 300658
rect 323485 300600 323490 300656
rect 323546 300600 381492 300656
rect 323485 300598 381492 300600
rect 323485 300595 323551 300598
rect 381486 300596 381492 300598
rect 381556 300596 381562 300660
rect 292389 300250 292455 300253
rect 302233 300252 302299 300253
rect 302182 300250 302188 300252
rect 292389 300248 302188 300250
rect 302252 300248 302299 300252
rect 292389 300192 292394 300248
rect 292450 300192 302188 300248
rect 302294 300192 302299 300248
rect 292389 300190 302188 300192
rect 292389 300187 292455 300190
rect 302182 300188 302188 300190
rect 302252 300188 302299 300192
rect 302233 300187 302299 300188
rect 238334 300052 238340 300116
rect 238404 300114 238410 300116
rect 298134 300114 298140 300116
rect 238404 300054 298140 300114
rect 238404 300052 238410 300054
rect 298134 300052 298140 300054
rect 298204 300052 298210 300116
rect 295149 299434 295215 299437
rect 368422 299434 368428 299436
rect 295149 299432 368428 299434
rect 295149 299376 295154 299432
rect 295210 299376 368428 299432
rect 295149 299374 368428 299376
rect 295149 299371 295215 299374
rect 368422 299372 368428 299374
rect 368492 299372 368498 299436
rect 310462 299236 310468 299300
rect 310532 299298 310538 299300
rect 311525 299298 311591 299301
rect 311750 299298 311756 299300
rect 310532 299296 311756 299298
rect 310532 299240 311530 299296
rect 311586 299240 311756 299296
rect 310532 299238 311756 299240
rect 310532 299236 310538 299238
rect 311525 299235 311591 299238
rect 311750 299236 311756 299238
rect 311820 299236 311826 299300
rect 316677 299298 316743 299301
rect 317270 299298 317276 299300
rect 316677 299296 317276 299298
rect 316677 299240 316682 299296
rect 316738 299240 317276 299296
rect 316677 299238 317276 299240
rect 316677 299235 316743 299238
rect 317270 299236 317276 299238
rect 317340 299236 317346 299300
rect 317413 299298 317479 299301
rect 318057 299298 318123 299301
rect 376886 299298 376892 299300
rect 317413 299296 376892 299298
rect 317413 299240 317418 299296
rect 317474 299240 318062 299296
rect 318118 299240 376892 299296
rect 317413 299238 376892 299240
rect 317278 299162 317338 299236
rect 317413 299235 317479 299238
rect 318057 299235 318123 299238
rect 376886 299236 376892 299238
rect 376956 299236 376962 299300
rect 375414 299162 375420 299164
rect 317278 299102 375420 299162
rect 375414 299100 375420 299102
rect 375484 299100 375490 299164
rect 228582 298964 228588 299028
rect 228652 299026 228658 299028
rect 287237 299026 287303 299029
rect 288249 299026 288315 299029
rect 228652 299024 288315 299026
rect 228652 298968 287242 299024
rect 287298 298968 288254 299024
rect 288310 298968 288315 299024
rect 228652 298966 288315 298968
rect 228652 298964 228658 298966
rect 287237 298963 287303 298966
rect 288249 298963 288315 298966
rect 235022 298828 235028 298892
rect 235092 298890 235098 298892
rect 293953 298890 294019 298893
rect 235092 298888 294019 298890
rect 235092 298832 293958 298888
rect 294014 298832 294019 298888
rect 235092 298830 294019 298832
rect 235092 298828 235098 298830
rect 293953 298827 294019 298830
rect 233918 298692 233924 298756
rect 233988 298754 233994 298756
rect 295006 298754 295012 298756
rect 233988 298694 295012 298754
rect 233988 298692 233994 298694
rect 295006 298692 295012 298694
rect 295076 298692 295082 298756
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect 304390 298074 304396 298076
rect 296670 298014 304396 298074
rect 211613 297394 211679 297397
rect 296670 297394 296730 298014
rect 304390 298012 304396 298014
rect 304460 298074 304466 298076
rect 364374 298074 364380 298076
rect 304460 298014 364380 298074
rect 304460 298012 304466 298014
rect 364374 298012 364380 298014
rect 364444 298012 364450 298076
rect 304165 297938 304231 297941
rect 359406 297938 359412 297940
rect 304165 297936 359412 297938
rect 304165 297880 304170 297936
rect 304226 297880 359412 297936
rect 304165 297878 359412 297880
rect 304165 297875 304231 297878
rect 359406 297876 359412 297878
rect 359476 297876 359482 297940
rect 302734 297604 302740 297668
rect 302804 297666 302810 297668
rect 303521 297666 303587 297669
rect 302804 297664 303587 297666
rect 302804 297608 303526 297664
rect 303582 297608 303587 297664
rect 302804 297606 303587 297608
rect 302804 297604 302810 297606
rect 303521 297603 303587 297606
rect 211613 297392 296730 297394
rect 211613 297336 211618 297392
rect 211674 297336 296730 297392
rect 211613 297334 296730 297336
rect 211613 297331 211679 297334
rect 238661 296850 238727 296853
rect 238886 296850 238892 296852
rect 238616 296848 238892 296850
rect 238616 296792 238666 296848
rect 238722 296792 238892 296848
rect 238616 296790 238892 296792
rect 238661 296787 238727 296790
rect 238886 296788 238892 296790
rect 238956 296788 238962 296852
rect 238661 296714 238727 296717
rect 238616 296712 238770 296714
rect 238616 296656 238666 296712
rect 238722 296656 238770 296712
rect 238616 296654 238770 296656
rect 238661 296651 238770 296654
rect 238710 296580 238770 296651
rect 238702 296516 238708 296580
rect 238772 296516 238778 296580
rect 226006 296380 226012 296444
rect 226076 296442 226082 296444
rect 284334 296442 284340 296444
rect 226076 296382 284340 296442
rect 226076 296380 226082 296382
rect 284334 296380 284340 296382
rect 284404 296380 284410 296444
rect 226374 296244 226380 296308
rect 226444 296306 226450 296308
rect 287973 296306 288039 296309
rect 226444 296304 288039 296306
rect 226444 296248 287978 296304
rect 288034 296248 288039 296304
rect 226444 296246 288039 296248
rect 226444 296244 226450 296246
rect 287973 296243 288039 296246
rect 223062 296108 223068 296172
rect 223132 296170 223138 296172
rect 283465 296170 283531 296173
rect 223132 296168 283531 296170
rect 223132 296112 283470 296168
rect 283526 296112 283531 296168
rect 223132 296110 283531 296112
rect 223132 296108 223138 296110
rect 283465 296107 283531 296110
rect 226558 295972 226564 296036
rect 226628 296034 226634 296036
rect 287789 296034 287855 296037
rect 226628 296032 287855 296034
rect 226628 295976 287794 296032
rect 287850 295976 287855 296032
rect 226628 295974 287855 295976
rect 226628 295972 226634 295974
rect 287789 295971 287855 295974
rect 223614 295292 223620 295356
rect 223684 295354 223690 295356
rect 225781 295354 225847 295357
rect 223684 295352 225847 295354
rect 223684 295296 225786 295352
rect 225842 295296 225847 295352
rect 223684 295294 225847 295296
rect 223684 295292 223690 295294
rect 225781 295291 225847 295294
rect 286593 295218 286659 295221
rect 286869 295218 286935 295221
rect 349102 295218 349108 295220
rect 286593 295216 349108 295218
rect 286593 295160 286598 295216
rect 286654 295160 286874 295216
rect 286930 295160 349108 295216
rect 286593 295158 349108 295160
rect 286593 295155 286659 295158
rect 286869 295155 286935 295158
rect 349102 295156 349108 295158
rect 349172 295156 349178 295220
rect 284661 295082 284727 295085
rect 345054 295082 345060 295084
rect 284661 295080 345060 295082
rect 284661 295024 284666 295080
rect 284722 295024 345060 295080
rect 284661 295022 345060 295024
rect 284661 295019 284727 295022
rect 345054 295020 345060 295022
rect 345124 295020 345130 295084
rect 229502 294884 229508 294948
rect 229572 294946 229578 294948
rect 288893 294946 288959 294949
rect 229572 294944 288959 294946
rect 229572 294888 288898 294944
rect 288954 294888 288959 294944
rect 229572 294886 288959 294888
rect 229572 294884 229578 294886
rect 288893 294883 288959 294886
rect 227294 294748 227300 294812
rect 227364 294810 227370 294812
rect 285806 294810 285812 294812
rect 227364 294750 285812 294810
rect 227364 294748 227370 294750
rect 285806 294748 285812 294750
rect 285876 294748 285882 294812
rect 225270 294612 225276 294676
rect 225340 294674 225346 294676
rect 285622 294674 285628 294676
rect 225340 294614 285628 294674
rect 225340 294612 225346 294614
rect 285622 294612 285628 294614
rect 285692 294612 285698 294676
rect 228398 294476 228404 294540
rect 228468 294538 228474 294540
rect 289629 294538 289695 294541
rect 228468 294536 289695 294538
rect 228468 294480 289634 294536
rect 289690 294480 289695 294536
rect 228468 294478 289695 294480
rect 228468 294476 228474 294478
rect 289629 294475 289695 294478
rect 232446 294340 232452 294404
rect 232516 294402 232522 294404
rect 291653 294402 291719 294405
rect 232516 294400 291719 294402
rect 232516 294344 291658 294400
rect 291714 294344 291719 294400
rect 232516 294342 291719 294344
rect 232516 294340 232522 294342
rect 291653 294339 291719 294342
rect 229870 294204 229876 294268
rect 229940 294266 229946 294268
rect 288382 294266 288388 294268
rect 229940 294206 288388 294266
rect 229940 294204 229946 294206
rect 288382 294204 288388 294206
rect 288452 294204 288458 294268
rect 284661 293994 284727 293997
rect 285121 293994 285187 293997
rect 284661 293992 285187 293994
rect 284661 293936 284666 293992
rect 284722 293936 285126 293992
rect 285182 293936 285187 293992
rect 284661 293934 285187 293936
rect 284661 293931 284727 293934
rect 285121 293931 285187 293934
rect 251950 293660 251956 293724
rect 252020 293722 252026 293724
rect 310646 293722 310652 293724
rect 252020 293662 310652 293722
rect 252020 293660 252026 293662
rect 310646 293660 310652 293662
rect 310716 293660 310722 293724
rect 242934 293524 242940 293588
rect 243004 293586 243010 293588
rect 302734 293586 302740 293588
rect 243004 293526 302740 293586
rect 243004 293524 243010 293526
rect 302734 293524 302740 293526
rect 302804 293524 302810 293588
rect 238150 293388 238156 293452
rect 238220 293450 238226 293452
rect 299289 293450 299355 293453
rect 238220 293448 299355 293450
rect 238220 293392 299294 293448
rect 299350 293392 299355 293448
rect 238220 293390 299355 293392
rect 238220 293388 238226 293390
rect 299289 293387 299355 293390
rect -960 293178 480 293268
rect 239070 293252 239076 293316
rect 239140 293314 239146 293316
rect 300577 293314 300643 293317
rect 239140 293312 300643 293314
rect 239140 293256 300582 293312
rect 300638 293256 300643 293312
rect 239140 293254 300643 293256
rect 239140 293252 239146 293254
rect 300577 293251 300643 293254
rect 3417 293178 3483 293181
rect -960 293176 3483 293178
rect -960 293120 3422 293176
rect 3478 293120 3483 293176
rect -960 293118 3483 293120
rect -960 293028 480 293118
rect 3417 293115 3483 293118
rect 235942 293116 235948 293180
rect 236012 293178 236018 293180
rect 297909 293178 297975 293181
rect 236012 293176 297975 293178
rect 236012 293120 297914 293176
rect 297970 293120 297975 293176
rect 236012 293118 297975 293120
rect 236012 293116 236018 293118
rect 297909 293115 297975 293118
rect 215886 292572 215892 292636
rect 215956 292634 215962 292636
rect 240869 292634 240935 292637
rect 215956 292632 240935 292634
rect 215956 292576 240874 292632
rect 240930 292576 240935 292632
rect 215956 292574 240935 292576
rect 215956 292572 215962 292574
rect 240869 292571 240935 292574
rect 242709 292498 242775 292501
rect 282126 292498 282132 292500
rect 242709 292496 282132 292498
rect 242709 292440 242714 292496
rect 242770 292440 282132 292496
rect 242709 292438 282132 292440
rect 242709 292435 242775 292438
rect 282126 292436 282132 292438
rect 282196 292436 282202 292500
rect 252645 292362 252711 292365
rect 253289 292362 253355 292365
rect 280654 292362 280660 292364
rect 238710 292360 253355 292362
rect 238710 292304 252650 292360
rect 252706 292304 253294 292360
rect 253350 292304 253355 292360
rect 238710 292302 253355 292304
rect 221038 292164 221044 292228
rect 221108 292226 221114 292228
rect 238710 292226 238770 292302
rect 252645 292299 252711 292302
rect 253289 292299 253355 292302
rect 258030 292302 280660 292362
rect 221108 292166 238770 292226
rect 251173 292226 251239 292229
rect 258030 292226 258090 292302
rect 280654 292300 280660 292302
rect 280724 292300 280730 292364
rect 251173 292224 258090 292226
rect 251173 292168 251178 292224
rect 251234 292168 258090 292224
rect 251173 292166 258090 292168
rect 221108 292164 221114 292166
rect 251173 292163 251239 292166
rect 218646 292028 218652 292092
rect 218716 292090 218722 292092
rect 251541 292090 251607 292093
rect 251909 292090 251975 292093
rect 218716 292088 251975 292090
rect 218716 292032 251546 292088
rect 251602 292032 251914 292088
rect 251970 292032 251975 292088
rect 218716 292030 251975 292032
rect 218716 292028 218722 292030
rect 251541 292027 251607 292030
rect 251909 292027 251975 292030
rect 249701 291954 249767 291957
rect 277894 291954 277900 291956
rect 249701 291952 277900 291954
rect 249701 291896 249706 291952
rect 249762 291896 277900 291952
rect 249701 291894 277900 291896
rect 249701 291891 249767 291894
rect 277894 291892 277900 291894
rect 277964 291892 277970 291956
rect 218053 291818 218119 291821
rect 219341 291818 219407 291821
rect 227713 291818 227779 291821
rect 218053 291816 227779 291818
rect 218053 291760 218058 291816
rect 218114 291760 219346 291816
rect 219402 291760 227718 291816
rect 227774 291760 227779 291816
rect 218053 291758 227779 291760
rect 218053 291755 218119 291758
rect 219341 291755 219407 291758
rect 227713 291755 227779 291758
rect 248086 291756 248092 291820
rect 248156 291818 248162 291820
rect 307845 291818 307911 291821
rect 248156 291816 307911 291818
rect 248156 291760 307850 291816
rect 307906 291760 307911 291816
rect 248156 291758 307911 291760
rect 248156 291756 248162 291758
rect 307845 291755 307911 291758
rect 310145 291818 310211 291821
rect 353886 291818 353892 291820
rect 310145 291816 353892 291818
rect 310145 291760 310150 291816
rect 310206 291760 353892 291816
rect 310145 291758 353892 291760
rect 310145 291755 310211 291758
rect 353886 291756 353892 291758
rect 353956 291756 353962 291820
rect 219985 291682 220051 291685
rect 247677 291682 247743 291685
rect 219985 291680 247743 291682
rect 219985 291624 219990 291680
rect 220046 291624 247682 291680
rect 247738 291624 247743 291680
rect 219985 291622 247743 291624
rect 219985 291619 220051 291622
rect 247677 291619 247743 291622
rect 220118 291484 220124 291548
rect 220188 291546 220194 291548
rect 250437 291546 250503 291549
rect 220188 291544 250503 291546
rect 220188 291488 250442 291544
rect 250498 291488 250503 291544
rect 220188 291486 250503 291488
rect 220188 291484 220194 291486
rect 250437 291483 250503 291486
rect 220302 291348 220308 291412
rect 220372 291410 220378 291412
rect 228357 291410 228423 291413
rect 220372 291408 228423 291410
rect 220372 291352 228362 291408
rect 228418 291352 228423 291408
rect 220372 291350 228423 291352
rect 220372 291348 220378 291350
rect 228357 291347 228423 291350
rect 221222 291212 221228 291276
rect 221292 291274 221298 291276
rect 226149 291274 226215 291277
rect 221292 291272 226215 291274
rect 221292 291216 226154 291272
rect 226210 291216 226215 291272
rect 221292 291214 226215 291216
rect 221292 291212 221298 291214
rect 226149 291211 226215 291214
rect 247677 291274 247743 291277
rect 248229 291274 248295 291277
rect 247677 291272 248295 291274
rect 247677 291216 247682 291272
rect 247738 291216 248234 291272
rect 248290 291216 248295 291272
rect 247677 291214 248295 291216
rect 247677 291211 247743 291214
rect 248229 291211 248295 291214
rect 250805 291138 250871 291141
rect 267089 291138 267155 291141
rect 250805 291136 267155 291138
rect 250805 291080 250810 291136
rect 250866 291080 267094 291136
rect 267150 291080 267155 291136
rect 250805 291078 267155 291080
rect 250805 291075 250871 291078
rect 267089 291075 267155 291078
rect 253054 290940 253060 291004
rect 253124 291002 253130 291004
rect 312118 291002 312124 291004
rect 253124 290942 312124 291002
rect 253124 290940 253130 290942
rect 312118 290940 312124 290942
rect 312188 290940 312194 291004
rect 245142 290804 245148 290868
rect 245212 290866 245218 290868
rect 304165 290866 304231 290869
rect 245212 290864 304231 290866
rect 245212 290808 304170 290864
rect 304226 290808 304231 290864
rect 245212 290806 304231 290808
rect 245212 290804 245218 290806
rect 304165 290803 304231 290806
rect 189165 290730 189231 290733
rect 246941 290730 247007 290733
rect 189165 290728 247007 290730
rect 189165 290672 189170 290728
rect 189226 290672 246946 290728
rect 247002 290672 247007 290728
rect 189165 290670 247007 290672
rect 189165 290667 189231 290670
rect 246941 290667 247007 290670
rect 253238 290668 253244 290732
rect 253308 290730 253314 290732
rect 313774 290730 313780 290732
rect 253308 290670 313780 290730
rect 253308 290668 253314 290670
rect 313774 290668 313780 290670
rect 313844 290668 313850 290732
rect 192017 290594 192083 290597
rect 251817 290594 251883 290597
rect 252093 290594 252159 290597
rect 192017 290592 252159 290594
rect 192017 290536 192022 290592
rect 192078 290536 251822 290592
rect 251878 290536 252098 290592
rect 252154 290536 252159 290592
rect 192017 290534 252159 290536
rect 192017 290531 192083 290534
rect 251817 290531 251883 290534
rect 252093 290531 252159 290534
rect 262070 290532 262076 290596
rect 262140 290594 262146 290596
rect 322749 290594 322815 290597
rect 262140 290592 322815 290594
rect 262140 290536 322754 290592
rect 322810 290536 322815 290592
rect 262140 290534 322815 290536
rect 262140 290532 262146 290534
rect 322749 290531 322815 290534
rect 220721 290458 220787 290461
rect 227621 290458 227687 290461
rect 220721 290456 227687 290458
rect 220721 290400 220726 290456
rect 220782 290400 227626 290456
rect 227682 290400 227687 290456
rect 220721 290398 227687 290400
rect 220721 290395 220787 290398
rect 227621 290395 227687 290398
rect 246246 290396 246252 290460
rect 246316 290458 246322 290460
rect 307569 290458 307635 290461
rect 246316 290456 307635 290458
rect 246316 290400 307574 290456
rect 307630 290400 307635 290456
rect 246316 290398 307635 290400
rect 246316 290396 246322 290398
rect 307569 290395 307635 290398
rect 224217 290186 224283 290189
rect 234153 290186 234219 290189
rect 238661 290186 238727 290189
rect 244273 290188 244339 290189
rect 238886 290186 238892 290188
rect 224217 290184 234219 290186
rect 224217 290128 224222 290184
rect 224278 290128 234158 290184
rect 234214 290128 234219 290184
rect 224217 290126 234219 290128
rect 238616 290184 238892 290186
rect 238616 290128 238666 290184
rect 238722 290128 238892 290184
rect 238616 290126 238892 290128
rect 224217 290123 224283 290126
rect 234153 290123 234219 290126
rect 238661 290123 238727 290126
rect 238886 290124 238892 290126
rect 238956 290124 238962 290188
rect 244222 290124 244228 290188
rect 244292 290186 244339 290188
rect 244292 290184 244384 290186
rect 244334 290128 244384 290184
rect 244292 290126 244384 290128
rect 244292 290124 244339 290126
rect 244273 290123 244339 290124
rect 190545 290050 190611 290053
rect 250621 290050 250687 290053
rect 190545 290048 250687 290050
rect 190545 289992 190550 290048
rect 190606 289992 250626 290048
rect 250682 289992 250687 290048
rect 190545 289990 250687 289992
rect 190545 289987 190611 289990
rect 250621 289987 250687 289990
rect 191833 289914 191899 289917
rect 224217 289914 224283 289917
rect 231577 289916 231643 289917
rect 191833 289912 224283 289914
rect 191833 289856 191838 289912
rect 191894 289856 224222 289912
rect 224278 289856 224283 289912
rect 191833 289854 224283 289856
rect 191833 289851 191899 289854
rect 224217 289851 224283 289854
rect 231526 289852 231532 289916
rect 231596 289914 231643 289916
rect 234153 289914 234219 289917
rect 251909 289914 251975 289917
rect 231596 289912 231688 289914
rect 231638 289856 231688 289912
rect 231596 289854 231688 289856
rect 234153 289912 251975 289914
rect 234153 289856 234158 289912
rect 234214 289856 251914 289912
rect 251970 289856 251975 289912
rect 234153 289854 251975 289856
rect 231596 289852 231643 289854
rect 231577 289851 231643 289852
rect 234153 289851 234219 289854
rect 251909 289851 251975 289854
rect 184197 289778 184263 289781
rect 241053 289778 241119 289781
rect 244222 289778 244228 289780
rect 184197 289776 241119 289778
rect 184197 289720 184202 289776
rect 184258 289720 241058 289776
rect 241114 289720 241119 289776
rect 184197 289718 241119 289720
rect 184197 289715 184263 289718
rect 241053 289715 241119 289718
rect 243862 289718 244228 289778
rect 186497 289642 186563 289645
rect 243862 289642 243922 289718
rect 244222 289716 244228 289718
rect 244292 289716 244298 289780
rect 244825 289778 244891 289781
rect 244414 289776 244891 289778
rect 244414 289720 244830 289776
rect 244886 289720 244891 289776
rect 244414 289718 244891 289720
rect 186497 289640 243922 289642
rect 186497 289584 186502 289640
rect 186558 289584 243922 289640
rect 186497 289582 243922 289584
rect 186497 289579 186563 289582
rect 186681 289506 186747 289509
rect 244414 289506 244474 289718
rect 244825 289715 244891 289718
rect 244958 289716 244964 289780
rect 245028 289778 245034 289780
rect 305453 289778 305519 289781
rect 245028 289776 305519 289778
rect 245028 289720 305458 289776
rect 305514 289720 305519 289776
rect 245028 289718 305519 289720
rect 245028 289716 245034 289718
rect 305453 289715 305519 289718
rect 248965 289642 249031 289645
rect 246622 289640 249031 289642
rect 246622 289584 248970 289640
rect 249026 289584 249031 289640
rect 246622 289582 249031 289584
rect 186681 289504 244474 289506
rect 186681 289448 186686 289504
rect 186742 289448 244474 289504
rect 186681 289446 244474 289448
rect 186681 289443 186747 289446
rect 245326 289444 245332 289508
rect 245396 289506 245402 289508
rect 245469 289506 245535 289509
rect 245396 289504 245535 289506
rect 245396 289448 245474 289504
rect 245530 289448 245535 289504
rect 245396 289446 245535 289448
rect 245396 289444 245402 289446
rect 245469 289443 245535 289446
rect 187785 289370 187851 289373
rect 246622 289370 246682 289582
rect 248965 289579 249031 289582
rect 247033 289506 247099 289509
rect 246990 289504 247099 289506
rect 246990 289448 247038 289504
rect 247094 289448 247099 289504
rect 246990 289443 247099 289448
rect 246990 289370 247050 289443
rect 247493 289370 247559 289373
rect 187785 289368 246682 289370
rect 187785 289312 187790 289368
rect 187846 289312 246682 289368
rect 187785 289310 246682 289312
rect 246806 289368 247559 289370
rect 246806 289312 247498 289368
rect 247554 289312 247559 289368
rect 246806 289310 247559 289312
rect 187785 289307 187851 289310
rect 186313 289234 186379 289237
rect 246806 289234 246866 289310
rect 247493 289307 247559 289310
rect 186313 289232 246866 289234
rect 186313 289176 186318 289232
rect 186374 289176 246866 289232
rect 186313 289174 246866 289176
rect 186313 289171 186379 289174
rect 249374 289172 249380 289236
rect 249444 289234 249450 289236
rect 310053 289234 310119 289237
rect 249444 289232 310119 289234
rect 249444 289176 310058 289232
rect 310114 289176 310119 289232
rect 249444 289174 310119 289176
rect 249444 289172 249450 289174
rect 310053 289171 310119 289174
rect 185025 289098 185091 289101
rect 245326 289098 245332 289100
rect 185025 289096 245332 289098
rect 185025 289040 185030 289096
rect 185086 289040 245332 289096
rect 185025 289038 245332 289040
rect 185025 289035 185091 289038
rect 245326 289036 245332 289038
rect 245396 289036 245402 289100
rect 231526 288356 231532 288420
rect 231596 288418 231602 288420
rect 274173 288418 274239 288421
rect 231596 288416 274239 288418
rect 231596 288360 274178 288416
rect 274234 288360 274239 288416
rect 231596 288358 274239 288360
rect 231596 288356 231602 288358
rect 274173 288355 274239 288358
rect 171317 287738 171383 287741
rect 231526 287738 231532 287740
rect 171317 287736 231532 287738
rect 171317 287680 171322 287736
rect 171378 287680 231532 287736
rect 171317 287678 231532 287680
rect 171317 287675 171383 287678
rect 231526 287676 231532 287678
rect 231596 287676 231602 287740
rect 269614 287676 269620 287740
rect 269684 287738 269690 287740
rect 323761 287738 323827 287741
rect 269684 287736 323827 287738
rect 269684 287680 323766 287736
rect 323822 287680 323827 287736
rect 269684 287678 323827 287680
rect 269684 287676 269690 287678
rect 323761 287675 323827 287678
rect 192109 286378 192175 286381
rect 221038 286378 221044 286380
rect 192109 286376 221044 286378
rect 192109 286320 192114 286376
rect 192170 286320 221044 286376
rect 192109 286318 221044 286320
rect 192109 286315 192175 286318
rect 221038 286316 221044 286318
rect 221108 286316 221114 286380
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 168465 278082 168531 278085
rect 220302 278082 220308 278084
rect 168465 278080 220308 278082
rect 168465 278024 168470 278080
rect 168526 278024 220308 278080
rect 168465 278022 220308 278024
rect 168465 278019 168531 278022
rect 220302 278020 220308 278022
rect 220372 278020 220378 278084
rect 190637 276722 190703 276725
rect 220118 276722 220124 276724
rect 190637 276720 220124 276722
rect 190637 276664 190642 276720
rect 190698 276664 220124 276720
rect 190637 276662 220124 276664
rect 190637 276659 190703 276662
rect 220118 276660 220124 276662
rect 220188 276660 220194 276724
rect 165797 275226 165863 275229
rect 221222 275226 221228 275228
rect 165797 275224 221228 275226
rect 165797 275168 165802 275224
rect 165858 275168 221228 275224
rect 165797 275166 221228 275168
rect 165797 275163 165863 275166
rect 221222 275164 221228 275166
rect 221292 275164 221298 275228
rect 271086 273804 271092 273868
rect 271156 273866 271162 273868
rect 322933 273866 322999 273869
rect 271156 273864 322999 273866
rect 271156 273808 322938 273864
rect 322994 273808 322999 273864
rect 271156 273806 322999 273808
rect 271156 273804 271162 273806
rect 322933 273803 322999 273806
rect 260598 272444 260604 272508
rect 260668 272506 260674 272508
rect 318926 272506 318932 272508
rect 260668 272446 318932 272506
rect 260668 272444 260674 272446
rect 318926 272444 318932 272446
rect 318996 272444 319002 272508
rect 580625 272234 580691 272237
rect 583520 272234 584960 272324
rect 580625 272232 584960 272234
rect 580625 272176 580630 272232
rect 580686 272176 584960 272232
rect 580625 272174 584960 272176
rect 580625 272171 580691 272174
rect 583520 272084 584960 272174
rect 266670 271084 266676 271148
rect 266740 271146 266746 271148
rect 326613 271146 326679 271149
rect 266740 271144 326679 271146
rect 266740 271088 326618 271144
rect 326674 271088 326679 271144
rect 266740 271086 326679 271088
rect 266740 271084 266746 271086
rect 326613 271083 326679 271086
rect 259310 268364 259316 268428
rect 259380 268426 259386 268428
rect 317638 268426 317644 268428
rect 259380 268366 317644 268426
rect 259380 268364 259386 268366
rect 317638 268364 317644 268366
rect 317708 268364 317714 268428
rect -960 267202 480 267292
rect 3049 267202 3115 267205
rect -960 267200 3115 267202
rect -960 267144 3054 267200
rect 3110 267144 3115 267200
rect -960 267142 3115 267144
rect -960 267052 480 267142
rect 3049 267139 3115 267142
rect 255630 267004 255636 267068
rect 255700 267066 255706 267068
rect 316861 267066 316927 267069
rect 255700 267064 316927 267066
rect 255700 267008 316866 267064
rect 316922 267008 316927 267064
rect 255700 267006 316927 267008
rect 255700 267004 255706 267006
rect 316861 267003 316927 267006
rect 268469 265570 268535 265573
rect 269113 265570 269179 265573
rect 268469 265568 269179 265570
rect 268469 265512 268474 265568
rect 268530 265512 269118 265568
rect 269174 265512 269179 265568
rect 268469 265510 269179 265512
rect 268469 265507 268535 265510
rect 269113 265507 269179 265510
rect 257102 264420 257108 264484
rect 257172 264482 257178 264484
rect 316350 264482 316356 264484
rect 257172 264422 316356 264482
rect 257172 264420 257178 264422
rect 316350 264420 316356 264422
rect 316420 264420 316426 264484
rect 264830 264284 264836 264348
rect 264900 264346 264906 264348
rect 325141 264346 325207 264349
rect 264900 264344 325207 264346
rect 264900 264288 325146 264344
rect 325202 264288 325207 264344
rect 264900 264286 325207 264288
rect 264900 264284 264906 264286
rect 325141 264283 325207 264286
rect 256366 264148 256372 264212
rect 256436 264210 256442 264212
rect 316769 264210 316835 264213
rect 256436 264208 316835 264210
rect 256436 264152 316774 264208
rect 316830 264152 316835 264208
rect 256436 264150 316835 264152
rect 256436 264148 256442 264150
rect 316769 264147 316835 264150
rect 259126 262788 259132 262852
rect 259196 262850 259202 262852
rect 318149 262850 318215 262853
rect 259196 262848 318215 262850
rect 259196 262792 318154 262848
rect 318210 262792 318215 262848
rect 259196 262790 318215 262792
rect 259196 262788 259202 262790
rect 318149 262787 318215 262790
rect 261886 261428 261892 261492
rect 261956 261490 261962 261492
rect 320398 261490 320404 261492
rect 261956 261430 320404 261490
rect 261956 261428 261962 261430
rect 320398 261428 320404 261430
rect 320468 261428 320474 261492
rect 267641 260130 267707 260133
rect 326521 260130 326587 260133
rect 267641 260128 326587 260130
rect 267641 260072 267646 260128
rect 267702 260072 326526 260128
rect 326582 260072 326587 260128
rect 267641 260070 326587 260072
rect 267641 260067 267707 260070
rect 326521 260067 326587 260070
rect 263542 258844 263548 258908
rect 263612 258906 263618 258908
rect 323342 258906 323348 258908
rect 263612 258846 323348 258906
rect 263612 258844 263618 258846
rect 323342 258844 323348 258846
rect 323412 258844 323418 258908
rect 580349 258906 580415 258909
rect 583520 258906 584960 258996
rect 580349 258904 584960 258906
rect 580349 258848 580354 258904
rect 580410 258848 584960 258904
rect 580349 258846 584960 258848
rect 580349 258843 580415 258846
rect 255446 258708 255452 258772
rect 255516 258770 255522 258772
rect 315389 258770 315455 258773
rect 255516 258768 315455 258770
rect 255516 258712 315394 258768
rect 315450 258712 315455 258768
rect 583520 258756 584960 258846
rect 255516 258710 315455 258712
rect 255516 258708 255522 258710
rect 315389 258707 315455 258710
rect 268561 257410 268627 257413
rect 269113 257410 269179 257413
rect 268561 257408 269179 257410
rect 268561 257352 268566 257408
rect 268622 257352 269118 257408
rect 269174 257352 269179 257408
rect 268561 257350 269179 257352
rect 268561 257347 268627 257350
rect 269113 257347 269179 257350
rect 260414 257212 260420 257276
rect 260484 257274 260490 257276
rect 321093 257274 321159 257277
rect 260484 257272 321159 257274
rect 260484 257216 321098 257272
rect 321154 257216 321159 257272
rect 260484 257214 321159 257216
rect 260484 257212 260490 257214
rect 321093 257211 321159 257214
rect 266118 255852 266124 255916
rect 266188 255914 266194 255916
rect 324446 255914 324452 255916
rect 266188 255854 324452 255914
rect 266188 255852 266194 255854
rect 324446 255852 324452 255854
rect 324516 255852 324522 255916
rect -960 254146 480 254236
rect 3417 254146 3483 254149
rect -960 254144 3483 254146
rect -960 254088 3422 254144
rect 3478 254088 3483 254144
rect -960 254086 3483 254088
rect -960 253996 480 254086
rect 3417 254083 3483 254086
rect 267406 253268 267412 253332
rect 267476 253330 267482 253332
rect 327165 253330 327231 253333
rect 267476 253328 327231 253330
rect 267476 253272 327170 253328
rect 327226 253272 327231 253328
rect 267476 253270 327231 253272
rect 267476 253268 267482 253270
rect 327165 253267 327231 253270
rect 261702 253132 261708 253196
rect 261772 253194 261778 253196
rect 322565 253194 322631 253197
rect 261772 253192 322631 253194
rect 261772 253136 322570 253192
rect 322626 253136 322631 253192
rect 261772 253134 322631 253136
rect 261772 253132 261778 253134
rect 322565 253131 322631 253134
rect 255998 251772 256004 251836
rect 256068 251834 256074 251836
rect 316677 251834 316743 251837
rect 256068 251832 316743 251834
rect 256068 251776 316682 251832
rect 316738 251776 316743 251832
rect 256068 251774 316743 251776
rect 256068 251772 256074 251774
rect 316677 251771 316743 251774
rect 269481 250746 269547 250749
rect 319529 250746 319595 250749
rect 269481 250744 319595 250746
rect 269481 250688 269486 250744
rect 269542 250688 319534 250744
rect 319590 250688 319595 250744
rect 269481 250686 319595 250688
rect 269481 250683 269547 250686
rect 319529 250683 319595 250686
rect 263542 250548 263548 250612
rect 263612 250610 263618 250612
rect 324630 250610 324636 250612
rect 263612 250550 324636 250610
rect 263612 250548 263618 250550
rect 324630 250548 324636 250550
rect 324700 250548 324706 250612
rect 267733 250474 267799 250477
rect 318241 250474 318307 250477
rect 267733 250472 318307 250474
rect 267733 250416 267738 250472
rect 267794 250416 318246 250472
rect 318302 250416 318307 250472
rect 267733 250414 318307 250416
rect 267733 250411 267799 250414
rect 318241 250411 318307 250414
rect 266118 249052 266124 249116
rect 266188 249114 266194 249116
rect 326337 249114 326403 249117
rect 266188 249112 326403 249114
rect 266188 249056 326342 249112
rect 326398 249056 326403 249112
rect 266188 249054 326403 249056
rect 266188 249052 266194 249054
rect 326337 249051 326403 249054
rect 258942 247964 258948 248028
rect 259012 248026 259018 248028
rect 290641 248026 290707 248029
rect 259012 248024 290707 248026
rect 259012 247968 290646 248024
rect 290702 247968 290707 248024
rect 259012 247966 290707 247968
rect 259012 247964 259018 247966
rect 290641 247963 290707 247966
rect 268745 247890 268811 247893
rect 327625 247890 327691 247893
rect 268745 247888 327691 247890
rect 268745 247832 268750 247888
rect 268806 247832 327630 247888
rect 327686 247832 327691 247888
rect 268745 247830 327691 247832
rect 268745 247827 268811 247830
rect 327625 247827 327691 247830
rect 263358 247692 263364 247756
rect 263428 247754 263434 247756
rect 323577 247754 323643 247757
rect 263428 247752 323643 247754
rect 263428 247696 323582 247752
rect 323638 247696 323643 247752
rect 263428 247694 323643 247696
rect 263428 247692 263434 247694
rect 323577 247691 323643 247694
rect 268009 247618 268075 247621
rect 321001 247618 321067 247621
rect 268009 247616 321067 247618
rect 268009 247560 268014 247616
rect 268070 247560 321006 247616
rect 321062 247560 321067 247616
rect 268009 247558 321067 247560
rect 268009 247555 268075 247558
rect 321001 247555 321067 247558
rect 265382 246604 265388 246668
rect 265452 246666 265458 246668
rect 269757 246666 269823 246669
rect 265452 246664 269823 246666
rect 265452 246608 269762 246664
rect 269818 246608 269823 246664
rect 265452 246606 269823 246608
rect 265452 246604 265458 246606
rect 269757 246603 269823 246606
rect 268837 246530 268903 246533
rect 317822 246530 317828 246532
rect 268837 246528 317828 246530
rect 268837 246472 268842 246528
rect 268898 246472 317828 246528
rect 268837 246470 317828 246472
rect 268837 246467 268903 246470
rect 317822 246468 317828 246470
rect 317892 246468 317898 246532
rect 221825 246394 221891 246397
rect 222009 246394 222075 246397
rect 221825 246392 222075 246394
rect 221825 246336 221830 246392
rect 221886 246336 222014 246392
rect 222070 246336 222075 246392
rect 221825 246334 222075 246336
rect 221825 246331 221891 246334
rect 222009 246331 222075 246334
rect 267917 246394 267983 246397
rect 322473 246394 322539 246397
rect 267917 246392 322539 246394
rect 267917 246336 267922 246392
rect 267978 246336 322478 246392
rect 322534 246336 322539 246392
rect 267917 246334 322539 246336
rect 267917 246331 267983 246334
rect 322473 246331 322539 246334
rect 266118 246196 266124 246260
rect 266188 246258 266194 246260
rect 326429 246258 326495 246261
rect 266188 246256 326495 246258
rect 266188 246200 326434 246256
rect 326490 246200 326495 246256
rect 266188 246198 326495 246200
rect 266188 246196 266194 246198
rect 326429 246195 326495 246198
rect 579613 245578 579679 245581
rect 583520 245578 584960 245668
rect 579613 245576 584960 245578
rect 579613 245520 579618 245576
rect 579674 245520 584960 245576
rect 579613 245518 584960 245520
rect 579613 245515 579679 245518
rect 583520 245428 584960 245518
rect 269941 245170 270007 245173
rect 323158 245170 323164 245172
rect 269941 245168 323164 245170
rect 269941 245112 269946 245168
rect 270002 245112 323164 245168
rect 269941 245110 323164 245112
rect 269941 245107 270007 245110
rect 323158 245108 323164 245110
rect 323228 245108 323234 245172
rect 264278 244972 264284 245036
rect 264348 245034 264354 245036
rect 325049 245034 325115 245037
rect 264348 245032 325115 245034
rect 264348 244976 325054 245032
rect 325110 244976 325115 245032
rect 264348 244974 325115 244976
rect 264348 244972 264354 244974
rect 325049 244971 325115 244974
rect 256918 244836 256924 244900
rect 256988 244898 256994 244900
rect 318057 244898 318123 244901
rect 256988 244896 318123 244898
rect 256988 244840 318062 244896
rect 318118 244840 318123 244896
rect 256988 244838 318123 244840
rect 256988 244836 256994 244838
rect 318057 244835 318123 244838
rect 268285 243674 268351 243677
rect 268469 243674 268535 243677
rect 268285 243672 268535 243674
rect 268285 243616 268290 243672
rect 268346 243616 268474 243672
rect 268530 243616 268535 243672
rect 268285 243614 268535 243616
rect 268285 243611 268351 243614
rect 268469 243611 268535 243614
rect 190729 243538 190795 243541
rect 218646 243538 218652 243540
rect 190729 243536 218652 243538
rect 190729 243480 190734 243536
rect 190790 243480 218652 243536
rect 190729 243478 218652 243480
rect 190729 243475 190795 243478
rect 218646 243476 218652 243478
rect 218716 243476 218722 243540
rect 268469 243538 268535 243541
rect 322197 243538 322263 243541
rect 268469 243536 322263 243538
rect 268469 243480 268474 243536
rect 268530 243480 322202 243536
rect 322258 243480 322263 243536
rect 268469 243478 322263 243480
rect 268469 243475 268535 243478
rect 322197 243475 322263 243478
rect 267406 242252 267412 242316
rect 267476 242314 267482 242316
rect 268101 242314 268167 242317
rect 267476 242312 268167 242314
rect 267476 242256 268106 242312
rect 268162 242256 268167 242312
rect 267476 242254 268167 242256
rect 267476 242252 267482 242254
rect 268101 242251 268167 242254
rect 259494 242116 259500 242180
rect 259564 242178 259570 242180
rect 319621 242178 319687 242181
rect 259564 242176 319687 242178
rect 259564 242120 319626 242176
rect 319682 242120 319687 242176
rect 259564 242118 319687 242120
rect 259564 242116 259570 242118
rect 319621 242115 319687 242118
rect 245694 241980 245700 242044
rect 245764 242042 245770 242044
rect 284385 242042 284451 242045
rect 245764 242040 284451 242042
rect 245764 241984 284390 242040
rect 284446 241984 284451 242040
rect 245764 241982 284451 241984
rect 245764 241980 245770 241982
rect 284385 241979 284451 241982
rect 153009 241906 153075 241909
rect 221181 241906 221247 241909
rect 153009 241904 221247 241906
rect 153009 241848 153014 241904
rect 153070 241848 221186 241904
rect 221242 241848 221247 241904
rect 153009 241846 221247 241848
rect 153009 241843 153075 241846
rect 221181 241843 221247 241846
rect 241830 241844 241836 241908
rect 241900 241906 241906 241908
rect 267549 241906 267615 241909
rect 241900 241904 267615 241906
rect 241900 241848 267554 241904
rect 267610 241848 267615 241904
rect 241900 241846 267615 241848
rect 241900 241844 241906 241846
rect 267549 241843 267615 241846
rect 151721 241770 151787 241773
rect 222694 241770 222700 241772
rect 151721 241768 222700 241770
rect 151721 241712 151726 241768
rect 151782 241712 222700 241768
rect 151721 241710 222700 241712
rect 151721 241707 151787 241710
rect 222694 241708 222700 241710
rect 222764 241708 222770 241772
rect 252686 241708 252692 241772
rect 252756 241770 252762 241772
rect 270125 241770 270191 241773
rect 252756 241768 270191 241770
rect 252756 241712 270130 241768
rect 270186 241712 270191 241768
rect 252756 241710 270191 241712
rect 252756 241708 252762 241710
rect 270125 241707 270191 241710
rect 151629 241634 151695 241637
rect 225454 241634 225460 241636
rect 151629 241632 225460 241634
rect 151629 241576 151634 241632
rect 151690 241576 225460 241632
rect 151629 241574 225460 241576
rect 151629 241571 151695 241574
rect 225454 241572 225460 241574
rect 225524 241572 225530 241636
rect 257286 241572 257292 241636
rect 257356 241634 257362 241636
rect 267733 241634 267799 241637
rect 257356 241632 267799 241634
rect 257356 241576 267738 241632
rect 267794 241576 267799 241632
rect 257356 241574 267799 241576
rect 257356 241572 257362 241574
rect 267733 241571 267799 241574
rect 268193 241634 268259 241637
rect 269614 241634 269620 241636
rect 268193 241632 269620 241634
rect 268193 241576 268198 241632
rect 268254 241576 269620 241632
rect 268193 241574 269620 241576
rect 268193 241571 268259 241574
rect 269614 241572 269620 241574
rect 269684 241572 269690 241636
rect 225638 241436 225644 241500
rect 225708 241498 225714 241500
rect 247534 241498 247540 241500
rect 225708 241438 247540 241498
rect 225708 241436 225714 241438
rect 247534 241436 247540 241438
rect 247604 241436 247610 241500
rect 258574 241436 258580 241500
rect 258644 241498 258650 241500
rect 269573 241498 269639 241501
rect 258644 241496 269639 241498
rect 258644 241440 269578 241496
rect 269634 241440 269639 241496
rect 258644 241438 269639 241440
rect 258644 241436 258650 241438
rect 269573 241435 269639 241438
rect 224166 241300 224172 241364
rect 224236 241362 224242 241364
rect 274541 241362 274607 241365
rect 224236 241360 274607 241362
rect 224236 241304 274546 241360
rect 274602 241304 274607 241360
rect 224236 241302 274607 241304
rect 224236 241300 224242 241302
rect 274541 241299 274607 241302
rect 217409 241226 217475 241229
rect 217409 241224 230674 241226
rect -960 241090 480 241180
rect 217409 241168 217414 241224
rect 217470 241168 230674 241224
rect 217409 241166 230674 241168
rect 217409 241163 217475 241166
rect 3325 241090 3391 241093
rect -960 241088 3391 241090
rect -960 241032 3330 241088
rect 3386 241032 3391 241088
rect -960 241030 3391 241032
rect 230614 241090 230674 241166
rect 230790 241164 230796 241228
rect 230860 241226 230866 241228
rect 284109 241226 284175 241229
rect 230860 241224 284175 241226
rect 230860 241168 284114 241224
rect 284170 241168 284175 241224
rect 230860 241166 284175 241168
rect 230860 241164 230866 241166
rect 284109 241163 284175 241166
rect 232078 241090 232084 241092
rect 230614 241030 232084 241090
rect -960 240940 480 241030
rect 3325 241027 3391 241030
rect 232078 241028 232084 241030
rect 232148 241028 232154 241092
rect 233366 241028 233372 241092
rect 233436 241090 233442 241092
rect 292614 241090 292620 241092
rect 233436 241030 292620 241090
rect 233436 241028 233442 241030
rect 292614 241028 292620 241030
rect 292684 241028 292690 241092
rect 157241 240954 157307 240957
rect 206369 240954 206435 240957
rect 221457 240954 221523 240957
rect 157241 240952 221523 240954
rect 157241 240896 157246 240952
rect 157302 240896 206374 240952
rect 206430 240896 221462 240952
rect 221518 240896 221523 240952
rect 157241 240894 221523 240896
rect 157241 240891 157307 240894
rect 206369 240891 206435 240894
rect 221457 240891 221523 240894
rect 227662 240892 227668 240956
rect 227732 240954 227738 240956
rect 284753 240954 284819 240957
rect 227732 240952 284819 240954
rect 227732 240896 284758 240952
rect 284814 240896 284819 240952
rect 227732 240894 284819 240896
rect 227732 240892 227738 240894
rect 284753 240891 284819 240894
rect 152917 240818 152983 240821
rect 209589 240818 209655 240821
rect 229134 240818 229140 240820
rect 152917 240816 229140 240818
rect 152917 240760 152922 240816
rect 152978 240760 209594 240816
rect 209650 240760 229140 240816
rect 152917 240758 229140 240760
rect 152917 240755 152983 240758
rect 209589 240755 209655 240758
rect 229134 240756 229140 240758
rect 229204 240756 229210 240820
rect 234838 240756 234844 240820
rect 234908 240818 234914 240820
rect 294454 240818 294460 240820
rect 234908 240758 294460 240818
rect 234908 240756 234914 240758
rect 294454 240756 294460 240758
rect 294524 240756 294530 240820
rect 157057 240682 157123 240685
rect 222193 240682 222259 240685
rect 233182 240682 233188 240684
rect 157057 240680 222072 240682
rect 157057 240624 157062 240680
rect 157118 240624 222072 240680
rect 157057 240622 222072 240624
rect 157057 240619 157123 240622
rect 222012 240546 222072 240622
rect 222193 240680 233188 240682
rect 222193 240624 222198 240680
rect 222254 240624 233188 240680
rect 222193 240622 233188 240624
rect 222193 240619 222259 240622
rect 233182 240620 233188 240622
rect 233252 240620 233258 240684
rect 233734 240620 233740 240684
rect 233804 240682 233810 240684
rect 234470 240682 234476 240684
rect 233804 240622 234476 240682
rect 233804 240620 233810 240622
rect 234470 240620 234476 240622
rect 234540 240620 234546 240684
rect 237966 240620 237972 240684
rect 238036 240682 238042 240684
rect 258390 240682 258396 240684
rect 238036 240622 258396 240682
rect 238036 240620 238042 240622
rect 258390 240620 258396 240622
rect 258460 240620 258466 240684
rect 259862 240620 259868 240684
rect 259932 240682 259938 240684
rect 268837 240682 268903 240685
rect 274582 240682 274588 240684
rect 259932 240680 268903 240682
rect 259932 240624 268842 240680
rect 268898 240624 268903 240680
rect 259932 240622 268903 240624
rect 259932 240620 259938 240622
rect 268837 240619 268903 240622
rect 273210 240622 274588 240682
rect 224166 240546 224172 240548
rect 222012 240486 224172 240546
rect 224166 240484 224172 240486
rect 224236 240484 224242 240548
rect 230422 240484 230428 240548
rect 230492 240546 230498 240548
rect 237782 240546 237788 240548
rect 230492 240486 237788 240546
rect 230492 240484 230498 240486
rect 237782 240484 237788 240486
rect 237852 240484 237858 240548
rect 269297 240546 269363 240549
rect 256650 240544 269363 240546
rect 256650 240488 269302 240544
rect 269358 240488 269363 240544
rect 256650 240486 269363 240488
rect 213453 240410 213519 240413
rect 222285 240410 222351 240413
rect 213453 240408 222351 240410
rect 213453 240352 213458 240408
rect 213514 240352 222290 240408
rect 222346 240352 222351 240408
rect 213453 240350 222351 240352
rect 213453 240347 213519 240350
rect 222285 240347 222351 240350
rect 222510 240348 222516 240412
rect 222580 240410 222586 240412
rect 232998 240410 233004 240412
rect 222580 240350 233004 240410
rect 222580 240348 222586 240350
rect 232998 240348 233004 240350
rect 233068 240348 233074 240412
rect 222101 240274 222167 240277
rect 239806 240274 239812 240276
rect 222101 240272 239812 240274
rect 222101 240216 222106 240272
rect 222162 240216 239812 240272
rect 222101 240214 239812 240216
rect 222101 240211 222167 240214
rect 239806 240212 239812 240214
rect 239876 240212 239882 240276
rect 256650 240274 256710 240486
rect 269297 240483 269363 240486
rect 265198 240348 265204 240412
rect 265268 240410 265274 240412
rect 273210 240410 273270 240622
rect 274582 240620 274588 240622
rect 274652 240620 274658 240684
rect 265268 240350 273270 240410
rect 265268 240348 265274 240350
rect 255270 240214 256710 240274
rect 225094 240078 227914 240138
rect 218881 240002 218947 240005
rect 222510 240002 222516 240004
rect 218881 240000 222516 240002
rect 218881 239944 218886 240000
rect 218942 239944 222516 240000
rect 218881 239942 222516 239944
rect 218881 239939 218947 239942
rect 222510 239940 222516 239942
rect 222580 239940 222586 240004
rect 223062 240002 223068 240004
rect 222702 239942 223068 240002
rect 222193 239866 222259 239869
rect 222702 239866 222762 239942
rect 223062 239940 223068 239942
rect 223132 240002 223138 240004
rect 223132 239942 223544 240002
rect 223132 239940 223138 239942
rect 223484 239869 223544 239942
rect 223798 239940 223804 240004
rect 223868 239940 223874 240004
rect 223982 239940 223988 240004
rect 224052 240002 224058 240004
rect 224052 239942 224970 240002
rect 224052 239940 224058 239942
rect 222193 239864 222762 239866
rect 222193 239808 222198 239864
rect 222254 239808 222762 239864
rect 222193 239806 222762 239808
rect 222883 239866 222949 239869
rect 223246 239866 223252 239868
rect 222883 239864 223252 239866
rect 222883 239808 222888 239864
rect 222944 239808 223252 239864
rect 222883 239806 223252 239808
rect 222193 239803 222259 239806
rect 222883 239803 222949 239806
rect 223246 239804 223252 239806
rect 223316 239804 223322 239868
rect 223484 239864 223593 239869
rect 223484 239808 223532 239864
rect 223588 239808 223593 239864
rect 223484 239806 223593 239808
rect 223806 239866 223866 239940
rect 224910 239869 224970 239942
rect 225094 239869 225154 240078
rect 226374 239940 226380 240004
rect 226444 240002 226450 240004
rect 227854 240002 227914 240078
rect 230974 240076 230980 240140
rect 231044 240138 231050 240140
rect 241830 240138 241836 240140
rect 231044 240078 241836 240138
rect 231044 240076 231050 240078
rect 241830 240076 241836 240078
rect 241900 240076 241906 240140
rect 242014 240076 242020 240140
rect 242084 240138 242090 240140
rect 246246 240138 246252 240140
rect 242084 240078 246252 240138
rect 242084 240076 242090 240078
rect 246246 240076 246252 240078
rect 246316 240138 246322 240140
rect 246316 240078 247050 240138
rect 246316 240076 246322 240078
rect 236678 240002 236684 240004
rect 226444 239942 227730 240002
rect 227854 239942 234630 240002
rect 226444 239940 226450 239942
rect 227670 239869 227730 239942
rect 223987 239866 224053 239869
rect 223806 239864 224053 239866
rect 223806 239808 223992 239864
rect 224048 239808 224053 239864
rect 223806 239806 224053 239808
rect 223527 239803 223593 239806
rect 223987 239803 224053 239806
rect 224125 239868 224191 239869
rect 224125 239864 224172 239868
rect 224236 239866 224242 239868
rect 224355 239866 224421 239869
rect 224718 239866 224724 239868
rect 224125 239808 224130 239864
rect 224125 239804 224172 239808
rect 224236 239806 224282 239866
rect 224355 239864 224724 239866
rect 224355 239808 224360 239864
rect 224416 239808 224724 239864
rect 224355 239806 224724 239808
rect 224236 239804 224242 239806
rect 224125 239803 224191 239804
rect 224355 239803 224421 239806
rect 224718 239804 224724 239806
rect 224788 239804 224794 239868
rect 224907 239864 224973 239869
rect 225091 239868 225157 239869
rect 224907 239808 224912 239864
rect 224968 239808 224973 239864
rect 224907 239803 224973 239808
rect 225086 239804 225092 239868
rect 225156 239866 225162 239868
rect 225781 239866 225847 239869
rect 226190 239866 226196 239868
rect 225156 239806 225248 239866
rect 225781 239864 226196 239866
rect 225781 239808 225786 239864
rect 225842 239808 226196 239864
rect 225781 239806 226196 239808
rect 225156 239804 225162 239806
rect 225091 239803 225157 239804
rect 225781 239803 225847 239806
rect 226190 239804 226196 239806
rect 226260 239804 226266 239868
rect 226563 239866 226629 239869
rect 227294 239866 227300 239868
rect 226563 239864 227300 239866
rect 226563 239808 226568 239864
rect 226624 239808 227300 239864
rect 226563 239806 227300 239808
rect 226563 239803 226629 239806
rect 227294 239804 227300 239806
rect 227364 239804 227370 239868
rect 227667 239864 227733 239869
rect 227667 239808 227672 239864
rect 227728 239808 227733 239864
rect 227667 239803 227733 239808
rect 228127 239866 228193 239869
rect 228449 239866 228515 239869
rect 229231 239866 229297 239869
rect 228127 239864 228236 239866
rect 228127 239808 228132 239864
rect 228188 239808 228236 239864
rect 228127 239803 228236 239808
rect 228449 239864 229297 239866
rect 228449 239808 228454 239864
rect 228510 239808 229236 239864
rect 229292 239808 229297 239864
rect 228449 239806 229297 239808
rect 228449 239803 228515 239806
rect 229231 239803 229297 239806
rect 229502 239804 229508 239868
rect 229572 239866 229578 239868
rect 229783 239866 229849 239869
rect 229572 239864 229849 239866
rect 229572 239808 229788 239864
rect 229844 239808 229849 239864
rect 229572 239806 229849 239808
rect 229572 239804 229578 239806
rect 229783 239803 229849 239806
rect 230054 239804 230060 239868
rect 230124 239866 230130 239868
rect 230335 239866 230401 239869
rect 230124 239864 230401 239866
rect 230124 239808 230340 239864
rect 230396 239808 230401 239864
rect 230124 239806 230401 239808
rect 230124 239804 230130 239806
rect 230335 239803 230401 239806
rect 230795 239866 230861 239869
rect 230974 239866 230980 239868
rect 230795 239864 230980 239866
rect 230795 239808 230800 239864
rect 230856 239808 230980 239864
rect 230795 239806 230980 239808
rect 230795 239803 230861 239806
rect 230974 239804 230980 239806
rect 231044 239804 231050 239868
rect 231163 239866 231229 239869
rect 231710 239866 231716 239868
rect 231163 239864 231716 239866
rect 231163 239808 231168 239864
rect 231224 239808 231716 239864
rect 231163 239806 231716 239808
rect 231163 239803 231229 239806
rect 231710 239804 231716 239806
rect 231780 239804 231786 239868
rect 231899 239866 231965 239869
rect 232630 239866 232636 239868
rect 231899 239864 232636 239866
rect 231899 239808 231904 239864
rect 231960 239808 232636 239864
rect 231899 239806 232636 239808
rect 231899 239803 231965 239806
rect 232630 239804 232636 239806
rect 232700 239804 232706 239868
rect 232814 239804 232820 239868
rect 232884 239866 232890 239868
rect 233187 239866 233253 239869
rect 233417 239868 233483 239869
rect 232884 239864 233253 239866
rect 232884 239808 233192 239864
rect 233248 239808 233253 239864
rect 232884 239806 233253 239808
rect 232884 239804 232890 239806
rect 233187 239803 233253 239806
rect 233366 239804 233372 239868
rect 233436 239866 233483 239868
rect 233436 239864 233528 239866
rect 233478 239808 233528 239864
rect 233436 239806 233528 239808
rect 233436 239804 233483 239806
rect 233918 239804 233924 239868
rect 233988 239866 233994 239868
rect 234291 239866 234357 239869
rect 233988 239864 234357 239866
rect 233988 239808 234296 239864
rect 234352 239808 234357 239864
rect 233988 239806 234357 239808
rect 233988 239804 233994 239806
rect 233417 239803 233483 239804
rect 234291 239803 234357 239806
rect 155769 239730 155835 239733
rect 210325 239730 210391 239733
rect 210785 239730 210851 239733
rect 155769 239728 210851 239730
rect 155769 239672 155774 239728
rect 155830 239672 210330 239728
rect 210386 239672 210790 239728
rect 210846 239672 210851 239728
rect 155769 239670 210851 239672
rect 155769 239667 155835 239670
rect 210325 239667 210391 239670
rect 210785 239667 210851 239670
rect 222377 239730 222443 239733
rect 223430 239730 223436 239732
rect 222377 239728 223436 239730
rect 222377 239672 222382 239728
rect 222438 239672 223436 239728
rect 222377 239670 223436 239672
rect 222377 239667 222443 239670
rect 223430 239668 223436 239670
rect 223500 239668 223506 239732
rect 223614 239668 223620 239732
rect 223684 239730 223690 239732
rect 223849 239730 223915 239733
rect 223684 239728 223915 239730
rect 223684 239672 223854 239728
rect 223910 239672 223915 239728
rect 223684 239670 223915 239672
rect 223684 239668 223690 239670
rect 223849 239667 223915 239670
rect 225094 239670 226258 239730
rect 155861 239594 155927 239597
rect 213085 239594 213151 239597
rect 155861 239592 213151 239594
rect 155861 239536 155866 239592
rect 155922 239536 213090 239592
rect 213146 239536 213151 239592
rect 155861 239534 213151 239536
rect 155861 239531 155927 239534
rect 213085 239531 213151 239534
rect 219985 239594 220051 239597
rect 225094 239594 225154 239670
rect 219985 239592 225154 239594
rect 219985 239536 219990 239592
rect 220046 239536 225154 239592
rect 219985 239534 225154 239536
rect 219985 239531 220051 239534
rect 225270 239532 225276 239596
rect 225340 239594 225346 239596
rect 225689 239594 225755 239597
rect 225340 239592 225755 239594
rect 225340 239536 225694 239592
rect 225750 239536 225755 239592
rect 225340 239534 225755 239536
rect 225340 239532 225346 239534
rect 225689 239531 225755 239534
rect 155493 239458 155559 239461
rect 207841 239458 207907 239461
rect 221457 239458 221523 239461
rect 155493 239456 221523 239458
rect 155493 239400 155498 239456
rect 155554 239400 207846 239456
rect 207902 239400 221462 239456
rect 221518 239400 221523 239456
rect 155493 239398 221523 239400
rect 155493 239395 155559 239398
rect 207841 239395 207907 239398
rect 221457 239395 221523 239398
rect 222694 239396 222700 239460
rect 222764 239458 222770 239460
rect 223481 239458 223547 239461
rect 222764 239456 223547 239458
rect 222764 239400 223486 239456
rect 223542 239400 223547 239456
rect 222764 239398 223547 239400
rect 222764 239396 222770 239398
rect 223481 239395 223547 239398
rect 225321 239458 225387 239461
rect 226006 239458 226012 239460
rect 225321 239456 226012 239458
rect 225321 239400 225326 239456
rect 225382 239400 226012 239456
rect 225321 239398 226012 239400
rect 225321 239395 225387 239398
rect 226006 239396 226012 239398
rect 226076 239396 226082 239460
rect 210785 239322 210851 239325
rect 220905 239322 220971 239325
rect 210785 239320 220971 239322
rect 210785 239264 210790 239320
rect 210846 239264 220910 239320
rect 220966 239264 220971 239320
rect 210785 239262 220971 239264
rect 210785 239259 210851 239262
rect 220905 239259 220971 239262
rect 225505 239322 225571 239325
rect 225638 239322 225644 239324
rect 225505 239320 225644 239322
rect 225505 239264 225510 239320
rect 225566 239264 225644 239320
rect 225505 239262 225644 239264
rect 225505 239259 225571 239262
rect 225638 239260 225644 239262
rect 225708 239260 225714 239324
rect 226198 239322 226258 239670
rect 226742 239668 226748 239732
rect 226812 239730 226818 239732
rect 227023 239730 227089 239733
rect 226812 239728 227089 239730
rect 226812 239672 227028 239728
rect 227084 239672 227089 239728
rect 226812 239670 227089 239672
rect 226812 239668 226818 239670
rect 227023 239667 227089 239670
rect 227437 239730 227503 239733
rect 227662 239730 227668 239732
rect 227437 239728 227668 239730
rect 227437 239672 227442 239728
rect 227498 239672 227668 239728
rect 227437 239670 227668 239672
rect 227437 239667 227503 239670
rect 227662 239668 227668 239670
rect 227732 239668 227738 239732
rect 227989 239730 228055 239733
rect 228176 239730 228236 239803
rect 227989 239728 228236 239730
rect 227989 239672 227994 239728
rect 228050 239672 228236 239728
rect 227989 239670 228236 239672
rect 228357 239730 228423 239733
rect 228582 239730 228588 239732
rect 228357 239728 228588 239730
rect 228357 239672 228362 239728
rect 228418 239672 228588 239728
rect 228357 239670 228588 239672
rect 227989 239667 228055 239670
rect 228357 239667 228423 239670
rect 228582 239668 228588 239670
rect 228652 239668 228658 239732
rect 229134 239668 229140 239732
rect 229204 239730 229210 239732
rect 229277 239730 229343 239733
rect 229204 239728 229343 239730
rect 229204 239672 229282 239728
rect 229338 239672 229343 239728
rect 229204 239670 229343 239672
rect 229204 239668 229210 239670
rect 229277 239667 229343 239670
rect 229461 239730 229527 239733
rect 229870 239730 229876 239732
rect 229461 239728 229876 239730
rect 229461 239672 229466 239728
rect 229522 239672 229876 239728
rect 229461 239670 229876 239672
rect 229461 239667 229527 239670
rect 229870 239668 229876 239670
rect 229940 239668 229946 239732
rect 230289 239730 230355 239733
rect 230790 239730 230796 239732
rect 230289 239728 230796 239730
rect 230289 239672 230294 239728
rect 230350 239672 230796 239728
rect 230289 239670 230796 239672
rect 230289 239667 230355 239670
rect 230790 239668 230796 239670
rect 230860 239668 230866 239732
rect 231117 239730 231183 239733
rect 231485 239732 231551 239733
rect 231342 239730 231348 239732
rect 231117 239728 231348 239730
rect 231117 239672 231122 239728
rect 231178 239672 231348 239728
rect 231117 239670 231348 239672
rect 231117 239667 231183 239670
rect 231342 239668 231348 239670
rect 231412 239668 231418 239732
rect 231485 239728 231532 239732
rect 231596 239730 231602 239732
rect 231485 239672 231490 239728
rect 231485 239668 231532 239672
rect 231596 239670 231642 239730
rect 231596 239668 231602 239670
rect 232078 239668 232084 239732
rect 232148 239730 232154 239732
rect 232313 239730 232379 239733
rect 232148 239728 232379 239730
rect 232148 239672 232318 239728
rect 232374 239672 232379 239728
rect 232148 239670 232379 239672
rect 232148 239668 232154 239670
rect 231485 239667 231551 239668
rect 232313 239667 232379 239670
rect 233182 239668 233188 239732
rect 233252 239730 233258 239732
rect 233417 239730 233483 239733
rect 233693 239732 233759 239733
rect 233693 239730 233740 239732
rect 233252 239728 233483 239730
rect 233252 239672 233422 239728
rect 233478 239672 233483 239728
rect 233252 239670 233483 239672
rect 233648 239728 233740 239730
rect 233648 239672 233698 239728
rect 233648 239670 233740 239672
rect 233252 239668 233258 239670
rect 233417 239667 233483 239670
rect 233693 239668 233740 239670
rect 233804 239668 233810 239732
rect 234102 239668 234108 239732
rect 234172 239730 234178 239732
rect 234429 239730 234495 239733
rect 234172 239728 234495 239730
rect 234172 239672 234434 239728
rect 234490 239672 234495 239728
rect 234172 239670 234495 239672
rect 234172 239668 234178 239670
rect 233693 239667 233759 239668
rect 234429 239667 234495 239670
rect 226374 239532 226380 239596
rect 226444 239594 226450 239596
rect 226517 239594 226583 239597
rect 228633 239594 228699 239597
rect 226444 239592 226583 239594
rect 226444 239536 226522 239592
rect 226578 239536 226583 239592
rect 226444 239534 226583 239536
rect 226444 239532 226450 239534
rect 226517 239531 226583 239534
rect 227992 239592 228699 239594
rect 227992 239536 228638 239592
rect 228694 239536 228699 239592
rect 227992 239534 228699 239536
rect 226558 239396 226564 239460
rect 226628 239458 226634 239460
rect 226977 239458 227043 239461
rect 226628 239456 227043 239458
rect 226628 239400 226982 239456
rect 227038 239400 227043 239456
rect 226628 239398 227043 239400
rect 226628 239396 226634 239398
rect 226977 239395 227043 239398
rect 227437 239460 227503 239461
rect 227437 239456 227484 239460
rect 227548 239458 227554 239460
rect 227437 239400 227442 239456
rect 227437 239396 227484 239400
rect 227548 239398 227594 239458
rect 227548 239396 227554 239398
rect 227846 239396 227852 239460
rect 227916 239458 227922 239460
rect 227992 239458 228052 239534
rect 228633 239531 228699 239534
rect 228950 239532 228956 239596
rect 229020 239594 229026 239596
rect 229277 239594 229343 239597
rect 229553 239596 229619 239597
rect 229020 239592 229343 239594
rect 229020 239536 229282 239592
rect 229338 239536 229343 239592
rect 229020 239534 229343 239536
rect 229020 239532 229026 239534
rect 229277 239531 229343 239534
rect 229502 239532 229508 239596
rect 229572 239594 229619 239596
rect 229572 239592 229664 239594
rect 229614 239536 229664 239592
rect 229572 239534 229664 239536
rect 229572 239532 229619 239534
rect 231158 239532 231164 239596
rect 231228 239594 231234 239596
rect 231761 239594 231827 239597
rect 231228 239592 231827 239594
rect 231228 239536 231766 239592
rect 231822 239536 231827 239592
rect 231228 239534 231827 239536
rect 231228 239532 231234 239534
rect 229553 239531 229619 239532
rect 231761 239531 231827 239534
rect 231945 239594 232011 239597
rect 232262 239594 232268 239596
rect 231945 239592 232268 239594
rect 231945 239536 231950 239592
rect 232006 239536 232268 239592
rect 231945 239534 232268 239536
rect 231945 239531 232011 239534
rect 232262 239532 232268 239534
rect 232332 239594 232338 239596
rect 232865 239594 232931 239597
rect 232332 239592 232931 239594
rect 232332 239536 232870 239592
rect 232926 239536 232931 239592
rect 232332 239534 232931 239536
rect 232332 239532 232338 239534
rect 232865 239531 232931 239534
rect 232998 239532 233004 239596
rect 233068 239594 233074 239596
rect 233325 239594 233391 239597
rect 233068 239592 233391 239594
rect 233068 239536 233330 239592
rect 233386 239536 233391 239592
rect 233068 239534 233391 239536
rect 234570 239594 234630 239942
rect 236318 239942 236684 240002
rect 236318 239869 236378 239942
rect 236678 239940 236684 239942
rect 236748 239940 236754 240004
rect 239622 240002 239628 240004
rect 238710 239942 239628 240002
rect 237327 239900 237393 239903
rect 237284 239898 237393 239900
rect 234843 239868 234909 239869
rect 234838 239866 234844 239868
rect 234752 239806 234844 239866
rect 234838 239804 234844 239806
rect 234908 239804 234914 239868
rect 236315 239864 236381 239869
rect 236315 239808 236320 239864
rect 236376 239808 236381 239864
rect 234843 239803 234909 239804
rect 236315 239803 236381 239808
rect 236499 239864 236565 239869
rect 236499 239808 236504 239864
rect 236560 239808 236565 239864
rect 236499 239803 236565 239808
rect 236862 239804 236868 239868
rect 236932 239866 236938 239868
rect 237284 239866 237332 239898
rect 236932 239842 237332 239866
rect 237388 239842 237393 239898
rect 238523 239898 238589 239903
rect 236932 239837 237393 239842
rect 236932 239806 237344 239837
rect 236932 239804 236938 239806
rect 237966 239804 237972 239868
rect 238036 239866 238042 239868
rect 238523 239866 238528 239898
rect 238036 239842 238528 239866
rect 238584 239842 238589 239898
rect 238036 239837 238589 239842
rect 238710 239866 238770 239942
rect 239622 239940 239628 239942
rect 239692 239940 239698 240004
rect 241191 239900 241257 239903
rect 241148 239898 241257 239900
rect 238891 239866 238957 239869
rect 238710 239864 238957 239866
rect 238036 239806 238586 239837
rect 238710 239808 238896 239864
rect 238952 239808 238957 239864
rect 238710 239806 238957 239808
rect 238036 239804 238042 239806
rect 238891 239803 238957 239806
rect 239070 239804 239076 239868
rect 239140 239866 239146 239868
rect 239535 239866 239601 239869
rect 239140 239864 239601 239866
rect 239140 239808 239540 239864
rect 239596 239808 239601 239864
rect 239140 239806 239601 239808
rect 239140 239804 239146 239806
rect 239535 239803 239601 239806
rect 240174 239804 240180 239868
rect 240244 239866 240250 239868
rect 240363 239866 240429 239869
rect 240244 239864 240429 239866
rect 240244 239808 240368 239864
rect 240424 239808 240429 239864
rect 240244 239806 240429 239808
rect 240244 239804 240250 239806
rect 240363 239803 240429 239806
rect 240542 239804 240548 239868
rect 240612 239866 240618 239868
rect 240823 239866 240889 239869
rect 241148 239868 241196 239898
rect 240612 239864 240889 239866
rect 240612 239808 240828 239864
rect 240884 239808 240889 239864
rect 240612 239806 240889 239808
rect 240612 239804 240618 239806
rect 240823 239803 240889 239806
rect 241094 239804 241100 239868
rect 241164 239842 241196 239868
rect 241252 239842 241257 239898
rect 243123 239898 243189 239903
rect 241164 239837 241257 239842
rect 241697 239866 241763 239869
rect 242111 239866 242177 239869
rect 241697 239864 242177 239866
rect 241164 239806 241208 239837
rect 241697 239808 241702 239864
rect 241758 239808 242116 239864
rect 242172 239808 242177 239864
rect 243123 239842 243128 239898
rect 243184 239842 243189 239898
rect 246343 239900 246409 239903
rect 246343 239898 246452 239900
rect 243123 239837 243189 239842
rect 244733 239866 244799 239869
rect 244958 239866 244964 239868
rect 244733 239864 244964 239866
rect 241697 239806 242177 239808
rect 241164 239804 241170 239806
rect 241697 239803 241763 239806
rect 242111 239803 242177 239806
rect 236502 239733 236562 239803
rect 235073 239732 235139 239733
rect 235022 239730 235028 239732
rect 234982 239670 235028 239730
rect 235092 239728 235139 239732
rect 235134 239672 235139 239728
rect 235022 239668 235028 239670
rect 235092 239668 235139 239672
rect 235390 239668 235396 239732
rect 235460 239730 235466 239732
rect 235533 239730 235599 239733
rect 235460 239728 235599 239730
rect 235460 239672 235538 239728
rect 235594 239672 235599 239728
rect 235460 239670 235599 239672
rect 235460 239668 235466 239670
rect 235073 239667 235139 239668
rect 235533 239667 235599 239670
rect 236085 239732 236151 239733
rect 236085 239728 236132 239732
rect 236196 239730 236202 239732
rect 236502 239730 236611 239733
rect 237230 239730 237236 239732
rect 236085 239672 236090 239728
rect 236085 239668 236132 239672
rect 236196 239670 236242 239730
rect 236502 239728 237236 239730
rect 236502 239672 236550 239728
rect 236606 239672 237236 239728
rect 236502 239670 237236 239672
rect 236196 239668 236202 239670
rect 236085 239667 236151 239668
rect 236545 239667 236611 239670
rect 237230 239668 237236 239670
rect 237300 239668 237306 239732
rect 237649 239730 237715 239733
rect 238334 239730 238340 239732
rect 237649 239728 238340 239730
rect 237649 239672 237654 239728
rect 237710 239672 238340 239728
rect 237649 239670 238340 239672
rect 237649 239667 237715 239670
rect 238334 239668 238340 239670
rect 238404 239668 238410 239732
rect 238702 239668 238708 239732
rect 238772 239730 238778 239732
rect 242934 239730 242940 239732
rect 238772 239670 242940 239730
rect 238772 239668 238778 239670
rect 242934 239668 242940 239670
rect 243004 239730 243010 239732
rect 243126 239730 243186 239837
rect 244733 239808 244738 239864
rect 244794 239808 244964 239864
rect 244733 239806 244964 239808
rect 244733 239803 244799 239806
rect 244958 239804 244964 239806
rect 245028 239804 245034 239868
rect 245142 239804 245148 239868
rect 245212 239866 245218 239868
rect 245377 239866 245443 239869
rect 245212 239864 245443 239866
rect 245212 239808 245382 239864
rect 245438 239808 245443 239864
rect 245212 239806 245443 239808
rect 245212 239804 245218 239806
rect 245377 239803 245443 239806
rect 245878 239804 245884 239868
rect 245948 239866 245954 239868
rect 246343 239866 246348 239898
rect 245948 239842 246348 239866
rect 246404 239868 246452 239898
rect 246990 239869 247050 240078
rect 249190 239940 249196 240004
rect 249260 240002 249266 240004
rect 249260 239942 249626 240002
rect 249260 239940 249266 239942
rect 246404 239842 246436 239868
rect 245948 239806 246436 239842
rect 245948 239804 245954 239806
rect 246430 239804 246436 239806
rect 246500 239804 246506 239868
rect 246987 239864 247053 239869
rect 246987 239808 246992 239864
rect 247048 239808 247053 239864
rect 246987 239803 247053 239808
rect 247539 239866 247605 239869
rect 248643 239868 248709 239869
rect 248270 239866 248276 239868
rect 247539 239864 248276 239866
rect 247539 239808 247544 239864
rect 247600 239808 248276 239864
rect 247539 239806 248276 239808
rect 247539 239803 247605 239806
rect 248270 239804 248276 239806
rect 248340 239804 248346 239868
rect 248638 239866 248644 239868
rect 248552 239806 248644 239866
rect 248638 239804 248644 239806
rect 248708 239804 248714 239868
rect 249374 239804 249380 239868
rect 249444 239804 249450 239868
rect 249566 239866 249626 239942
rect 250299 239898 250365 239903
rect 249747 239866 249813 239869
rect 249566 239864 249813 239866
rect 249566 239808 249752 239864
rect 249808 239808 249813 239864
rect 250299 239842 250304 239898
rect 250360 239866 250365 239898
rect 252599 239900 252665 239903
rect 252599 239898 252708 239900
rect 250846 239866 250852 239868
rect 250360 239842 250852 239866
rect 250299 239837 250852 239842
rect 249566 239806 249813 239808
rect 250302 239806 250852 239837
rect 248643 239803 248709 239804
rect 243004 239670 243186 239730
rect 243261 239730 243327 239733
rect 243445 239730 243511 239733
rect 243261 239728 243511 239730
rect 243261 239672 243266 239728
rect 243322 239672 243450 239728
rect 243506 239672 243511 239728
rect 243261 239670 243511 239672
rect 243004 239668 243010 239670
rect 243261 239667 243327 239670
rect 243445 239667 243511 239670
rect 244590 239668 244596 239732
rect 244660 239730 244666 239732
rect 245326 239730 245332 239732
rect 244660 239670 245332 239730
rect 244660 239668 244666 239670
rect 245326 239668 245332 239670
rect 245396 239730 245402 239732
rect 245653 239730 245719 239733
rect 245396 239728 245719 239730
rect 245396 239672 245658 239728
rect 245714 239672 245719 239728
rect 245396 239670 245719 239672
rect 245396 239668 245402 239670
rect 245653 239667 245719 239670
rect 246389 239730 246455 239733
rect 246798 239730 246804 239732
rect 246389 239728 246804 239730
rect 246389 239672 246394 239728
rect 246450 239672 246804 239728
rect 246389 239670 246804 239672
rect 246389 239667 246455 239670
rect 246798 239668 246804 239670
rect 246868 239668 246874 239732
rect 247902 239668 247908 239732
rect 247972 239730 247978 239732
rect 248137 239730 248203 239733
rect 247972 239728 248203 239730
rect 247972 239672 248142 239728
rect 248198 239672 248203 239728
rect 247972 239670 248203 239672
rect 247972 239668 247978 239670
rect 248137 239667 248203 239670
rect 248454 239668 248460 239732
rect 248524 239730 248530 239732
rect 248873 239730 248939 239733
rect 249382 239730 249442 239804
rect 249747 239803 249813 239806
rect 250846 239804 250852 239806
rect 250916 239804 250922 239868
rect 251817 239866 251883 239869
rect 251950 239866 251956 239868
rect 251817 239864 251956 239866
rect 251817 239808 251822 239864
rect 251878 239808 251956 239864
rect 251817 239806 251956 239808
rect 251817 239803 251883 239806
rect 251950 239804 251956 239806
rect 252020 239804 252026 239868
rect 252599 239842 252604 239898
rect 252660 239868 252708 239898
rect 252660 239842 252692 239868
rect 252599 239837 252692 239842
rect 252648 239806 252692 239837
rect 252686 239804 252692 239806
rect 252756 239804 252762 239868
rect 254715 239866 254781 239869
rect 254894 239866 254900 239868
rect 254715 239864 254900 239866
rect 254715 239808 254720 239864
rect 254776 239808 254900 239864
rect 254715 239806 254900 239808
rect 254715 239803 254781 239806
rect 254894 239804 254900 239806
rect 254964 239804 254970 239868
rect 248524 239728 249442 239730
rect 248524 239672 248878 239728
rect 248934 239672 249442 239728
rect 248524 239670 249442 239672
rect 249885 239730 249951 239733
rect 250110 239730 250116 239732
rect 249885 239728 250116 239730
rect 249885 239672 249890 239728
rect 249946 239672 250116 239728
rect 249885 239670 250116 239672
rect 248524 239668 248530 239670
rect 248873 239667 248939 239670
rect 249885 239667 249951 239670
rect 250110 239668 250116 239670
rect 250180 239668 250186 239732
rect 250989 239730 251055 239733
rect 251449 239730 251515 239733
rect 250989 239728 251515 239730
rect 250989 239672 250994 239728
rect 251050 239672 251454 239728
rect 251510 239672 251515 239728
rect 250989 239670 251515 239672
rect 250989 239667 251055 239670
rect 251449 239667 251515 239670
rect 251766 239668 251772 239732
rect 251836 239730 251842 239732
rect 251909 239730 251975 239733
rect 251836 239728 251975 239730
rect 251836 239672 251914 239728
rect 251970 239672 251975 239728
rect 251836 239670 251975 239672
rect 251836 239668 251842 239670
rect 251909 239667 251975 239670
rect 252737 239730 252803 239733
rect 253422 239730 253428 239732
rect 252737 239728 253428 239730
rect 252737 239672 252742 239728
rect 252798 239672 253428 239728
rect 252737 239670 253428 239672
rect 252737 239667 252803 239670
rect 253422 239668 253428 239670
rect 253492 239668 253498 239732
rect 255129 239730 255195 239733
rect 255270 239730 255330 240214
rect 258390 240212 258396 240276
rect 258460 240274 258466 240276
rect 267733 240274 267799 240277
rect 258460 240272 267799 240274
rect 258460 240216 267738 240272
rect 267794 240216 267799 240272
rect 258460 240214 267799 240216
rect 258460 240212 258466 240214
rect 267733 240211 267799 240214
rect 269481 240274 269547 240277
rect 277485 240274 277551 240277
rect 277853 240274 277919 240277
rect 269481 240272 277919 240274
rect 269481 240216 269486 240272
rect 269542 240216 277490 240272
rect 277546 240216 277858 240272
rect 277914 240216 277919 240272
rect 269481 240214 277919 240216
rect 269481 240211 269547 240214
rect 277485 240211 277551 240214
rect 277853 240211 277919 240214
rect 267917 240138 267983 240141
rect 259502 240136 267983 240138
rect 259502 240080 267922 240136
rect 267978 240080 267983 240136
rect 259502 240078 267983 240080
rect 258390 240002 258396 240004
rect 257846 239942 258396 240002
rect 256095 239900 256161 239903
rect 256052 239898 256161 239900
rect 256052 239868 256100 239898
rect 255998 239804 256004 239868
rect 256068 239842 256100 239868
rect 256156 239842 256161 239898
rect 256068 239837 256161 239842
rect 256068 239806 256112 239837
rect 256068 239804 256074 239806
rect 255129 239728 255330 239730
rect 255129 239672 255134 239728
rect 255190 239672 255330 239728
rect 255129 239670 255330 239672
rect 255129 239667 255195 239670
rect 255446 239668 255452 239732
rect 255516 239730 255522 239732
rect 256049 239730 256115 239733
rect 257153 239732 257219 239733
rect 255516 239728 256115 239730
rect 255516 239672 256054 239728
rect 256110 239672 256115 239728
rect 255516 239670 256115 239672
rect 255516 239668 255522 239670
rect 256049 239667 256115 239670
rect 257102 239668 257108 239732
rect 257172 239730 257219 239732
rect 257846 239730 257906 239942
rect 258390 239940 258396 239942
rect 258460 239940 258466 240004
rect 258119 239866 258185 239869
rect 259502 239866 259562 240078
rect 267917 240075 267983 240078
rect 268009 240002 268075 240005
rect 260790 240000 268075 240002
rect 260790 239944 268014 240000
rect 268070 239944 268075 240000
rect 260790 239942 268075 239944
rect 260790 239869 260850 239942
rect 268009 239939 268075 239942
rect 258119 239864 259562 239866
rect 258119 239808 258124 239864
rect 258180 239808 259562 239864
rect 258119 239806 259562 239808
rect 260511 239866 260577 239869
rect 260511 239864 260620 239866
rect 260511 239808 260516 239864
rect 260572 239808 260620 239864
rect 258119 239803 258185 239806
rect 260511 239803 260620 239808
rect 260787 239864 260853 239869
rect 260787 239808 260792 239864
rect 260848 239808 260853 239864
rect 260787 239803 260853 239808
rect 261431 239866 261497 239869
rect 261702 239866 261708 239868
rect 261431 239864 261708 239866
rect 261431 239808 261436 239864
rect 261492 239808 261708 239864
rect 261431 239806 261708 239808
rect 261431 239803 261497 239806
rect 261702 239804 261708 239806
rect 261772 239804 261778 239868
rect 262438 239804 262444 239868
rect 262508 239866 262514 239868
rect 262627 239866 262693 239869
rect 262508 239864 262693 239866
rect 262508 239808 262632 239864
rect 262688 239808 262693 239864
rect 262508 239806 262693 239808
rect 262508 239804 262514 239806
rect 262627 239803 262693 239806
rect 262990 239804 262996 239868
rect 263060 239866 263066 239868
rect 263179 239866 263245 239869
rect 263060 239864 263245 239866
rect 263060 239808 263184 239864
rect 263240 239808 263245 239864
rect 263060 239806 263245 239808
rect 263060 239804 263066 239806
rect 263179 239803 263245 239806
rect 263542 239804 263548 239868
rect 263612 239866 263618 239868
rect 263910 239866 263916 239868
rect 263612 239806 263916 239866
rect 263612 239804 263618 239806
rect 263910 239804 263916 239806
rect 263980 239866 263986 239868
rect 264099 239866 264165 239869
rect 263980 239864 264165 239866
rect 263980 239808 264104 239864
rect 264160 239808 264165 239864
rect 263980 239806 264165 239808
rect 263980 239804 263986 239806
rect 264099 239803 264165 239806
rect 264651 239866 264717 239869
rect 265387 239868 265453 239869
rect 264830 239866 264836 239868
rect 264651 239864 264836 239866
rect 264651 239808 264656 239864
rect 264712 239808 264836 239864
rect 264651 239806 264836 239808
rect 264651 239803 264717 239806
rect 264830 239804 264836 239806
rect 264900 239804 264906 239868
rect 265382 239866 265388 239868
rect 265296 239806 265388 239866
rect 265382 239804 265388 239806
rect 265452 239804 265458 239868
rect 266031 239866 266097 239869
rect 266302 239866 266308 239868
rect 266031 239864 266308 239866
rect 266031 239808 266036 239864
rect 266092 239808 266308 239864
rect 266031 239806 266308 239808
rect 265387 239803 265453 239804
rect 266031 239803 266097 239806
rect 266302 239804 266308 239806
rect 266372 239804 266378 239868
rect 258533 239730 258599 239733
rect 259453 239732 259519 239733
rect 259453 239730 259500 239732
rect 257172 239728 257264 239730
rect 257214 239672 257264 239728
rect 257172 239670 257264 239672
rect 257846 239728 258599 239730
rect 257846 239672 258538 239728
rect 258594 239672 258599 239728
rect 257846 239670 258599 239672
rect 259408 239728 259500 239730
rect 259408 239672 259458 239728
rect 259408 239670 259500 239672
rect 257172 239668 257219 239670
rect 257153 239667 257219 239668
rect 258533 239667 258599 239670
rect 259453 239668 259500 239670
rect 259564 239668 259570 239732
rect 259678 239668 259684 239732
rect 259748 239730 259754 239732
rect 260414 239730 260420 239732
rect 259748 239670 260420 239730
rect 259748 239668 259754 239670
rect 260414 239668 260420 239670
rect 260484 239730 260490 239732
rect 260560 239730 260620 239803
rect 260484 239670 260620 239730
rect 261385 239730 261451 239733
rect 261518 239730 261524 239732
rect 261385 239728 261524 239730
rect 261385 239672 261390 239728
rect 261446 239672 261524 239728
rect 261385 239670 261524 239672
rect 260484 239668 260490 239670
rect 259453 239667 259519 239668
rect 261385 239667 261451 239670
rect 261518 239668 261524 239670
rect 261588 239668 261594 239732
rect 261661 239730 261727 239733
rect 262070 239730 262076 239732
rect 261661 239728 262076 239730
rect 261661 239672 261666 239728
rect 261722 239672 262076 239728
rect 261661 239670 262076 239672
rect 261661 239667 261727 239670
rect 262070 239668 262076 239670
rect 262140 239668 262146 239732
rect 262254 239668 262260 239732
rect 262324 239730 262330 239732
rect 263358 239730 263364 239732
rect 262324 239670 263364 239730
rect 262324 239668 262330 239670
rect 263358 239668 263364 239670
rect 263428 239730 263434 239732
rect 263593 239730 263659 239733
rect 263428 239728 263659 239730
rect 263428 239672 263598 239728
rect 263654 239672 263659 239728
rect 263428 239670 263659 239672
rect 263428 239668 263434 239670
rect 263593 239667 263659 239670
rect 264094 239668 264100 239732
rect 264164 239730 264170 239732
rect 264654 239730 264714 239803
rect 264164 239670 264714 239730
rect 264881 239730 264947 239733
rect 265198 239730 265204 239732
rect 264881 239728 265204 239730
rect 264881 239672 264886 239728
rect 264942 239672 265204 239728
rect 264881 239670 265204 239672
rect 264164 239668 264170 239670
rect 264881 239667 264947 239670
rect 265198 239668 265204 239670
rect 265268 239668 265274 239732
rect 265525 239730 265591 239733
rect 265750 239730 265756 239732
rect 265525 239728 265756 239730
rect 265525 239672 265530 239728
rect 265586 239672 265756 239728
rect 265525 239670 265756 239672
rect 265525 239667 265591 239670
rect 265750 239668 265756 239670
rect 265820 239668 265826 239732
rect 266118 239668 266124 239732
rect 266188 239730 266194 239732
rect 266307 239730 266373 239733
rect 266188 239728 266373 239730
rect 266188 239672 266312 239728
rect 266368 239672 266373 239728
rect 266188 239670 266373 239672
rect 266188 239668 266194 239670
rect 266307 239667 266373 239670
rect 266670 239668 266676 239732
rect 266740 239730 266746 239732
rect 266813 239730 266879 239733
rect 266740 239728 266879 239730
rect 266740 239672 266818 239728
rect 266874 239672 266879 239728
rect 266740 239670 266879 239672
rect 266740 239668 266746 239670
rect 266813 239667 266879 239670
rect 285121 239594 285187 239597
rect 234570 239592 285187 239594
rect 234570 239536 285126 239592
rect 285182 239536 285187 239592
rect 234570 239534 285187 239536
rect 233068 239532 233074 239534
rect 233325 239531 233391 239534
rect 285121 239531 285187 239534
rect 227916 239398 228052 239458
rect 227916 239396 227922 239398
rect 228214 239396 228220 239460
rect 228284 239458 228290 239460
rect 228817 239458 228883 239461
rect 228284 239456 228883 239458
rect 228284 239400 228822 239456
rect 228878 239400 228883 239456
rect 228284 239398 228883 239400
rect 228284 239396 228290 239398
rect 227437 239395 227503 239396
rect 228817 239395 228883 239398
rect 229318 239396 229324 239460
rect 229388 239458 229394 239460
rect 230013 239458 230079 239461
rect 229388 239456 230079 239458
rect 229388 239400 230018 239456
rect 230074 239400 230079 239456
rect 229388 239398 230079 239400
rect 229388 239396 229394 239398
rect 230013 239395 230079 239398
rect 230289 239458 230355 239461
rect 230422 239458 230428 239460
rect 230289 239456 230428 239458
rect 230289 239400 230294 239456
rect 230350 239400 230428 239456
rect 230289 239398 230428 239400
rect 230289 239395 230355 239398
rect 230422 239396 230428 239398
rect 230492 239396 230498 239460
rect 233233 239458 233299 239461
rect 233785 239458 233851 239461
rect 233233 239456 233851 239458
rect 233233 239400 233238 239456
rect 233294 239400 233790 239456
rect 233846 239400 233851 239456
rect 233233 239398 233851 239400
rect 233233 239395 233299 239398
rect 233785 239395 233851 239398
rect 233969 239458 234035 239461
rect 234286 239458 234292 239460
rect 233969 239456 234292 239458
rect 233969 239400 233974 239456
rect 234030 239400 234292 239456
rect 233969 239398 234292 239400
rect 233969 239395 234035 239398
rect 234286 239396 234292 239398
rect 234356 239458 234362 239460
rect 234889 239458 234955 239461
rect 234356 239456 234955 239458
rect 234356 239400 234894 239456
rect 234950 239400 234955 239456
rect 234356 239398 234955 239400
rect 234356 239396 234362 239398
rect 234889 239395 234955 239398
rect 235206 239396 235212 239460
rect 235276 239458 235282 239460
rect 235901 239458 235967 239461
rect 235276 239456 235967 239458
rect 235276 239400 235906 239456
rect 235962 239400 235967 239456
rect 235276 239398 235967 239400
rect 235276 239396 235282 239398
rect 235901 239395 235967 239398
rect 236177 239458 236243 239461
rect 237005 239460 237071 239461
rect 236310 239458 236316 239460
rect 236177 239456 236316 239458
rect 236177 239400 236182 239456
rect 236238 239400 236316 239456
rect 236177 239398 236316 239400
rect 236177 239395 236243 239398
rect 236310 239396 236316 239398
rect 236380 239396 236386 239460
rect 237005 239458 237052 239460
rect 236960 239456 237052 239458
rect 236960 239400 237010 239456
rect 236960 239398 237052 239400
rect 237005 239396 237052 239398
rect 237116 239396 237122 239460
rect 238150 239396 238156 239460
rect 238220 239458 238226 239460
rect 238293 239458 238359 239461
rect 238220 239456 238359 239458
rect 238220 239400 238298 239456
rect 238354 239400 238359 239456
rect 238220 239398 238359 239400
rect 238220 239396 238226 239398
rect 237005 239395 237071 239396
rect 238293 239395 238359 239398
rect 238518 239396 238524 239460
rect 238588 239458 238594 239460
rect 238661 239458 238727 239461
rect 238937 239460 239003 239461
rect 239305 239460 239371 239461
rect 238588 239456 238727 239458
rect 238588 239400 238666 239456
rect 238722 239400 238727 239456
rect 238588 239398 238727 239400
rect 238588 239396 238594 239398
rect 238661 239395 238727 239398
rect 238886 239396 238892 239460
rect 238956 239458 239003 239460
rect 238956 239456 239048 239458
rect 238998 239400 239048 239456
rect 238956 239398 239048 239400
rect 238956 239396 239003 239398
rect 239254 239396 239260 239460
rect 239324 239458 239371 239460
rect 239324 239456 239416 239458
rect 239366 239400 239416 239456
rect 239324 239398 239416 239400
rect 239324 239396 239371 239398
rect 239806 239396 239812 239460
rect 239876 239458 239882 239460
rect 242893 239458 242959 239461
rect 239876 239456 242959 239458
rect 239876 239400 242898 239456
rect 242954 239400 242959 239456
rect 239876 239398 242959 239400
rect 239876 239396 239882 239398
rect 238937 239395 239003 239396
rect 239305 239395 239371 239396
rect 242893 239395 242959 239398
rect 243118 239396 243124 239460
rect 243188 239458 243194 239460
rect 243261 239458 243327 239461
rect 243188 239456 243327 239458
rect 243188 239400 243266 239456
rect 243322 239400 243327 239456
rect 243188 239398 243327 239400
rect 243188 239396 243194 239398
rect 243261 239395 243327 239398
rect 244457 239458 244523 239461
rect 244774 239458 244780 239460
rect 244457 239456 244780 239458
rect 244457 239400 244462 239456
rect 244518 239400 244780 239456
rect 244457 239398 244780 239400
rect 244457 239395 244523 239398
rect 244774 239396 244780 239398
rect 244844 239458 244850 239460
rect 245285 239458 245351 239461
rect 244844 239456 245351 239458
rect 244844 239400 245290 239456
rect 245346 239400 245351 239456
rect 244844 239398 245351 239400
rect 244844 239396 244850 239398
rect 245285 239395 245351 239398
rect 247309 239458 247375 239461
rect 247534 239458 247540 239460
rect 247309 239456 247540 239458
rect 247309 239400 247314 239456
rect 247370 239400 247540 239456
rect 247309 239398 247540 239400
rect 247309 239395 247375 239398
rect 247534 239396 247540 239398
rect 247604 239396 247610 239460
rect 247861 239458 247927 239461
rect 249517 239460 249583 239461
rect 248086 239458 248092 239460
rect 247861 239456 248092 239458
rect 247861 239400 247866 239456
rect 247922 239400 248092 239456
rect 247861 239398 248092 239400
rect 247861 239395 247927 239398
rect 248086 239396 248092 239398
rect 248156 239396 248162 239460
rect 249517 239458 249564 239460
rect 249472 239456 249564 239458
rect 249472 239400 249522 239456
rect 249472 239398 249564 239400
rect 249517 239396 249564 239398
rect 249628 239396 249634 239460
rect 252318 239396 252324 239460
rect 252388 239458 252394 239460
rect 252553 239458 252619 239461
rect 253013 239460 253079 239461
rect 253013 239458 253060 239460
rect 252388 239456 252619 239458
rect 252388 239400 252558 239456
rect 252614 239400 252619 239456
rect 252388 239398 252619 239400
rect 252968 239456 253060 239458
rect 252968 239400 253018 239456
rect 252968 239398 253060 239400
rect 252388 239396 252394 239398
rect 249517 239395 249583 239396
rect 252553 239395 252619 239398
rect 253013 239396 253060 239398
rect 253124 239396 253130 239460
rect 253238 239396 253244 239460
rect 253308 239458 253314 239460
rect 253841 239458 253907 239461
rect 253308 239456 253907 239458
rect 253308 239400 253846 239456
rect 253902 239400 253907 239456
rect 253308 239398 253907 239400
rect 253308 239396 253314 239398
rect 253013 239395 253079 239396
rect 253841 239395 253907 239398
rect 255957 239458 256023 239461
rect 256366 239458 256372 239460
rect 255957 239456 256372 239458
rect 255957 239400 255962 239456
rect 256018 239400 256372 239456
rect 255957 239398 256372 239400
rect 255957 239395 256023 239398
rect 256366 239396 256372 239398
rect 256436 239396 256442 239460
rect 257286 239396 257292 239460
rect 257356 239458 257362 239460
rect 257613 239458 257679 239461
rect 257356 239456 257679 239458
rect 257356 239400 257618 239456
rect 257674 239400 257679 239456
rect 257356 239398 257679 239400
rect 257356 239396 257362 239398
rect 257613 239395 257679 239398
rect 258073 239458 258139 239461
rect 258574 239458 258580 239460
rect 258073 239456 258580 239458
rect 258073 239400 258078 239456
rect 258134 239400 258580 239456
rect 258073 239398 258580 239400
rect 258073 239395 258139 239398
rect 258574 239396 258580 239398
rect 258644 239396 258650 239460
rect 258809 239458 258875 239461
rect 259126 239458 259132 239460
rect 258809 239456 259132 239458
rect 258809 239400 258814 239456
rect 258870 239400 259132 239456
rect 258809 239398 259132 239400
rect 258809 239395 258875 239398
rect 259126 239396 259132 239398
rect 259196 239396 259202 239460
rect 259310 239396 259316 239460
rect 259380 239458 259386 239460
rect 259729 239458 259795 239461
rect 259380 239456 259795 239458
rect 259380 239400 259734 239456
rect 259790 239400 259795 239456
rect 259380 239398 259795 239400
rect 259380 239396 259386 239398
rect 259729 239395 259795 239398
rect 260465 239458 260531 239461
rect 260649 239458 260715 239461
rect 260465 239456 260715 239458
rect 260465 239400 260470 239456
rect 260526 239400 260654 239456
rect 260710 239400 260715 239456
rect 260465 239398 260715 239400
rect 260465 239395 260531 239398
rect 260649 239395 260715 239398
rect 261150 239396 261156 239460
rect 261220 239458 261226 239460
rect 261937 239458 262003 239461
rect 261220 239456 262003 239458
rect 261220 239400 261942 239456
rect 261998 239400 262003 239456
rect 261220 239398 262003 239400
rect 261220 239396 261226 239398
rect 261937 239395 262003 239398
rect 262397 239458 262463 239461
rect 263358 239458 263364 239460
rect 262397 239456 263364 239458
rect 262397 239400 262402 239456
rect 262458 239400 263364 239456
rect 262397 239398 263364 239400
rect 262397 239395 262463 239398
rect 263358 239396 263364 239398
rect 263428 239396 263434 239460
rect 263726 239396 263732 239460
rect 263796 239458 263802 239460
rect 264697 239458 264763 239461
rect 263796 239456 264763 239458
rect 263796 239400 264702 239456
rect 264758 239400 264763 239456
rect 263796 239398 264763 239400
rect 263796 239396 263802 239398
rect 264697 239395 264763 239398
rect 264881 239458 264947 239461
rect 289169 239458 289235 239461
rect 264881 239456 289235 239458
rect 264881 239400 264886 239456
rect 264942 239400 289174 239456
rect 289230 239400 289235 239456
rect 264881 239398 289235 239400
rect 264881 239395 264947 239398
rect 289169 239395 289235 239398
rect 228173 239322 228239 239325
rect 270217 239322 270283 239325
rect 226198 239320 270283 239322
rect 226198 239264 228178 239320
rect 228234 239264 270222 239320
rect 270278 239264 270283 239320
rect 226198 239262 270283 239264
rect 228173 239259 228239 239262
rect 270217 239259 270283 239262
rect 211705 239186 211771 239189
rect 255681 239186 255747 239189
rect 303153 239186 303219 239189
rect 211705 239184 303219 239186
rect 211705 239128 211710 239184
rect 211766 239128 255686 239184
rect 255742 239128 303158 239184
rect 303214 239128 303219 239184
rect 211705 239126 303219 239128
rect 211705 239123 211771 239126
rect 255681 239123 255747 239126
rect 303153 239123 303219 239126
rect 219893 239050 219959 239053
rect 223798 239050 223804 239052
rect 219893 239048 223804 239050
rect 219893 238992 219898 239048
rect 219954 238992 223804 239048
rect 219893 238990 223804 238992
rect 219893 238987 219959 238990
rect 223798 238988 223804 238990
rect 223868 238988 223874 239052
rect 225454 238988 225460 239052
rect 225524 239050 225530 239052
rect 226609 239050 226675 239053
rect 225524 239048 226675 239050
rect 225524 238992 226614 239048
rect 226670 238992 226675 239048
rect 225524 238990 226675 238992
rect 225524 238988 225530 238990
rect 226609 238987 226675 238990
rect 226977 239050 227043 239053
rect 282453 239050 282519 239053
rect 226977 239048 282519 239050
rect 226977 238992 226982 239048
rect 227038 238992 282458 239048
rect 282514 238992 282519 239048
rect 226977 238990 282519 238992
rect 226977 238987 227043 238990
rect 282453 238987 282519 238990
rect 220629 238914 220695 238917
rect 223113 238914 223179 238917
rect 220629 238912 223179 238914
rect 220629 238856 220634 238912
rect 220690 238856 223118 238912
rect 223174 238856 223179 238912
rect 220629 238854 223179 238856
rect 220629 238851 220695 238854
rect 223113 238851 223179 238854
rect 223757 238914 223823 238917
rect 282913 238914 282979 238917
rect 223757 238912 282979 238914
rect 223757 238856 223762 238912
rect 223818 238856 282918 238912
rect 282974 238856 282979 238912
rect 223757 238854 282979 238856
rect 223757 238851 223823 238854
rect 282913 238851 282979 238854
rect 217501 238778 217567 238781
rect 227989 238778 228055 238781
rect 228398 238778 228404 238780
rect 217501 238776 224970 238778
rect 217501 238720 217506 238776
rect 217562 238720 224970 238776
rect 217501 238718 224970 238720
rect 217501 238715 217567 238718
rect 224910 238642 224970 238718
rect 227989 238776 228404 238778
rect 227989 238720 227994 238776
rect 228050 238720 228404 238776
rect 227989 238718 228404 238720
rect 227989 238715 228055 238718
rect 228398 238716 228404 238718
rect 228468 238778 228474 238780
rect 229185 238778 229251 238781
rect 228468 238776 229251 238778
rect 228468 238720 229190 238776
rect 229246 238720 229251 238776
rect 228468 238718 229251 238720
rect 228468 238716 228474 238718
rect 229185 238715 229251 238718
rect 231117 238780 231183 238781
rect 231117 238776 231164 238780
rect 231228 238778 231234 238780
rect 232037 238778 232103 238781
rect 232446 238778 232452 238780
rect 231117 238720 231122 238776
rect 231117 238716 231164 238720
rect 231228 238718 231274 238778
rect 232037 238776 232452 238778
rect 232037 238720 232042 238776
rect 232098 238720 232452 238776
rect 232037 238718 232452 238720
rect 231228 238716 231234 238718
rect 231117 238715 231183 238716
rect 232037 238715 232103 238718
rect 232446 238716 232452 238718
rect 232516 238716 232522 238780
rect 233233 238778 233299 238781
rect 233734 238778 233740 238780
rect 233233 238776 233740 238778
rect 233233 238720 233238 238776
rect 233294 238720 233740 238776
rect 233233 238718 233740 238720
rect 233233 238715 233299 238718
rect 233734 238716 233740 238718
rect 233804 238716 233810 238780
rect 235441 238778 235507 238781
rect 235574 238778 235580 238780
rect 235441 238776 235580 238778
rect 235441 238720 235446 238776
rect 235502 238720 235580 238776
rect 235441 238718 235580 238720
rect 235441 238715 235507 238718
rect 235574 238716 235580 238718
rect 235644 238716 235650 238780
rect 236453 238778 236519 238781
rect 236729 238778 236795 238781
rect 236453 238776 236795 238778
rect 236453 238720 236458 238776
rect 236514 238720 236734 238776
rect 236790 238720 236795 238776
rect 236453 238718 236795 238720
rect 236453 238715 236519 238718
rect 236729 238715 236795 238718
rect 239438 238716 239444 238780
rect 239508 238778 239514 238780
rect 240133 238778 240199 238781
rect 239508 238776 240199 238778
rect 239508 238720 240138 238776
rect 240194 238720 240199 238776
rect 239508 238718 240199 238720
rect 239508 238716 239514 238718
rect 240133 238715 240199 238718
rect 240685 238778 240751 238781
rect 240910 238778 240916 238780
rect 240685 238776 240916 238778
rect 240685 238720 240690 238776
rect 240746 238720 240916 238776
rect 240685 238718 240916 238720
rect 240685 238715 240751 238718
rect 240910 238716 240916 238718
rect 240980 238716 240986 238780
rect 245694 238778 245700 238780
rect 244230 238718 245700 238778
rect 232773 238642 232839 238645
rect 224910 238640 232839 238642
rect 224910 238584 232778 238640
rect 232834 238584 232839 238640
rect 224910 238582 232839 238584
rect 232773 238579 232839 238582
rect 233601 238642 233667 238645
rect 233918 238642 233924 238644
rect 233601 238640 233924 238642
rect 233601 238584 233606 238640
rect 233662 238584 233924 238640
rect 233601 238582 233924 238584
rect 233601 238579 233667 238582
rect 233918 238580 233924 238582
rect 233988 238580 233994 238644
rect 234153 238642 234219 238645
rect 240317 238642 240383 238645
rect 241145 238644 241211 238645
rect 234153 238640 240383 238642
rect 234153 238584 234158 238640
rect 234214 238584 240322 238640
rect 240378 238584 240383 238640
rect 234153 238582 240383 238584
rect 234153 238579 234219 238582
rect 240317 238579 240383 238582
rect 241094 238580 241100 238644
rect 241164 238642 241211 238644
rect 241421 238642 241487 238645
rect 244230 238642 244290 238718
rect 245694 238716 245700 238718
rect 245764 238716 245770 238780
rect 249926 238716 249932 238780
rect 249996 238778 250002 238780
rect 250989 238778 251055 238781
rect 249996 238776 251055 238778
rect 249996 238720 250994 238776
rect 251050 238720 251055 238776
rect 249996 238718 251055 238720
rect 249996 238716 250002 238718
rect 250989 238715 251055 238718
rect 255865 238778 255931 238781
rect 255865 238776 256802 238778
rect 255865 238720 255870 238776
rect 255926 238720 256802 238776
rect 255865 238718 256802 238720
rect 255865 238715 255931 238718
rect 245377 238644 245443 238645
rect 241164 238640 241256 238642
rect 241206 238584 241256 238640
rect 241164 238582 241256 238584
rect 241421 238640 244290 238642
rect 241421 238584 241426 238640
rect 241482 238584 244290 238640
rect 241421 238582 244290 238584
rect 241164 238580 241211 238582
rect 241145 238579 241211 238580
rect 241421 238579 241487 238582
rect 245326 238580 245332 238644
rect 245396 238642 245443 238644
rect 245396 238640 245488 238642
rect 245438 238584 245488 238640
rect 245396 238582 245488 238584
rect 245396 238580 245443 238582
rect 250294 238580 250300 238644
rect 250364 238642 250370 238644
rect 250713 238642 250779 238645
rect 250364 238640 250779 238642
rect 250364 238584 250718 238640
rect 250774 238584 250779 238640
rect 250364 238582 250779 238584
rect 250364 238580 250370 238582
rect 245377 238579 245443 238580
rect 250713 238579 250779 238582
rect 255129 238642 255195 238645
rect 255630 238642 255636 238644
rect 255129 238640 255636 238642
rect 255129 238584 255134 238640
rect 255190 238584 255636 238640
rect 255129 238582 255636 238584
rect 255129 238579 255195 238582
rect 255630 238580 255636 238582
rect 255700 238580 255706 238644
rect 256742 238642 256802 238718
rect 256918 238716 256924 238780
rect 256988 238778 256994 238780
rect 257245 238778 257311 238781
rect 256988 238776 257311 238778
rect 256988 238720 257250 238776
rect 257306 238720 257311 238776
rect 256988 238718 257311 238720
rect 256988 238716 256994 238718
rect 257245 238715 257311 238718
rect 259085 238778 259151 238781
rect 260373 238780 260439 238781
rect 259494 238778 259500 238780
rect 259085 238776 259500 238778
rect 259085 238720 259090 238776
rect 259146 238720 259500 238776
rect 259085 238718 259500 238720
rect 259085 238715 259151 238718
rect 259494 238716 259500 238718
rect 259564 238716 259570 238780
rect 260373 238776 260420 238780
rect 260484 238778 260490 238780
rect 260373 238720 260378 238776
rect 260373 238716 260420 238720
rect 260484 238718 260530 238778
rect 260484 238716 260490 238718
rect 260598 238716 260604 238780
rect 260668 238778 260674 238780
rect 262581 238778 262647 238781
rect 264145 238780 264211 238781
rect 260668 238776 262647 238778
rect 260668 238720 262586 238776
rect 262642 238720 262647 238776
rect 260668 238718 262647 238720
rect 260668 238716 260674 238718
rect 260373 238715 260439 238716
rect 262581 238715 262647 238718
rect 264094 238716 264100 238780
rect 264164 238778 264211 238780
rect 265157 238778 265223 238781
rect 265382 238778 265388 238780
rect 264164 238776 264256 238778
rect 264206 238720 264256 238776
rect 264164 238718 264256 238720
rect 265157 238776 265388 238778
rect 265157 238720 265162 238776
rect 265218 238720 265388 238776
rect 265157 238718 265388 238720
rect 264164 238716 264211 238718
rect 264145 238715 264211 238716
rect 265157 238715 265223 238718
rect 265382 238716 265388 238718
rect 265452 238716 265458 238780
rect 266169 238778 266235 238781
rect 268653 238778 268719 238781
rect 271822 238778 271828 238780
rect 266169 238776 271828 238778
rect 266169 238720 266174 238776
rect 266230 238720 268658 238776
rect 268714 238720 271828 238776
rect 266169 238718 271828 238720
rect 266169 238715 266235 238718
rect 268653 238715 268719 238718
rect 271822 238716 271828 238718
rect 271892 238716 271898 238780
rect 260373 238642 260439 238645
rect 256742 238640 260439 238642
rect 256742 238584 260378 238640
rect 260434 238584 260439 238640
rect 256742 238582 260439 238584
rect 260373 238579 260439 238582
rect 260649 238642 260715 238645
rect 261017 238642 261083 238645
rect 260649 238640 261083 238642
rect 260649 238584 260654 238640
rect 260710 238584 261022 238640
rect 261078 238584 261083 238640
rect 260649 238582 261083 238584
rect 260649 238579 260715 238582
rect 261017 238579 261083 238582
rect 261293 238642 261359 238645
rect 270585 238642 270651 238645
rect 261293 238640 270651 238642
rect 261293 238584 261298 238640
rect 261354 238584 270590 238640
rect 270646 238584 270651 238640
rect 261293 238582 270651 238584
rect 261293 238579 261359 238582
rect 270585 238579 270651 238582
rect 204897 238506 204963 238509
rect 223665 238506 223731 238509
rect 204897 238504 223731 238506
rect 204897 238448 204902 238504
rect 204958 238448 223670 238504
rect 223726 238448 223731 238504
rect 204897 238446 223731 238448
rect 204897 238443 204963 238446
rect 223665 238443 223731 238446
rect 234286 238444 234292 238508
rect 234356 238506 234362 238508
rect 259310 238506 259316 238508
rect 234356 238446 259316 238506
rect 234356 238444 234362 238446
rect 259310 238444 259316 238446
rect 259380 238444 259386 238508
rect 259637 238506 259703 238509
rect 271045 238506 271111 238509
rect 259637 238504 271111 238506
rect 259637 238448 259642 238504
rect 259698 238448 271050 238504
rect 271106 238448 271111 238504
rect 259637 238446 271111 238448
rect 186814 238308 186820 238372
rect 186884 238370 186890 238372
rect 212073 238370 212139 238373
rect 229369 238370 229435 238373
rect 186884 238368 229435 238370
rect 186884 238312 212078 238368
rect 212134 238312 229374 238368
rect 229430 238312 229435 238368
rect 186884 238310 229435 238312
rect 186884 238308 186890 238310
rect 212073 238307 212139 238310
rect 229369 238307 229435 238310
rect 229737 238370 229803 238373
rect 258257 238370 258323 238373
rect 258390 238370 258396 238372
rect 229737 238368 255514 238370
rect 229737 238312 229742 238368
rect 229798 238312 255514 238368
rect 229737 238310 255514 238312
rect 229737 238307 229803 238310
rect 175958 238172 175964 238236
rect 176028 238234 176034 238236
rect 206645 238234 206711 238237
rect 176028 238232 206711 238234
rect 176028 238176 206650 238232
rect 206706 238176 206711 238232
rect 176028 238174 206711 238176
rect 176028 238172 176034 238174
rect 206645 238171 206711 238174
rect 208945 238234 209011 238237
rect 223481 238234 223547 238237
rect 208945 238232 223547 238234
rect 208945 238176 208950 238232
rect 209006 238176 223486 238232
rect 223542 238176 223547 238232
rect 208945 238174 223547 238176
rect 208945 238171 209011 238174
rect 223481 238171 223547 238174
rect 223665 238234 223731 238237
rect 223982 238234 223988 238236
rect 223665 238232 223988 238234
rect 223665 238176 223670 238232
rect 223726 238176 223988 238232
rect 223665 238174 223988 238176
rect 223665 238171 223731 238174
rect 223982 238172 223988 238174
rect 224052 238172 224058 238236
rect 226609 238234 226675 238237
rect 227294 238234 227300 238236
rect 226609 238232 227300 238234
rect 226609 238176 226614 238232
rect 226670 238176 227300 238232
rect 226609 238174 227300 238176
rect 226609 238171 226675 238174
rect 227294 238172 227300 238174
rect 227364 238172 227370 238236
rect 231117 238234 231183 238237
rect 231710 238234 231716 238236
rect 231117 238232 231716 238234
rect 231117 238176 231122 238232
rect 231178 238176 231716 238232
rect 231117 238174 231716 238176
rect 231117 238171 231183 238174
rect 231710 238172 231716 238174
rect 231780 238172 231786 238236
rect 233550 238172 233556 238236
rect 233620 238234 233626 238236
rect 234521 238234 234587 238237
rect 233620 238232 234587 238234
rect 233620 238176 234526 238232
rect 234582 238176 234587 238232
rect 233620 238174 234587 238176
rect 233620 238172 233626 238174
rect 234521 238171 234587 238174
rect 236126 238172 236132 238236
rect 236196 238234 236202 238236
rect 236453 238234 236519 238237
rect 236196 238232 236519 238234
rect 236196 238176 236458 238232
rect 236514 238176 236519 238232
rect 236196 238174 236519 238176
rect 236196 238172 236202 238174
rect 236453 238171 236519 238174
rect 236678 238172 236684 238236
rect 236748 238234 236754 238236
rect 236913 238234 236979 238237
rect 236748 238232 236979 238234
rect 236748 238176 236918 238232
rect 236974 238176 236979 238232
rect 236748 238174 236979 238176
rect 236748 238172 236754 238174
rect 236913 238171 236979 238174
rect 238845 238234 238911 238237
rect 239254 238234 239260 238236
rect 238845 238232 239260 238234
rect 238845 238176 238850 238232
rect 238906 238176 239260 238232
rect 238845 238174 239260 238176
rect 238845 238171 238911 238174
rect 239254 238172 239260 238174
rect 239324 238172 239330 238236
rect 240869 238234 240935 238237
rect 241278 238234 241284 238236
rect 240869 238232 241284 238234
rect 240869 238176 240874 238232
rect 240930 238176 241284 238232
rect 240869 238174 241284 238176
rect 240869 238171 240935 238174
rect 241278 238172 241284 238174
rect 241348 238172 241354 238236
rect 242382 238172 242388 238236
rect 242452 238234 242458 238236
rect 244733 238234 244799 238237
rect 242452 238232 244799 238234
rect 242452 238176 244738 238232
rect 244794 238176 244799 238232
rect 242452 238174 244799 238176
rect 255454 238234 255514 238310
rect 258257 238368 258396 238370
rect 258257 238312 258262 238368
rect 258318 238312 258396 238368
rect 258257 238310 258396 238312
rect 258257 238307 258323 238310
rect 258390 238308 258396 238310
rect 258460 238308 258466 238372
rect 258942 238234 258948 238236
rect 255454 238174 258948 238234
rect 242452 238172 242458 238174
rect 244733 238171 244799 238174
rect 258942 238172 258948 238174
rect 259012 238172 259018 238236
rect 259318 238234 259378 238444
rect 259637 238443 259703 238446
rect 271045 238443 271111 238446
rect 259729 238370 259795 238373
rect 259862 238370 259868 238372
rect 259729 238368 259868 238370
rect 259729 238312 259734 238368
rect 259790 238312 259868 238368
rect 259729 238310 259868 238312
rect 259729 238307 259795 238310
rect 259862 238308 259868 238310
rect 259932 238308 259938 238372
rect 260598 238308 260604 238372
rect 260668 238370 260674 238372
rect 260741 238370 260807 238373
rect 260668 238368 260807 238370
rect 260668 238312 260746 238368
rect 260802 238312 260807 238368
rect 260668 238310 260807 238312
rect 260668 238308 260674 238310
rect 260741 238307 260807 238310
rect 261017 238370 261083 238373
rect 268377 238370 268443 238373
rect 261017 238368 268443 238370
rect 261017 238312 261022 238368
rect 261078 238312 268382 238368
rect 268438 238312 268443 238368
rect 261017 238310 268443 238312
rect 261017 238307 261083 238310
rect 268377 238307 268443 238310
rect 262121 238234 262187 238237
rect 263593 238236 263659 238237
rect 259318 238232 262187 238234
rect 259318 238176 262126 238232
rect 262182 238176 262187 238232
rect 259318 238174 262187 238176
rect 262121 238171 262187 238174
rect 263542 238172 263548 238236
rect 263612 238234 263659 238236
rect 266353 238234 266419 238237
rect 273437 238234 273503 238237
rect 263612 238232 263704 238234
rect 263654 238176 263704 238232
rect 263612 238174 263704 238176
rect 266353 238232 273503 238234
rect 266353 238176 266358 238232
rect 266414 238176 273442 238232
rect 273498 238176 273503 238232
rect 266353 238174 273503 238176
rect 263612 238172 263659 238174
rect 263593 238171 263659 238172
rect 266353 238171 266419 238174
rect 273437 238171 273503 238174
rect 185158 238036 185164 238100
rect 185228 238098 185234 238100
rect 222009 238098 222075 238101
rect 185228 238096 222075 238098
rect 185228 238040 222014 238096
rect 222070 238040 222075 238096
rect 185228 238038 222075 238040
rect 185228 238036 185234 238038
rect 222009 238035 222075 238038
rect 227110 238036 227116 238100
rect 227180 238098 227186 238100
rect 234286 238098 234292 238100
rect 227180 238038 234292 238098
rect 227180 238036 227186 238038
rect 234286 238036 234292 238038
rect 234356 238036 234362 238100
rect 234429 238098 234495 238101
rect 241421 238098 241487 238101
rect 234429 238096 241487 238098
rect 234429 238040 234434 238096
rect 234490 238040 241426 238096
rect 241482 238040 241487 238096
rect 234429 238038 241487 238040
rect 234429 238035 234495 238038
rect 241421 238035 241487 238038
rect 253289 238098 253355 238101
rect 258349 238098 258415 238101
rect 258758 238098 258764 238100
rect 253289 238096 256710 238098
rect 253289 238040 253294 238096
rect 253350 238040 256710 238096
rect 253289 238038 256710 238040
rect 253289 238035 253355 238038
rect 175774 237900 175780 237964
rect 175844 237962 175850 237964
rect 229737 237962 229803 237965
rect 175844 237960 229803 237962
rect 175844 237904 229742 237960
rect 229798 237904 229803 237960
rect 175844 237902 229803 237904
rect 175844 237900 175850 237902
rect 229737 237899 229803 237902
rect 230606 237900 230612 237964
rect 230676 237962 230682 237964
rect 250805 237962 250871 237965
rect 255405 237964 255471 237965
rect 255405 237962 255452 237964
rect 230676 237960 250871 237962
rect 230676 237904 250810 237960
rect 250866 237904 250871 237960
rect 230676 237902 250871 237904
rect 255360 237960 255452 237962
rect 255360 237904 255410 237960
rect 255360 237902 255452 237904
rect 230676 237900 230682 237902
rect 250805 237899 250871 237902
rect 255405 237900 255452 237902
rect 255516 237900 255522 237964
rect 256650 237962 256710 238038
rect 258349 238096 258764 238098
rect 258349 238040 258354 238096
rect 258410 238040 258764 238096
rect 258349 238038 258764 238040
rect 258349 238035 258415 238038
rect 258758 238036 258764 238038
rect 258828 238036 258834 238100
rect 260557 238098 260623 238101
rect 271229 238098 271295 238101
rect 260557 238096 271295 238098
rect 260557 238040 260562 238096
rect 260618 238040 271234 238096
rect 271290 238040 271295 238096
rect 260557 238038 271295 238040
rect 260557 238035 260623 238038
rect 271229 238035 271295 238038
rect 262806 237962 262812 237964
rect 256650 237902 262812 237962
rect 262806 237900 262812 237902
rect 262876 237900 262882 237964
rect 268326 237900 268332 237964
rect 268396 237962 268402 237964
rect 334249 237962 334315 237965
rect 268396 237960 334315 237962
rect 268396 237904 334254 237960
rect 334310 237904 334315 237960
rect 268396 237902 334315 237904
rect 268396 237900 268402 237902
rect 255405 237899 255471 237900
rect 334249 237899 334315 237902
rect 227253 237826 227319 237829
rect 215250 237824 227319 237826
rect 215250 237768 227258 237824
rect 227314 237768 227319 237824
rect 215250 237766 227319 237768
rect 206645 237690 206711 237693
rect 215250 237690 215310 237766
rect 227253 237763 227319 237766
rect 229686 237764 229692 237828
rect 229756 237826 229762 237828
rect 237189 237826 237255 237829
rect 229756 237824 237255 237826
rect 229756 237768 237194 237824
rect 237250 237768 237255 237824
rect 229756 237766 237255 237768
rect 229756 237764 229762 237766
rect 237189 237763 237255 237766
rect 251030 237764 251036 237828
rect 251100 237826 251106 237828
rect 254853 237826 254919 237829
rect 251100 237824 254919 237826
rect 251100 237768 254858 237824
rect 254914 237768 254919 237824
rect 251100 237766 254919 237768
rect 251100 237764 251106 237766
rect 254853 237763 254919 237766
rect 255589 237826 255655 237829
rect 266997 237826 267063 237829
rect 255589 237824 267063 237826
rect 255589 237768 255594 237824
rect 255650 237768 267002 237824
rect 267058 237768 267063 237824
rect 255589 237766 267063 237768
rect 255589 237763 255655 237766
rect 266997 237763 267063 237766
rect 206645 237688 215310 237690
rect 206645 237632 206650 237688
rect 206706 237632 215310 237688
rect 206645 237630 215310 237632
rect 224585 237690 224651 237693
rect 224585 237688 244290 237690
rect 224585 237632 224590 237688
rect 224646 237632 244290 237688
rect 224585 237630 244290 237632
rect 206645 237627 206711 237630
rect 224585 237627 224651 237630
rect 225689 237554 225755 237557
rect 230054 237554 230060 237556
rect 225689 237552 230060 237554
rect 225689 237496 225694 237552
rect 225750 237496 230060 237552
rect 225689 237494 230060 237496
rect 225689 237491 225755 237494
rect 230054 237492 230060 237494
rect 230124 237492 230130 237556
rect 236361 237554 236427 237557
rect 236862 237554 236868 237556
rect 236361 237552 236868 237554
rect 236361 237496 236366 237552
rect 236422 237496 236868 237552
rect 236361 237494 236868 237496
rect 236361 237491 236427 237494
rect 236862 237492 236868 237494
rect 236932 237492 236938 237556
rect 238937 237554 239003 237557
rect 239622 237554 239628 237556
rect 238937 237552 239628 237554
rect 238937 237496 238942 237552
rect 238998 237496 239628 237552
rect 238937 237494 239628 237496
rect 238937 237491 239003 237494
rect 239622 237492 239628 237494
rect 239692 237492 239698 237556
rect 244230 237554 244290 237630
rect 263174 237628 263180 237692
rect 263244 237690 263250 237692
rect 263501 237690 263567 237693
rect 263244 237688 263567 237690
rect 263244 237632 263506 237688
rect 263562 237632 263567 237688
rect 263244 237630 263567 237632
rect 263244 237628 263250 237630
rect 263501 237627 263567 237630
rect 263777 237690 263843 237693
rect 271086 237690 271092 237692
rect 263777 237688 271092 237690
rect 263777 237632 263782 237688
rect 263838 237632 271092 237688
rect 263777 237630 271092 237632
rect 263777 237627 263843 237630
rect 271086 237628 271092 237630
rect 271156 237628 271162 237692
rect 244230 237494 267290 237554
rect 232221 237418 232287 237421
rect 228406 237416 232287 237418
rect 228406 237360 232226 237416
rect 232282 237360 232287 237416
rect 228406 237358 232287 237360
rect 217409 237282 217475 237285
rect 217777 237282 217843 237285
rect 217409 237280 217843 237282
rect 217409 237224 217414 237280
rect 217470 237224 217782 237280
rect 217838 237224 217843 237280
rect 217409 237222 217843 237224
rect 217409 237219 217475 237222
rect 217777 237219 217843 237222
rect 218605 237282 218671 237285
rect 228406 237282 228466 237358
rect 232221 237355 232287 237358
rect 218605 237280 228466 237282
rect 218605 237224 218610 237280
rect 218666 237224 228466 237280
rect 218605 237222 228466 237224
rect 229645 237282 229711 237285
rect 253381 237282 253447 237285
rect 229645 237280 253447 237282
rect 229645 237224 229650 237280
rect 229706 237224 253386 237280
rect 253442 237224 253447 237280
rect 229645 237222 253447 237224
rect 267230 237282 267290 237494
rect 271781 237418 271847 237421
rect 267598 237416 271847 237418
rect 267598 237360 271786 237416
rect 271842 237360 271847 237416
rect 267598 237358 271847 237360
rect 267598 237282 267658 237358
rect 271781 237355 271847 237358
rect 284753 237418 284819 237421
rect 287646 237418 287652 237420
rect 284753 237416 287652 237418
rect 284753 237360 284758 237416
rect 284814 237360 287652 237416
rect 284753 237358 287652 237360
rect 284753 237355 284819 237358
rect 287646 237356 287652 237358
rect 287716 237356 287722 237420
rect 267230 237222 267658 237282
rect 268929 237282 268995 237285
rect 270125 237282 270191 237285
rect 333513 237282 333579 237285
rect 268929 237280 333579 237282
rect 268929 237224 268934 237280
rect 268990 237224 270130 237280
rect 270186 237224 333518 237280
rect 333574 237224 333579 237280
rect 268929 237222 333579 237224
rect 218605 237219 218671 237222
rect 229645 237219 229711 237222
rect 253381 237219 253447 237222
rect 268929 237219 268995 237222
rect 270125 237219 270191 237222
rect 333513 237219 333579 237222
rect 214649 237146 214715 237149
rect 237281 237146 237347 237149
rect 214649 237144 237347 237146
rect 214649 237088 214654 237144
rect 214710 237088 237286 237144
rect 237342 237088 237347 237144
rect 214649 237086 237347 237088
rect 214649 237083 214715 237086
rect 237281 237083 237347 237086
rect 265709 237148 265775 237149
rect 265709 237144 265756 237148
rect 265820 237146 265826 237148
rect 266905 237146 266971 237149
rect 268326 237146 268332 237148
rect 265709 237088 265714 237144
rect 265709 237084 265756 237088
rect 265820 237086 265866 237146
rect 266905 237144 268332 237146
rect 266905 237088 266910 237144
rect 266966 237088 268332 237144
rect 266905 237086 268332 237088
rect 265820 237084 265826 237086
rect 265709 237083 265775 237084
rect 266905 237083 266971 237086
rect 268326 237084 268332 237086
rect 268396 237084 268402 237148
rect 216121 237010 216187 237013
rect 236177 237010 236243 237013
rect 237925 237010 237991 237013
rect 216121 237008 236243 237010
rect 216121 236952 216126 237008
rect 216182 236952 236182 237008
rect 236238 236952 236243 237008
rect 216121 236950 236243 236952
rect 216121 236947 216187 236950
rect 236177 236947 236243 236950
rect 236364 237008 237991 237010
rect 236364 236952 237930 237008
rect 237986 236952 237991 237008
rect 236364 236950 237991 236952
rect 215109 236874 215175 236877
rect 217409 236874 217475 236877
rect 236364 236874 236424 236950
rect 237925 236947 237991 236950
rect 238385 237010 238451 237013
rect 279785 237010 279851 237013
rect 238385 237008 279851 237010
rect 238385 236952 238390 237008
rect 238446 236952 279790 237008
rect 279846 236952 279851 237008
rect 238385 236950 279851 236952
rect 238385 236947 238451 236950
rect 279785 236947 279851 236950
rect 215109 236872 215310 236874
rect 215109 236816 215114 236872
rect 215170 236816 215310 236872
rect 215109 236814 215310 236816
rect 215109 236811 215175 236814
rect 215250 236738 215310 236814
rect 217409 236872 236424 236874
rect 217409 236816 217414 236872
rect 217470 236816 236424 236872
rect 217409 236814 236424 236816
rect 217409 236811 217475 236814
rect 236494 236812 236500 236876
rect 236564 236874 236570 236876
rect 243261 236874 243327 236877
rect 283465 236874 283531 236877
rect 236564 236872 283531 236874
rect 236564 236816 243266 236872
rect 243322 236816 283470 236872
rect 283526 236816 283531 236872
rect 236564 236814 283531 236816
rect 236564 236812 236570 236814
rect 243261 236811 243327 236814
rect 283465 236811 283531 236814
rect 235165 236738 235231 236741
rect 215250 236736 235231 236738
rect 215250 236680 235170 236736
rect 235226 236680 235231 236736
rect 215250 236678 235231 236680
rect 235165 236675 235231 236678
rect 238109 236738 238175 236741
rect 239070 236738 239076 236740
rect 238109 236736 239076 236738
rect 238109 236680 238114 236736
rect 238170 236680 239076 236736
rect 238109 236678 239076 236680
rect 238109 236675 238175 236678
rect 239070 236676 239076 236678
rect 239140 236676 239146 236740
rect 240726 236676 240732 236740
rect 240796 236738 240802 236740
rect 241237 236738 241303 236741
rect 241881 236740 241947 236741
rect 241830 236738 241836 236740
rect 240796 236736 241303 236738
rect 240796 236680 241242 236736
rect 241298 236680 241303 236736
rect 240796 236678 241303 236680
rect 241790 236678 241836 236738
rect 241900 236736 241947 236740
rect 249885 236740 249951 236741
rect 249885 236738 249932 236740
rect 241942 236680 241947 236736
rect 240796 236676 240802 236678
rect 241237 236675 241303 236678
rect 241830 236676 241836 236678
rect 241900 236676 241947 236680
rect 249840 236736 249932 236738
rect 249840 236680 249890 236736
rect 249840 236678 249932 236680
rect 241881 236675 241947 236676
rect 249885 236676 249932 236678
rect 249996 236676 250002 236740
rect 252502 236676 252508 236740
rect 252572 236738 252578 236740
rect 253105 236738 253171 236741
rect 252572 236736 253171 236738
rect 252572 236680 253110 236736
rect 253166 236680 253171 236736
rect 252572 236678 253171 236680
rect 252572 236676 252578 236678
rect 249885 236675 249951 236676
rect 253105 236675 253171 236678
rect 255773 236738 255839 236741
rect 256366 236738 256372 236740
rect 255773 236736 256372 236738
rect 255773 236680 255778 236736
rect 255834 236680 256372 236736
rect 255773 236678 256372 236680
rect 255773 236675 255839 236678
rect 256366 236676 256372 236678
rect 256436 236676 256442 236740
rect 258574 236676 258580 236740
rect 258644 236738 258650 236740
rect 258993 236738 259059 236741
rect 258644 236736 259059 236738
rect 258644 236680 258998 236736
rect 259054 236680 259059 236736
rect 258644 236678 259059 236680
rect 258644 236676 258650 236678
rect 258993 236675 259059 236678
rect 264973 236738 265039 236741
rect 266118 236738 266124 236740
rect 264973 236736 266124 236738
rect 264973 236680 264978 236736
rect 265034 236680 266124 236736
rect 264973 236678 266124 236680
rect 264973 236675 265039 236678
rect 266118 236676 266124 236678
rect 266188 236676 266194 236740
rect 266629 236738 266695 236741
rect 298185 236738 298251 236741
rect 299013 236738 299079 236741
rect 266629 236736 299079 236738
rect 266629 236680 266634 236736
rect 266690 236680 298190 236736
rect 298246 236680 299018 236736
rect 299074 236680 299079 236736
rect 266629 236678 299079 236680
rect 266629 236675 266695 236678
rect 298185 236675 298251 236678
rect 299013 236675 299079 236678
rect 210969 236602 211035 236605
rect 229921 236602 229987 236605
rect 210969 236600 229987 236602
rect 210969 236544 210974 236600
rect 211030 236544 229926 236600
rect 229982 236544 229987 236600
rect 210969 236542 229987 236544
rect 210969 236539 211035 236542
rect 229921 236539 229987 236542
rect 232446 236540 232452 236604
rect 232516 236602 232522 236604
rect 252921 236602 252987 236605
rect 232516 236600 252987 236602
rect 232516 236544 252926 236600
rect 252982 236544 252987 236600
rect 232516 236542 252987 236544
rect 232516 236540 232522 236542
rect 252921 236539 252987 236542
rect 264053 236602 264119 236605
rect 294597 236602 294663 236605
rect 332041 236602 332107 236605
rect 264053 236600 332107 236602
rect 264053 236544 264058 236600
rect 264114 236544 294602 236600
rect 294658 236544 332046 236600
rect 332102 236544 332107 236600
rect 264053 236542 332107 236544
rect 264053 236539 264119 236542
rect 294597 236539 294663 236542
rect 332041 236539 332107 236542
rect 212165 236466 212231 236469
rect 229686 236466 229692 236468
rect 212165 236464 229692 236466
rect 212165 236408 212170 236464
rect 212226 236408 229692 236464
rect 212165 236406 229692 236408
rect 212165 236403 212231 236406
rect 229686 236404 229692 236406
rect 229756 236404 229762 236468
rect 248638 236404 248644 236468
rect 248708 236466 248714 236468
rect 248781 236466 248847 236469
rect 248708 236464 248847 236466
rect 248708 236408 248786 236464
rect 248842 236408 248847 236464
rect 248708 236406 248847 236408
rect 248708 236404 248714 236406
rect 248781 236403 248847 236406
rect 252093 236466 252159 236469
rect 252870 236466 252876 236468
rect 252093 236464 252876 236466
rect 252093 236408 252098 236464
rect 252154 236408 252876 236464
rect 252093 236406 252876 236408
rect 252093 236403 252159 236406
rect 252870 236404 252876 236406
rect 252940 236404 252946 236468
rect 260465 236466 260531 236469
rect 274541 236466 274607 236469
rect 260465 236464 274607 236466
rect 260465 236408 260470 236464
rect 260526 236408 274546 236464
rect 274602 236408 274607 236464
rect 260465 236406 274607 236408
rect 260465 236403 260531 236406
rect 274541 236403 274607 236406
rect 224718 236268 224724 236332
rect 224788 236330 224794 236332
rect 225873 236330 225939 236333
rect 224788 236328 225939 236330
rect 224788 236272 225878 236328
rect 225934 236272 225939 236328
rect 224788 236270 225939 236272
rect 224788 236268 224794 236270
rect 225873 236267 225939 236270
rect 234981 236330 235047 236333
rect 235206 236330 235212 236332
rect 234981 236328 235212 236330
rect 234981 236272 234986 236328
rect 235042 236272 235212 236328
rect 234981 236270 235212 236272
rect 234981 236267 235047 236270
rect 235206 236268 235212 236270
rect 235276 236330 235282 236332
rect 277945 236330 278011 236333
rect 235276 236328 278011 236330
rect 235276 236272 277950 236328
rect 278006 236272 278011 236328
rect 235276 236270 278011 236272
rect 235276 236268 235282 236270
rect 277945 236267 278011 236270
rect 220445 236194 220511 236197
rect 229645 236194 229711 236197
rect 220445 236192 229711 236194
rect 220445 236136 220450 236192
rect 220506 236136 229650 236192
rect 229706 236136 229711 236192
rect 220445 236134 229711 236136
rect 220445 236131 220511 236134
rect 229645 236131 229711 236134
rect 236177 236194 236243 236197
rect 261385 236196 261451 236197
rect 237046 236194 237052 236196
rect 236177 236192 237052 236194
rect 236177 236136 236182 236192
rect 236238 236136 237052 236192
rect 236177 236134 237052 236136
rect 236177 236131 236243 236134
rect 237046 236132 237052 236134
rect 237116 236132 237122 236196
rect 261334 236194 261340 236196
rect 261294 236134 261340 236194
rect 261404 236192 261451 236196
rect 261446 236136 261451 236192
rect 261334 236132 261340 236134
rect 261404 236132 261451 236136
rect 261385 236131 261451 236132
rect 229645 236058 229711 236061
rect 229870 236058 229876 236060
rect 229645 236056 229876 236058
rect 229645 236000 229650 236056
rect 229706 236000 229876 236056
rect 229645 235998 229876 236000
rect 229645 235995 229711 235998
rect 229870 235996 229876 235998
rect 229940 235996 229946 236060
rect 233734 235996 233740 236060
rect 233804 236058 233810 236060
rect 233877 236058 233943 236061
rect 233804 236056 233943 236058
rect 233804 236000 233882 236056
rect 233938 236000 233943 236056
rect 233804 235998 233943 236000
rect 233804 235996 233810 235998
rect 233877 235995 233943 235998
rect 234061 236058 234127 236061
rect 234470 236058 234476 236060
rect 234061 236056 234476 236058
rect 234061 236000 234066 236056
rect 234122 236000 234476 236056
rect 234061 235998 234476 236000
rect 234061 235995 234127 235998
rect 234470 235996 234476 235998
rect 234540 235996 234546 236060
rect 282913 236058 282979 236061
rect 283465 236058 283531 236061
rect 282913 236056 283531 236058
rect 282913 236000 282918 236056
rect 282974 236000 283470 236056
rect 283526 236000 283531 236056
rect 282913 235998 283531 236000
rect 282913 235995 282979 235998
rect 283465 235995 283531 235998
rect 226517 235922 226583 235925
rect 226742 235922 226748 235924
rect 226517 235920 226748 235922
rect 226517 235864 226522 235920
rect 226578 235864 226748 235920
rect 226517 235862 226748 235864
rect 226517 235859 226583 235862
rect 226742 235860 226748 235862
rect 226812 235860 226818 235924
rect 243077 235922 243143 235925
rect 274357 235922 274423 235925
rect 243077 235920 274423 235922
rect 243077 235864 243082 235920
rect 243138 235864 274362 235920
rect 274418 235864 274423 235920
rect 243077 235862 274423 235864
rect 243077 235859 243143 235862
rect 274357 235859 274423 235862
rect 274582 235860 274588 235924
rect 274652 235922 274658 235924
rect 275369 235922 275435 235925
rect 274652 235920 275435 235922
rect 274652 235864 275374 235920
rect 275430 235864 275435 235920
rect 274652 235862 275435 235864
rect 274652 235860 274658 235862
rect 275369 235859 275435 235862
rect 295333 235922 295399 235925
rect 296621 235922 296687 235925
rect 328678 235922 328684 235924
rect 295333 235920 328684 235922
rect 295333 235864 295338 235920
rect 295394 235864 296626 235920
rect 296682 235864 328684 235920
rect 295333 235862 328684 235864
rect 295333 235859 295399 235862
rect 296621 235859 296687 235862
rect 328678 235860 328684 235862
rect 328748 235860 328754 235924
rect 203977 235786 204043 235789
rect 228449 235786 228515 235789
rect 203977 235784 228515 235786
rect 203977 235728 203982 235784
rect 204038 235728 228454 235784
rect 228510 235728 228515 235784
rect 203977 235726 228515 235728
rect 203977 235723 204043 235726
rect 228449 235723 228515 235726
rect 230473 235786 230539 235789
rect 230606 235786 230612 235788
rect 230473 235784 230612 235786
rect 230473 235728 230478 235784
rect 230534 235728 230612 235784
rect 230473 235726 230612 235728
rect 230473 235723 230539 235726
rect 230606 235724 230612 235726
rect 230676 235724 230682 235788
rect 232630 235724 232636 235788
rect 232700 235786 232706 235788
rect 232865 235786 232931 235789
rect 232700 235784 232931 235786
rect 232700 235728 232870 235784
rect 232926 235728 232931 235784
rect 232700 235726 232931 235728
rect 232700 235724 232706 235726
rect 232865 235723 232931 235726
rect 237465 235786 237531 235789
rect 238518 235786 238524 235788
rect 237465 235784 238524 235786
rect 237465 235728 237470 235784
rect 237526 235728 238524 235784
rect 237465 235726 238524 235728
rect 237465 235723 237531 235726
rect 238518 235724 238524 235726
rect 238588 235724 238594 235788
rect 253238 235724 253244 235788
rect 253308 235786 253314 235788
rect 253657 235786 253723 235789
rect 253308 235784 253723 235786
rect 253308 235728 253662 235784
rect 253718 235728 253723 235784
rect 253308 235726 253723 235728
rect 253308 235724 253314 235726
rect 253657 235723 253723 235726
rect 257245 235786 257311 235789
rect 269113 235786 269179 235789
rect 257245 235784 269179 235786
rect 257245 235728 257250 235784
rect 257306 235728 269118 235784
rect 269174 235728 269179 235784
rect 257245 235726 269179 235728
rect 257245 235723 257311 235726
rect 269113 235723 269179 235726
rect 183134 235588 183140 235652
rect 183204 235650 183210 235652
rect 209681 235650 209747 235653
rect 238753 235650 238819 235653
rect 183204 235648 238819 235650
rect 183204 235592 209686 235648
rect 209742 235592 238758 235648
rect 238814 235592 238819 235648
rect 183204 235590 238819 235592
rect 183204 235588 183210 235590
rect 209681 235587 209747 235590
rect 238753 235587 238819 235590
rect 261702 235588 261708 235652
rect 261772 235650 261778 235652
rect 269573 235650 269639 235653
rect 261772 235648 269639 235650
rect 261772 235592 269578 235648
rect 269634 235592 269639 235648
rect 261772 235590 269639 235592
rect 261772 235588 261778 235590
rect 269573 235587 269639 235590
rect 169518 235452 169524 235516
rect 169588 235514 169594 235516
rect 203977 235514 204043 235517
rect 235022 235514 235028 235516
rect 169588 235512 204043 235514
rect 169588 235456 203982 235512
rect 204038 235456 204043 235512
rect 169588 235454 204043 235456
rect 169588 235452 169594 235454
rect 203977 235451 204043 235454
rect 215250 235454 235028 235514
rect 158345 235378 158411 235381
rect 214833 235378 214899 235381
rect 158345 235376 214899 235378
rect 158345 235320 158350 235376
rect 158406 235320 214838 235376
rect 214894 235320 214899 235376
rect 158345 235318 214899 235320
rect 158345 235315 158411 235318
rect 214833 235315 214899 235318
rect 176510 235180 176516 235244
rect 176580 235242 176586 235244
rect 215250 235242 215310 235454
rect 235022 235452 235028 235454
rect 235092 235452 235098 235516
rect 238661 235514 238727 235517
rect 239622 235514 239628 235516
rect 238661 235512 239628 235514
rect 238661 235456 238666 235512
rect 238722 235456 239628 235512
rect 238661 235454 239628 235456
rect 238661 235451 238727 235454
rect 239622 235452 239628 235454
rect 239692 235452 239698 235516
rect 266905 235514 266971 235517
rect 267917 235514 267983 235517
rect 328862 235514 328868 235516
rect 266905 235512 328868 235514
rect 266905 235456 266910 235512
rect 266966 235456 267922 235512
rect 267978 235456 328868 235512
rect 266905 235454 328868 235456
rect 266905 235451 266971 235454
rect 267917 235451 267983 235454
rect 328862 235452 328868 235454
rect 328932 235452 328938 235516
rect 233049 235378 233115 235381
rect 243077 235378 243143 235381
rect 233049 235376 243143 235378
rect 233049 235320 233054 235376
rect 233110 235320 243082 235376
rect 243138 235320 243143 235376
rect 233049 235318 243143 235320
rect 233049 235315 233115 235318
rect 243077 235315 243143 235318
rect 244774 235316 244780 235380
rect 244844 235378 244850 235380
rect 257245 235378 257311 235381
rect 244844 235376 257311 235378
rect 244844 235320 257250 235376
rect 257306 235320 257311 235376
rect 244844 235318 257311 235320
rect 244844 235316 244850 235318
rect 257245 235315 257311 235318
rect 265801 235378 265867 235381
rect 270953 235378 271019 235381
rect 332685 235378 332751 235381
rect 265801 235376 332751 235378
rect 265801 235320 265806 235376
rect 265862 235320 270958 235376
rect 271014 235320 332690 235376
rect 332746 235320 332751 235376
rect 265801 235318 332751 235320
rect 265801 235315 265867 235318
rect 270953 235315 271019 235318
rect 332685 235315 332751 235318
rect 176580 235182 215310 235242
rect 236637 235242 236703 235245
rect 253013 235242 253079 235245
rect 236637 235240 253079 235242
rect 236637 235184 236642 235240
rect 236698 235184 253018 235240
rect 253074 235184 253079 235240
rect 236637 235182 253079 235184
rect 176580 235180 176586 235182
rect 236637 235179 236703 235182
rect 253013 235179 253079 235182
rect 263317 235242 263383 235245
rect 267825 235242 267891 235245
rect 331489 235242 331555 235245
rect 263317 235240 331555 235242
rect 263317 235184 263322 235240
rect 263378 235184 267830 235240
rect 267886 235184 331494 235240
rect 331550 235184 331555 235240
rect 263317 235182 331555 235184
rect 263317 235179 263383 235182
rect 267825 235179 267891 235182
rect 331489 235179 331555 235182
rect 257102 235044 257108 235108
rect 257172 235106 257178 235108
rect 257521 235106 257587 235109
rect 257172 235104 257587 235106
rect 257172 235048 257526 235104
rect 257582 235048 257587 235104
rect 257172 235046 257587 235048
rect 257172 235044 257178 235046
rect 257521 235043 257587 235046
rect 261518 235044 261524 235108
rect 261588 235106 261594 235108
rect 261845 235106 261911 235109
rect 261588 235104 261911 235106
rect 261588 235048 261850 235104
rect 261906 235048 261911 235104
rect 261588 235046 261911 235048
rect 261588 235044 261594 235046
rect 261845 235043 261911 235046
rect 266997 235106 267063 235109
rect 268101 235106 268167 235109
rect 282085 235106 282151 235109
rect 266997 235104 282151 235106
rect 266997 235048 267002 235104
rect 267058 235048 268106 235104
rect 268162 235048 282090 235104
rect 282146 235048 282151 235104
rect 266997 235046 282151 235048
rect 266997 235043 267063 235046
rect 268101 235043 268167 235046
rect 282085 235043 282151 235046
rect 183318 234636 183324 234700
rect 183388 234698 183394 234700
rect 243118 234698 243124 234700
rect 183388 234638 243124 234698
rect 183388 234636 183394 234638
rect 243118 234636 243124 234638
rect 243188 234636 243194 234700
rect 182950 234500 182956 234564
rect 183020 234562 183026 234564
rect 208761 234562 208827 234565
rect 209405 234562 209471 234565
rect 183020 234560 209471 234562
rect 183020 234504 208766 234560
rect 208822 234504 209410 234560
rect 209466 234504 209471 234560
rect 183020 234502 209471 234504
rect 183020 234500 183026 234502
rect 208761 234499 208827 234502
rect 209405 234499 209471 234502
rect 261150 234500 261156 234564
rect 261220 234562 261226 234564
rect 262489 234562 262555 234565
rect 261220 234560 262555 234562
rect 261220 234504 262494 234560
rect 262550 234504 262555 234560
rect 261220 234502 262555 234504
rect 261220 234500 261226 234502
rect 262489 234499 262555 234502
rect 181478 234364 181484 234428
rect 181548 234426 181554 234428
rect 210141 234426 210207 234429
rect 241789 234426 241855 234429
rect 181548 234424 241855 234426
rect 181548 234368 210146 234424
rect 210202 234368 241794 234424
rect 241850 234368 241855 234424
rect 181548 234366 241855 234368
rect 181548 234364 181554 234366
rect 210141 234363 210207 234366
rect 241789 234363 241855 234366
rect 254894 234364 254900 234428
rect 254964 234426 254970 234428
rect 270309 234426 270375 234429
rect 254964 234424 270375 234426
rect 254964 234368 270314 234424
rect 270370 234368 270375 234424
rect 254964 234366 270375 234368
rect 254964 234364 254970 234366
rect 270309 234363 270375 234366
rect 181294 234228 181300 234292
rect 181364 234290 181370 234292
rect 240869 234290 240935 234293
rect 181364 234288 240935 234290
rect 181364 234232 240874 234288
rect 240930 234232 240935 234288
rect 181364 234230 240935 234232
rect 181364 234228 181370 234230
rect 240869 234227 240935 234230
rect 248321 234290 248387 234293
rect 250110 234290 250116 234292
rect 248321 234288 250116 234290
rect 248321 234232 248326 234288
rect 248382 234232 250116 234288
rect 248321 234230 250116 234232
rect 248321 234227 248387 234230
rect 250110 234228 250116 234230
rect 250180 234290 250186 234292
rect 310145 234290 310211 234293
rect 250180 234288 310211 234290
rect 250180 234232 310150 234288
rect 310206 234232 310211 234288
rect 250180 234230 310211 234232
rect 250180 234228 250186 234230
rect 310145 234227 310211 234230
rect 182766 234092 182772 234156
rect 182836 234154 182842 234156
rect 242801 234154 242867 234157
rect 182836 234152 242867 234154
rect 182836 234096 242806 234152
rect 242862 234096 242867 234152
rect 182836 234094 242867 234096
rect 182836 234092 182842 234094
rect 242801 234091 242867 234094
rect 173750 233956 173756 234020
rect 173820 234018 173826 234020
rect 233366 234018 233372 234020
rect 173820 233958 233372 234018
rect 173820 233956 173826 233958
rect 233366 233956 233372 233958
rect 233436 233956 233442 234020
rect 266813 234018 266879 234021
rect 282453 234018 282519 234021
rect 331305 234018 331371 234021
rect 266813 234016 331371 234018
rect 266813 233960 266818 234016
rect 266874 233960 282458 234016
rect 282514 233960 331310 234016
rect 331366 233960 331371 234016
rect 266813 233958 331371 233960
rect 266813 233955 266879 233958
rect 282453 233955 282519 233958
rect 331305 233955 331371 233958
rect 180558 233820 180564 233884
rect 180628 233882 180634 233884
rect 240685 233882 240751 233885
rect 180628 233880 240751 233882
rect 180628 233824 240690 233880
rect 240746 233824 240751 233880
rect 180628 233822 240751 233824
rect 180628 233820 180634 233822
rect 240685 233819 240751 233822
rect 247677 233882 247743 233885
rect 263777 233882 263843 233885
rect 247677 233880 263843 233882
rect 247677 233824 247682 233880
rect 247738 233824 263782 233880
rect 263838 233824 263843 233880
rect 247677 233822 263843 233824
rect 247677 233819 247743 233822
rect 263777 233819 263843 233822
rect 266077 233882 266143 233885
rect 285121 233882 285187 233885
rect 335537 233882 335603 233885
rect 266077 233880 335603 233882
rect 266077 233824 266082 233880
rect 266138 233824 285126 233880
rect 285182 233824 335542 233880
rect 335598 233824 335603 233880
rect 266077 233822 335603 233824
rect 266077 233819 266143 233822
rect 285121 233819 285187 233822
rect 335537 233819 335603 233822
rect 184422 233684 184428 233748
rect 184492 233746 184498 233748
rect 208485 233746 208551 233749
rect 184492 233744 208551 233746
rect 184492 233688 208490 233744
rect 208546 233688 208551 233744
rect 184492 233686 208551 233688
rect 184492 233684 184498 233686
rect 208485 233683 208551 233686
rect 221457 233746 221523 233749
rect 235390 233746 235396 233748
rect 221457 233744 235396 233746
rect 221457 233688 221462 233744
rect 221518 233688 235396 233744
rect 221457 233686 235396 233688
rect 221457 233683 221523 233686
rect 235390 233684 235396 233686
rect 235460 233684 235466 233748
rect 208761 233610 208827 233613
rect 243353 233610 243419 233613
rect 208761 233608 243419 233610
rect 208761 233552 208766 233608
rect 208822 233552 243358 233608
rect 243414 233552 243419 233608
rect 208761 233550 243419 233552
rect 208761 233547 208827 233550
rect 243353 233547 243419 233550
rect 258574 233276 258580 233340
rect 258644 233338 258650 233340
rect 259177 233338 259243 233341
rect 258644 233336 259243 233338
rect 258644 233280 259182 233336
rect 259238 233280 259243 233336
rect 258644 233278 259243 233280
rect 258644 233276 258650 233278
rect 259177 233275 259243 233278
rect 165470 233140 165476 233204
rect 165540 233202 165546 233204
rect 193765 233202 193831 233205
rect 165540 233200 193831 233202
rect 165540 233144 193770 233200
rect 193826 233144 193831 233200
rect 165540 233142 193831 233144
rect 165540 233140 165546 233142
rect 193765 233139 193831 233142
rect 240542 233140 240548 233204
rect 240612 233202 240618 233204
rect 240685 233202 240751 233205
rect 240612 233200 240751 233202
rect 240612 233144 240690 233200
rect 240746 233144 240751 233200
rect 240612 233142 240751 233144
rect 240612 233140 240618 233142
rect 240685 233139 240751 233142
rect 245929 233202 245995 233205
rect 246430 233202 246436 233204
rect 245929 233200 246436 233202
rect 245929 233144 245934 233200
rect 245990 233144 246436 233200
rect 245929 233142 246436 233144
rect 245929 233139 245995 233142
rect 246430 233140 246436 233142
rect 246500 233140 246506 233204
rect 255221 233202 255287 233205
rect 332869 233202 332935 233205
rect 255221 233200 332935 233202
rect 255221 233144 255226 233200
rect 255282 233144 332874 233200
rect 332930 233144 332935 233200
rect 255221 233142 332935 233144
rect 255221 233139 255287 233142
rect 332869 233139 332935 233142
rect 190862 233004 190868 233068
rect 190932 233066 190938 233068
rect 222009 233066 222075 233069
rect 190932 233064 222075 233066
rect 190932 233008 222014 233064
rect 222070 233008 222075 233064
rect 190932 233006 222075 233008
rect 190932 233004 190938 233006
rect 222009 233003 222075 233006
rect 261661 233066 261727 233069
rect 333973 233066 334039 233069
rect 261661 233064 334039 233066
rect 261661 233008 261666 233064
rect 261722 233008 333978 233064
rect 334034 233008 334039 233064
rect 261661 233006 334039 233008
rect 261661 233003 261727 233006
rect 333973 233003 334039 233006
rect 175038 232868 175044 232932
rect 175108 232930 175114 232932
rect 233969 232930 234035 232933
rect 175108 232928 234035 232930
rect 175108 232872 233974 232928
rect 234030 232872 234035 232928
rect 175108 232870 234035 232872
rect 175108 232868 175114 232870
rect 233969 232867 234035 232870
rect 162894 232732 162900 232796
rect 162964 232794 162970 232796
rect 192477 232794 192543 232797
rect 162964 232792 192543 232794
rect 162964 232736 192482 232792
rect 192538 232736 192543 232792
rect 162964 232734 192543 232736
rect 162964 232732 162970 232734
rect 192477 232731 192543 232734
rect 193622 232732 193628 232796
rect 193692 232794 193698 232796
rect 220445 232794 220511 232797
rect 193692 232792 220511 232794
rect 193692 232736 220450 232792
rect 220506 232736 220511 232792
rect 193692 232734 220511 232736
rect 193692 232732 193698 232734
rect 220445 232731 220511 232734
rect 250897 232794 250963 232797
rect 299974 232794 299980 232796
rect 250897 232792 299980 232794
rect 250897 232736 250902 232792
rect 250958 232736 299980 232792
rect 250897 232734 299980 232736
rect 250897 232731 250963 232734
rect 299974 232732 299980 232734
rect 300044 232732 300050 232796
rect 163814 232596 163820 232660
rect 163884 232658 163890 232660
rect 223573 232658 223639 232661
rect 163884 232656 223639 232658
rect 163884 232600 223578 232656
rect 223634 232600 223639 232656
rect 163884 232598 223639 232600
rect 163884 232596 163890 232598
rect 223573 232595 223639 232598
rect 265750 232596 265756 232660
rect 265820 232658 265826 232660
rect 330334 232658 330340 232660
rect 265820 232598 330340 232658
rect 265820 232596 265826 232598
rect 330334 232596 330340 232598
rect 330404 232596 330410 232660
rect 168230 232460 168236 232524
rect 168300 232522 168306 232524
rect 228357 232522 228423 232525
rect 168300 232520 228423 232522
rect 168300 232464 228362 232520
rect 228418 232464 228423 232520
rect 168300 232462 228423 232464
rect 168300 232460 168306 232462
rect 228357 232459 228423 232462
rect 191414 232324 191420 232388
rect 191484 232386 191490 232388
rect 218697 232386 218763 232389
rect 191484 232384 218763 232386
rect 191484 232328 218702 232384
rect 218758 232328 218763 232384
rect 191484 232326 218763 232328
rect 191484 232324 191490 232326
rect 218697 232323 218763 232326
rect 221917 232386 221983 232389
rect 254485 232386 254551 232389
rect 221917 232384 254551 232386
rect 221917 232328 221922 232384
rect 221978 232328 254490 232384
rect 254546 232328 254551 232384
rect 221917 232326 254551 232328
rect 221917 232323 221983 232326
rect 254485 232323 254551 232326
rect 259269 232386 259335 232389
rect 259494 232386 259500 232388
rect 259269 232384 259500 232386
rect 259269 232328 259274 232384
rect 259330 232328 259500 232384
rect 259269 232326 259500 232328
rect 259269 232323 259335 232326
rect 259494 232324 259500 232326
rect 259564 232324 259570 232388
rect 579613 232386 579679 232389
rect 583520 232386 584960 232476
rect 579613 232384 584960 232386
rect 579613 232328 579618 232384
rect 579674 232328 584960 232384
rect 579613 232326 584960 232328
rect 579613 232323 579679 232326
rect 192702 232188 192708 232252
rect 192772 232250 192778 232252
rect 252134 232250 252140 232252
rect 192772 232190 252140 232250
rect 192772 232188 192778 232190
rect 252134 232188 252140 232190
rect 252204 232188 252210 232252
rect 259729 232250 259795 232253
rect 262438 232250 262444 232252
rect 259729 232248 262444 232250
rect 259729 232192 259734 232248
rect 259790 232192 262444 232248
rect 259729 232190 262444 232192
rect 259729 232187 259795 232190
rect 262438 232188 262444 232190
rect 262508 232188 262514 232252
rect 583520 232236 584960 232326
rect 250069 231978 250135 231981
rect 250897 231978 250963 231981
rect 250069 231976 250963 231978
rect 250069 231920 250074 231976
rect 250130 231920 250902 231976
rect 250958 231920 250963 231976
rect 250069 231918 250963 231920
rect 250069 231915 250135 231918
rect 250897 231915 250963 231918
rect 168046 231780 168052 231844
rect 168116 231842 168122 231844
rect 205449 231842 205515 231845
rect 227161 231842 227227 231845
rect 168116 231840 227227 231842
rect 168116 231784 205454 231840
rect 205510 231784 227166 231840
rect 227222 231784 227227 231840
rect 168116 231782 227227 231784
rect 168116 231780 168122 231782
rect 205449 231779 205515 231782
rect 227161 231779 227227 231782
rect 265249 231842 265315 231845
rect 265709 231842 265775 231845
rect 331213 231842 331279 231845
rect 265249 231840 331279 231842
rect 265249 231784 265254 231840
rect 265310 231784 265714 231840
rect 265770 231784 331218 231840
rect 331274 231784 331279 231840
rect 265249 231782 331279 231784
rect 265249 231779 265315 231782
rect 265709 231779 265775 231782
rect 331213 231779 331279 231782
rect 159817 231706 159883 231709
rect 202505 231706 202571 231709
rect 227846 231706 227852 231708
rect 159817 231704 227852 231706
rect 159817 231648 159822 231704
rect 159878 231648 202510 231704
rect 202566 231648 227852 231704
rect 159817 231646 227852 231648
rect 159817 231643 159883 231646
rect 202505 231643 202571 231646
rect 227846 231644 227852 231646
rect 227916 231644 227922 231708
rect 234470 231644 234476 231708
rect 234540 231706 234546 231708
rect 281073 231706 281139 231709
rect 234540 231704 281139 231706
rect 234540 231648 281078 231704
rect 281134 231648 281139 231704
rect 234540 231646 281139 231648
rect 234540 231644 234546 231646
rect 281073 231643 281139 231646
rect 172278 231508 172284 231572
rect 172348 231570 172354 231572
rect 231117 231570 231183 231573
rect 172348 231568 231183 231570
rect 172348 231512 231122 231568
rect 231178 231512 231183 231568
rect 172348 231510 231183 231512
rect 172348 231508 172354 231510
rect 231117 231507 231183 231510
rect 256969 231570 257035 231573
rect 295926 231570 295932 231572
rect 256969 231568 295932 231570
rect 256969 231512 256974 231568
rect 257030 231512 295932 231568
rect 256969 231510 295932 231512
rect 256969 231507 257035 231510
rect 295926 231508 295932 231510
rect 295996 231508 296002 231572
rect 174854 231372 174860 231436
rect 174924 231434 174930 231436
rect 233785 231434 233851 231437
rect 174924 231432 233851 231434
rect 174924 231376 233790 231432
rect 233846 231376 233851 231432
rect 174924 231374 233851 231376
rect 174924 231372 174930 231374
rect 233785 231371 233851 231374
rect 252553 231434 252619 231437
rect 255681 231434 255747 231437
rect 271689 231434 271755 231437
rect 252553 231432 271755 231434
rect 252553 231376 252558 231432
rect 252614 231376 255686 231432
rect 255742 231376 271694 231432
rect 271750 231376 271755 231432
rect 252553 231374 271755 231376
rect 252553 231371 252619 231374
rect 255681 231371 255747 231374
rect 271689 231371 271755 231374
rect 166758 231236 166764 231300
rect 166828 231298 166834 231300
rect 225597 231298 225663 231301
rect 166828 231296 225663 231298
rect 166828 231240 225602 231296
rect 225658 231240 225663 231296
rect 166828 231238 225663 231240
rect 166828 231236 166834 231238
rect 225597 231235 225663 231238
rect 170622 231100 170628 231164
rect 170692 231162 170698 231164
rect 230841 231162 230907 231165
rect 170692 231160 230907 231162
rect 170692 231104 230846 231160
rect 230902 231104 230907 231160
rect 170692 231102 230907 231104
rect 170692 231100 170698 231102
rect 230841 231099 230907 231102
rect 258809 231162 258875 231165
rect 272609 231162 272675 231165
rect 286685 231162 286751 231165
rect 258809 231160 286751 231162
rect 258809 231104 258814 231160
rect 258870 231104 272614 231160
rect 272670 231104 286690 231160
rect 286746 231104 286751 231160
rect 258809 231102 286751 231104
rect 258809 231099 258875 231102
rect 272609 231099 272675 231102
rect 286685 231099 286751 231102
rect 262305 230890 262371 230893
rect 262990 230890 262996 230892
rect 262305 230888 262996 230890
rect 262305 230832 262310 230888
rect 262366 230832 262996 230888
rect 262305 230830 262996 230832
rect 262305 230827 262371 230830
rect 262990 230828 262996 230830
rect 263060 230828 263066 230892
rect 226885 230482 226951 230485
rect 209730 230480 226951 230482
rect 209730 230424 226890 230480
rect 226946 230424 226951 230480
rect 209730 230422 226951 230424
rect 166574 230012 166580 230076
rect 166644 230074 166650 230076
rect 205265 230074 205331 230077
rect 209730 230074 209790 230422
rect 226885 230419 226951 230422
rect 255773 230482 255839 230485
rect 256141 230482 256207 230485
rect 272793 230482 272859 230485
rect 255773 230480 272859 230482
rect 255773 230424 255778 230480
rect 255834 230424 256146 230480
rect 256202 230424 272798 230480
rect 272854 230424 272859 230480
rect 255773 230422 272859 230424
rect 255773 230419 255839 230422
rect 256141 230419 256207 230422
rect 272793 230419 272859 230422
rect 241830 230346 241836 230348
rect 166644 230072 209790 230074
rect 166644 230016 205270 230072
rect 205326 230016 209790 230072
rect 166644 230014 209790 230016
rect 238710 230286 241836 230346
rect 166644 230012 166650 230014
rect 205265 230011 205331 230014
rect 173566 229876 173572 229940
rect 173636 229938 173642 229940
rect 233233 229938 233299 229941
rect 173636 229936 233299 229938
rect 173636 229880 233238 229936
rect 233294 229880 233299 229936
rect 173636 229878 233299 229880
rect 173636 229876 173642 229878
rect 233233 229875 233299 229878
rect 150341 229802 150407 229805
rect 225086 229802 225092 229804
rect 150341 229800 225092 229802
rect 150341 229744 150346 229800
rect 150402 229744 225092 229800
rect 150341 229742 225092 229744
rect 150341 229739 150407 229742
rect 225086 229740 225092 229742
rect 225156 229740 225162 229804
rect 235349 229802 235415 229805
rect 238710 229802 238770 230286
rect 241830 230284 241836 230286
rect 241900 230346 241906 230348
rect 300301 230346 300367 230349
rect 241900 230344 300367 230346
rect 241900 230288 300306 230344
rect 300362 230288 300367 230344
rect 241900 230286 300367 230288
rect 241900 230284 241906 230286
rect 300301 230283 300367 230286
rect 262857 230212 262923 230213
rect 262806 230210 262812 230212
rect 262730 230150 262812 230210
rect 262876 230210 262923 230212
rect 310462 230210 310468 230212
rect 262876 230208 310468 230210
rect 262918 230152 310468 230208
rect 262806 230148 262812 230150
rect 262876 230150 310468 230152
rect 262876 230148 262923 230150
rect 310462 230148 310468 230150
rect 310532 230148 310538 230212
rect 262857 230147 262923 230148
rect 252461 230076 252527 230077
rect 252461 230074 252508 230076
rect 252380 230072 252508 230074
rect 252572 230074 252578 230076
rect 294781 230074 294847 230077
rect 252572 230072 294847 230074
rect 252380 230016 252466 230072
rect 252572 230016 294786 230072
rect 294842 230016 294847 230072
rect 252380 230014 252508 230016
rect 252461 230012 252508 230014
rect 252572 230014 294847 230016
rect 252572 230012 252578 230014
rect 252461 230011 252527 230012
rect 294781 230011 294847 230014
rect 267181 229938 267247 229941
rect 268009 229938 268075 229941
rect 327533 229938 327599 229941
rect 267181 229936 327599 229938
rect 267181 229880 267186 229936
rect 267242 229880 268014 229936
rect 268070 229880 327538 229936
rect 327594 229880 327599 229936
rect 267181 229878 327599 229880
rect 267181 229875 267247 229878
rect 268009 229875 268075 229878
rect 327533 229875 327599 229878
rect 235349 229800 238770 229802
rect 235349 229744 235354 229800
rect 235410 229744 238770 229800
rect 235349 229742 238770 229744
rect 235349 229739 235415 229742
rect 262438 229740 262444 229804
rect 262508 229802 262514 229804
rect 322381 229802 322447 229805
rect 262508 229800 322447 229802
rect 262508 229744 322386 229800
rect 322442 229744 322447 229800
rect 262508 229742 322447 229744
rect 262508 229740 262514 229742
rect 322381 229739 322447 229742
rect 224493 229530 224559 229533
rect 224493 229528 224602 229530
rect 224493 229472 224498 229528
rect 224554 229472 224602 229528
rect 224493 229467 224602 229472
rect 224542 229397 224602 229467
rect 224493 229392 224602 229397
rect 224493 229336 224498 229392
rect 224554 229336 224602 229392
rect 224493 229334 224602 229336
rect 224493 229331 224559 229334
rect 205357 228986 205423 228989
rect 228173 228986 228239 228989
rect 205357 228984 228239 228986
rect 205357 228928 205362 228984
rect 205418 228928 228178 228984
rect 228234 228928 228239 228984
rect 205357 228926 228239 228928
rect 205357 228923 205423 228926
rect 228173 228923 228239 228926
rect 265617 228986 265683 228989
rect 329833 228986 329899 228989
rect 265617 228984 329899 228986
rect 265617 228928 265622 228984
rect 265678 228928 329838 228984
rect 329894 228928 329899 228984
rect 265617 228926 329899 228928
rect 265617 228923 265683 228926
rect 329833 228923 329899 228926
rect 265617 228850 265683 228853
rect 265985 228850 266051 228853
rect 326337 228850 326403 228853
rect 265617 228848 326403 228850
rect 265617 228792 265622 228848
rect 265678 228792 265990 228848
rect 266046 228792 326342 228848
rect 326398 228792 326403 228848
rect 265617 228790 326403 228792
rect 265617 228787 265683 228790
rect 265985 228787 266051 228790
rect 326337 228787 326403 228790
rect 267365 228714 267431 228717
rect 327574 228714 327580 228716
rect 267365 228712 327580 228714
rect 267365 228656 267370 228712
rect 267426 228656 327580 228712
rect 267365 228654 327580 228656
rect 267365 228651 267431 228654
rect 327574 228652 327580 228654
rect 327644 228652 327650 228716
rect 248781 228578 248847 228581
rect 248965 228578 249031 228581
rect 307702 228578 307708 228580
rect 248781 228576 307708 228578
rect 248781 228520 248786 228576
rect 248842 228520 248970 228576
rect 249026 228520 307708 228576
rect 248781 228518 307708 228520
rect 248781 228515 248847 228518
rect 248965 228515 249031 228518
rect 307702 228516 307708 228518
rect 307772 228516 307778 228580
rect 249333 228442 249399 228445
rect 252870 228442 252876 228444
rect 249333 228440 252876 228442
rect 249333 228384 249338 228440
rect 249394 228384 252876 228440
rect 249333 228382 252876 228384
rect 249333 228379 249399 228382
rect 252870 228380 252876 228382
rect 252940 228442 252946 228444
rect 307109 228442 307175 228445
rect 252940 228440 307175 228442
rect 252940 228384 307114 228440
rect 307170 228384 307175 228440
rect 252940 228382 307175 228384
rect 252940 228380 252946 228382
rect 307109 228379 307175 228382
rect 158253 228306 158319 228309
rect 205357 228306 205423 228309
rect 158253 228304 205423 228306
rect 158253 228248 158258 228304
rect 158314 228248 205362 228304
rect 205418 228248 205423 228304
rect 158253 228246 205423 228248
rect 158253 228243 158319 228246
rect 205357 228243 205423 228246
rect 220077 228306 220143 228309
rect 242382 228306 242388 228308
rect 220077 228304 242388 228306
rect 220077 228248 220082 228304
rect 220138 228248 242388 228304
rect 220077 228246 242388 228248
rect 220077 228243 220143 228246
rect 242382 228244 242388 228246
rect 242452 228244 242458 228308
rect 249742 228244 249748 228308
rect 249812 228306 249818 228308
rect 250846 228306 250852 228308
rect 249812 228246 250852 228306
rect 249812 228244 249818 228246
rect 250846 228244 250852 228246
rect 250916 228306 250922 228308
rect 278865 228306 278931 228309
rect 250916 228304 278931 228306
rect 250916 228248 278870 228304
rect 278926 228248 278931 228304
rect 250916 228246 278931 228248
rect 250916 228244 250922 228246
rect 278865 228243 278931 228246
rect -960 227884 480 228124
rect 258574 227564 258580 227628
rect 258644 227626 258650 227628
rect 336825 227626 336891 227629
rect 258644 227624 336891 227626
rect 258644 227568 336830 227624
rect 336886 227568 336891 227624
rect 258644 227566 336891 227568
rect 258644 227564 258650 227566
rect 336825 227563 336891 227566
rect 267273 227490 267339 227493
rect 336733 227490 336799 227493
rect 267273 227488 336799 227490
rect 267273 227432 267278 227488
rect 267334 227432 336738 227488
rect 336794 227432 336799 227488
rect 267273 227430 336799 227432
rect 267273 227427 267339 227430
rect 336733 227427 336799 227430
rect 229737 227354 229803 227357
rect 249742 227354 249748 227356
rect 229737 227352 249748 227354
rect 229737 227296 229742 227352
rect 229798 227296 249748 227352
rect 229737 227294 249748 227296
rect 229737 227291 229803 227294
rect 249742 227292 249748 227294
rect 249812 227292 249818 227356
rect 259913 227354 259979 227357
rect 328494 227354 328500 227356
rect 259913 227352 328500 227354
rect 259913 227296 259918 227352
rect 259974 227296 328500 227352
rect 259913 227294 328500 227296
rect 259913 227291 259979 227294
rect 328494 227292 328500 227294
rect 328564 227292 328570 227356
rect 249190 227156 249196 227220
rect 249260 227218 249266 227220
rect 295057 227218 295123 227221
rect 249260 227216 295123 227218
rect 249260 227160 295062 227216
rect 295118 227160 295123 227216
rect 249260 227158 295123 227160
rect 249260 227156 249266 227158
rect 295057 227155 295123 227158
rect 241973 227082 242039 227085
rect 285305 227082 285371 227085
rect 241973 227080 285371 227082
rect 241973 227024 241978 227080
rect 242034 227024 285310 227080
rect 285366 227024 285371 227080
rect 241973 227022 285371 227024
rect 241973 227019 242039 227022
rect 285305 227019 285371 227022
rect 190310 226884 190316 226948
rect 190380 226946 190386 226948
rect 249190 226946 249196 226948
rect 190380 226886 249196 226946
rect 190380 226884 190386 226886
rect 249190 226884 249196 226886
rect 249260 226884 249266 226948
rect 236821 226810 236887 226813
rect 264605 226810 264671 226813
rect 236821 226808 264671 226810
rect 236821 226752 236826 226808
rect 236882 226752 264610 226808
rect 264666 226752 264671 226808
rect 236821 226750 264671 226752
rect 236821 226747 236887 226750
rect 264605 226747 264671 226750
rect 181110 226340 181116 226404
rect 181180 226402 181186 226404
rect 241237 226402 241303 226405
rect 241973 226402 242039 226405
rect 181180 226400 242039 226402
rect 181180 226344 241242 226400
rect 241298 226344 241978 226400
rect 242034 226344 242039 226400
rect 181180 226342 242039 226344
rect 181180 226340 181186 226342
rect 241237 226339 241303 226342
rect 241973 226339 242039 226342
rect 201309 226266 201375 226269
rect 224309 226266 224375 226269
rect 200070 226264 224375 226266
rect 200070 226208 201314 226264
rect 201370 226208 224314 226264
rect 224370 226208 224375 226264
rect 200070 226206 224375 226208
rect 163446 225660 163452 225724
rect 163516 225722 163522 225724
rect 200070 225722 200130 226206
rect 201309 226203 201375 226206
rect 224309 226203 224375 226206
rect 246982 226204 246988 226268
rect 247052 226266 247058 226268
rect 248270 226266 248276 226268
rect 247052 226206 248276 226266
rect 247052 226204 247058 226206
rect 248270 226204 248276 226206
rect 248340 226204 248346 226268
rect 260414 226204 260420 226268
rect 260484 226266 260490 226268
rect 260925 226266 260991 226269
rect 260484 226264 260991 226266
rect 260484 226208 260930 226264
rect 260986 226208 260991 226264
rect 260484 226206 260991 226208
rect 260484 226204 260490 226206
rect 260925 226203 260991 226206
rect 264329 226266 264395 226269
rect 323526 226266 323532 226268
rect 264329 226264 323532 226266
rect 264329 226208 264334 226264
rect 264390 226208 323532 226264
rect 264329 226206 323532 226208
rect 264329 226203 264395 226206
rect 323526 226204 323532 226206
rect 323596 226204 323602 226268
rect 243118 226068 243124 226132
rect 243188 226130 243194 226132
rect 302550 226130 302556 226132
rect 243188 226070 302556 226130
rect 243188 226068 243194 226070
rect 302550 226068 302556 226070
rect 302620 226068 302626 226132
rect 225413 225994 225479 225997
rect 227662 225994 227668 225996
rect 225413 225992 227668 225994
rect 225413 225936 225418 225992
rect 225474 225936 227668 225992
rect 225413 225934 227668 225936
rect 225413 225931 225479 225934
rect 227662 225932 227668 225934
rect 227732 225932 227738 225996
rect 248270 225932 248276 225996
rect 248340 225994 248346 225996
rect 306414 225994 306420 225996
rect 248340 225934 306420 225994
rect 248340 225932 248346 225934
rect 306414 225932 306420 225934
rect 306484 225932 306490 225996
rect 233734 225796 233740 225860
rect 233804 225858 233810 225860
rect 283925 225858 283991 225861
rect 233804 225856 283991 225858
rect 233804 225800 283930 225856
rect 283986 225800 283991 225856
rect 233804 225798 283991 225800
rect 233804 225796 233810 225798
rect 283925 225795 283991 225798
rect 163516 225662 200130 225722
rect 163516 225660 163522 225662
rect 159541 225586 159607 225589
rect 234470 225586 234476 225588
rect 159541 225584 234476 225586
rect 159541 225528 159546 225584
rect 159602 225528 234476 225584
rect 159541 225526 234476 225528
rect 159541 225523 159607 225526
rect 234470 225524 234476 225526
rect 234540 225524 234546 225588
rect 242801 225042 242867 225045
rect 243118 225042 243124 225044
rect 242801 225040 243124 225042
rect 242801 224984 242806 225040
rect 242862 224984 243124 225040
rect 242801 224982 243124 224984
rect 242801 224979 242867 224982
rect 243118 224980 243124 224982
rect 243188 224980 243194 225044
rect 240174 224906 240180 224908
rect 209730 224846 240180 224906
rect 180374 224300 180380 224364
rect 180444 224362 180450 224364
rect 208301 224362 208367 224365
rect 209730 224362 209790 224846
rect 240174 224844 240180 224846
rect 240244 224844 240250 224908
rect 300117 224906 300183 224909
rect 248370 224904 300183 224906
rect 248370 224848 300122 224904
rect 300178 224848 300183 224904
rect 248370 224846 300183 224848
rect 236913 224770 236979 224773
rect 240685 224770 240751 224773
rect 248370 224770 248430 224846
rect 300117 224843 300183 224846
rect 236913 224768 248430 224770
rect 236913 224712 236918 224768
rect 236974 224712 240690 224768
rect 240746 224712 248430 224768
rect 236913 224710 248430 224712
rect 236913 224707 236979 224710
rect 240685 224707 240751 224710
rect 261334 224708 261340 224772
rect 261404 224770 261410 224772
rect 320214 224770 320220 224772
rect 261404 224710 320220 224770
rect 261404 224708 261410 224710
rect 320214 224708 320220 224710
rect 320284 224708 320290 224772
rect 304206 224634 304212 224636
rect 248370 224574 304212 224634
rect 224217 224498 224283 224501
rect 246430 224498 246436 224500
rect 224217 224496 246436 224498
rect 224217 224440 224222 224496
rect 224278 224440 246436 224496
rect 224217 224438 246436 224440
rect 224217 224435 224283 224438
rect 246430 224436 246436 224438
rect 246500 224498 246506 224500
rect 248370 224498 248430 224574
rect 304206 224572 304212 224574
rect 304276 224572 304282 224636
rect 246500 224438 248430 224498
rect 246500 224436 246506 224438
rect 180444 224360 209790 224362
rect 180444 224304 208306 224360
rect 208362 224304 209790 224360
rect 180444 224302 209790 224304
rect 223021 224362 223087 224365
rect 251582 224362 251588 224364
rect 223021 224360 251588 224362
rect 223021 224304 223026 224360
rect 223082 224304 251588 224360
rect 223021 224302 251588 224304
rect 180444 224300 180450 224302
rect 208301 224299 208367 224302
rect 223021 224299 223087 224302
rect 251582 224300 251588 224302
rect 251652 224300 251658 224364
rect 165286 224164 165292 224228
rect 165356 224226 165362 224228
rect 225045 224226 225111 224229
rect 165356 224224 225111 224226
rect 165356 224168 225050 224224
rect 225106 224168 225111 224224
rect 165356 224166 225111 224168
rect 165356 224164 165362 224166
rect 225045 224163 225111 224166
rect 225781 224226 225847 224229
rect 246982 224226 246988 224228
rect 225781 224224 246988 224226
rect 225781 224168 225786 224224
rect 225842 224168 246988 224224
rect 225781 224166 246988 224168
rect 225781 224163 225847 224166
rect 246982 224164 246988 224166
rect 247052 224164 247058 224228
rect 205633 223546 205699 223549
rect 206645 223546 206711 223549
rect 225086 223546 225092 223548
rect 205633 223544 225092 223546
rect 205633 223488 205638 223544
rect 205694 223488 206650 223544
rect 206706 223488 225092 223544
rect 205633 223486 225092 223488
rect 205633 223483 205699 223486
rect 206645 223483 206711 223486
rect 225086 223484 225092 223486
rect 225156 223484 225162 223548
rect 263041 223546 263107 223549
rect 263174 223546 263180 223548
rect 263041 223544 263180 223546
rect 263041 223488 263046 223544
rect 263102 223488 263180 223544
rect 263041 223486 263180 223488
rect 263041 223483 263107 223486
rect 263174 223484 263180 223486
rect 263244 223546 263250 223548
rect 340873 223546 340939 223549
rect 263244 223544 340939 223546
rect 263244 223488 340878 223544
rect 340934 223488 340939 223544
rect 263244 223486 340939 223488
rect 263244 223484 263250 223486
rect 340873 223483 340939 223486
rect 260097 223410 260163 223413
rect 320766 223410 320772 223412
rect 260097 223408 320772 223410
rect 260097 223352 260102 223408
rect 260158 223352 320772 223408
rect 260097 223350 320772 223352
rect 260097 223347 260163 223350
rect 320766 223348 320772 223350
rect 320836 223348 320842 223412
rect 242249 223274 242315 223277
rect 300894 223274 300900 223276
rect 242249 223272 300900 223274
rect 242249 223216 242254 223272
rect 242310 223216 300900 223272
rect 242249 223214 300900 223216
rect 242249 223211 242315 223214
rect 300894 223212 300900 223214
rect 300964 223212 300970 223276
rect 253933 223138 253999 223141
rect 254393 223138 254459 223141
rect 314326 223138 314332 223140
rect 253933 223136 314332 223138
rect 253933 223080 253938 223136
rect 253994 223080 254398 223136
rect 254454 223080 314332 223136
rect 253933 223078 314332 223080
rect 253933 223075 253999 223078
rect 254393 223075 254459 223078
rect 314326 223076 314332 223078
rect 314396 223076 314402 223140
rect 239622 223002 239628 223004
rect 219390 222942 239628 223002
rect 178902 222804 178908 222868
rect 178972 222866 178978 222868
rect 219390 222866 219450 222942
rect 239622 222940 239628 222942
rect 239692 223002 239698 223004
rect 285213 223002 285279 223005
rect 239692 223000 285279 223002
rect 239692 222944 285218 223000
rect 285274 222944 285279 223000
rect 239692 222942 285279 222944
rect 239692 222940 239698 222942
rect 285213 222939 285279 222942
rect 178972 222806 219450 222866
rect 178972 222804 178978 222806
rect 240726 222804 240732 222868
rect 240796 222866 240802 222868
rect 278037 222866 278103 222869
rect 240796 222864 278103 222866
rect 240796 222808 278042 222864
rect 278098 222808 278103 222864
rect 240796 222806 278103 222808
rect 240796 222804 240802 222806
rect 278037 222803 278103 222806
rect 250529 222186 250595 222189
rect 251030 222186 251036 222188
rect 250529 222184 251036 222186
rect 250529 222128 250534 222184
rect 250590 222128 251036 222184
rect 250529 222126 251036 222128
rect 250529 222123 250595 222126
rect 251030 222124 251036 222126
rect 251100 222186 251106 222188
rect 315481 222186 315547 222189
rect 251100 222184 315547 222186
rect 251100 222128 315486 222184
rect 315542 222128 315547 222184
rect 251100 222126 315547 222128
rect 251100 222124 251106 222126
rect 315481 222123 315547 222126
rect 256049 222050 256115 222053
rect 256366 222050 256372 222052
rect 256049 222048 256372 222050
rect 256049 221992 256054 222048
rect 256110 221992 256372 222048
rect 256049 221990 256372 221992
rect 256049 221987 256115 221990
rect 256366 221988 256372 221990
rect 256436 222050 256442 222052
rect 308254 222050 308260 222052
rect 256436 221990 308260 222050
rect 256436 221988 256442 221990
rect 308254 221988 308260 221990
rect 308324 221988 308330 222052
rect 233182 221852 233188 221916
rect 233252 221914 233258 221916
rect 233550 221914 233556 221916
rect 233252 221854 233556 221914
rect 233252 221852 233258 221854
rect 233550 221852 233556 221854
rect 233620 221914 233626 221916
rect 280153 221914 280219 221917
rect 233620 221912 280219 221914
rect 233620 221856 280158 221912
rect 280214 221856 280219 221912
rect 233620 221854 280219 221856
rect 233620 221852 233626 221854
rect 280153 221851 280219 221854
rect 263358 221716 263364 221780
rect 263428 221778 263434 221780
rect 305821 221778 305887 221781
rect 263428 221776 305887 221778
rect 263428 221720 305826 221776
rect 305882 221720 305887 221776
rect 263428 221718 305887 221720
rect 263428 221716 263434 221718
rect 305821 221715 305887 221718
rect 180926 221580 180932 221644
rect 180996 221642 181002 221644
rect 241145 221642 241211 221645
rect 180996 221640 241211 221642
rect 180996 221584 241150 221640
rect 241206 221584 241211 221640
rect 180996 221582 241211 221584
rect 180996 221580 181002 221582
rect 241145 221579 241211 221582
rect 158161 221506 158227 221509
rect 233182 221506 233188 221508
rect 158161 221504 233188 221506
rect 158161 221448 158166 221504
rect 158222 221448 233188 221504
rect 158161 221446 233188 221448
rect 158161 221443 158227 221446
rect 233182 221444 233188 221446
rect 233252 221444 233258 221508
rect 238293 221506 238359 221509
rect 260966 221506 260972 221508
rect 238293 221504 260972 221506
rect 238293 221448 238298 221504
rect 238354 221448 260972 221504
rect 238293 221446 260972 221448
rect 238293 221443 238359 221446
rect 260966 221444 260972 221446
rect 261036 221444 261042 221508
rect 231301 221370 231367 221373
rect 264094 221370 264100 221372
rect 231301 221368 264100 221370
rect 231301 221312 231306 221368
rect 231362 221312 264100 221368
rect 231301 221310 264100 221312
rect 231301 221307 231367 221310
rect 264094 221308 264100 221310
rect 264164 221308 264170 221372
rect 230197 220826 230263 220829
rect 290549 220826 290615 220829
rect 219390 220824 290615 220826
rect 219390 220768 230202 220824
rect 230258 220768 290554 220824
rect 290610 220768 290615 220824
rect 219390 220766 290615 220768
rect 170070 220356 170076 220420
rect 170140 220418 170146 220420
rect 219390 220418 219450 220766
rect 230197 220763 230263 220766
rect 290549 220763 290615 220766
rect 230422 220628 230428 220692
rect 230492 220690 230498 220692
rect 231158 220690 231164 220692
rect 230492 220630 231164 220690
rect 230492 220628 230498 220630
rect 231158 220628 231164 220630
rect 231228 220690 231234 220692
rect 292297 220690 292363 220693
rect 231228 220688 292363 220690
rect 231228 220632 292302 220688
rect 292358 220632 292363 220688
rect 231228 220630 292363 220632
rect 231228 220628 231234 220630
rect 292297 220627 292363 220630
rect 230974 220492 230980 220556
rect 231044 220554 231050 220556
rect 231526 220554 231532 220556
rect 231044 220494 231532 220554
rect 231044 220492 231050 220494
rect 231526 220492 231532 220494
rect 231596 220554 231602 220556
rect 292113 220554 292179 220557
rect 231596 220552 292179 220554
rect 231596 220496 292118 220552
rect 292174 220496 292179 220552
rect 231596 220494 292179 220496
rect 231596 220492 231602 220494
rect 292113 220491 292179 220494
rect 170140 220358 219450 220418
rect 230473 220418 230539 220421
rect 290590 220418 290596 220420
rect 230473 220416 290596 220418
rect 230473 220360 230478 220416
rect 230534 220360 290596 220416
rect 230473 220358 290596 220360
rect 170140 220356 170146 220358
rect 230473 220355 230539 220358
rect 290590 220356 290596 220358
rect 290660 220356 290666 220420
rect 174670 220220 174676 220284
rect 174740 220282 174746 220284
rect 233601 220282 233667 220285
rect 174740 220280 233667 220282
rect 174740 220224 233606 220280
rect 233662 220224 233667 220280
rect 174740 220222 233667 220224
rect 174740 220220 174746 220222
rect 233601 220219 233667 220222
rect 256233 220282 256299 220285
rect 314878 220282 314884 220284
rect 256233 220280 314884 220282
rect 256233 220224 256238 220280
rect 256294 220224 314884 220280
rect 256233 220222 314884 220224
rect 256233 220219 256299 220222
rect 314878 220220 314884 220222
rect 314948 220220 314954 220284
rect 154113 220146 154179 220149
rect 230422 220146 230428 220148
rect 154113 220144 230428 220146
rect 154113 220088 154118 220144
rect 154174 220088 230428 220144
rect 154113 220086 230428 220088
rect 154113 220083 154179 220086
rect 230422 220084 230428 220086
rect 230492 220084 230498 220148
rect 202781 219330 202847 219333
rect 223757 219330 223823 219333
rect 202781 219328 223823 219330
rect 202781 219272 202786 219328
rect 202842 219272 223762 219328
rect 223818 219272 223823 219328
rect 202781 219270 223823 219272
rect 202781 219267 202847 219270
rect 223757 219267 223823 219270
rect 250294 219268 250300 219332
rect 250364 219330 250370 219332
rect 342345 219330 342411 219333
rect 250364 219328 342411 219330
rect 250364 219272 342350 219328
rect 342406 219272 342411 219328
rect 250364 219270 342411 219272
rect 250364 219268 250370 219270
rect 342345 219267 342411 219270
rect 255037 219194 255103 219197
rect 315062 219194 315068 219196
rect 255037 219192 315068 219194
rect 255037 219136 255042 219192
rect 255098 219136 315068 219192
rect 255037 219134 315068 219136
rect 255037 219131 255103 219134
rect 315062 219132 315068 219134
rect 315132 219132 315138 219196
rect 306966 219058 306972 219060
rect 248370 218998 306972 219058
rect 165102 218860 165108 218924
rect 165172 218922 165178 218924
rect 202781 218922 202847 218925
rect 165172 218920 202847 218922
rect 165172 218864 202786 218920
rect 202842 218864 202847 218920
rect 165172 218862 202847 218864
rect 165172 218860 165178 218862
rect 202781 218859 202847 218862
rect 236729 218922 236795 218925
rect 247534 218922 247540 218924
rect 236729 218920 247540 218922
rect 236729 218864 236734 218920
rect 236790 218864 247540 218920
rect 236729 218862 247540 218864
rect 236729 218859 236795 218862
rect 247534 218860 247540 218862
rect 247604 218922 247610 218924
rect 248370 218922 248430 218998
rect 306966 218996 306972 218998
rect 307036 218996 307042 219060
rect 580533 219058 580599 219061
rect 583520 219058 584960 219148
rect 580533 219056 584960 219058
rect 580533 219000 580538 219056
rect 580594 219000 584960 219056
rect 580533 218998 584960 219000
rect 580533 218995 580599 218998
rect 247604 218862 248430 218922
rect 247604 218860 247610 218862
rect 253422 218860 253428 218924
rect 253492 218922 253498 218924
rect 312302 218922 312308 218924
rect 253492 218862 312308 218922
rect 253492 218860 253498 218862
rect 312302 218860 312308 218862
rect 312372 218860 312378 218924
rect 583520 218908 584960 218998
rect 163630 218724 163636 218788
rect 163700 218786 163706 218788
rect 222193 218786 222259 218789
rect 163700 218784 222259 218786
rect 163700 218728 222198 218784
rect 222254 218728 222259 218784
rect 163700 218726 222259 218728
rect 163700 218724 163706 218726
rect 222193 218723 222259 218726
rect 231209 218786 231275 218789
rect 250294 218786 250300 218788
rect 231209 218784 250300 218786
rect 231209 218728 231214 218784
rect 231270 218728 250300 218784
rect 231209 218726 250300 218728
rect 231209 218723 231275 218726
rect 250294 218724 250300 218726
rect 250364 218724 250370 218788
rect 179086 218588 179092 218652
rect 179156 218650 179162 218652
rect 238886 218650 238892 218652
rect 179156 218590 238892 218650
rect 179156 218588 179162 218590
rect 238886 218588 238892 218590
rect 238956 218588 238962 218652
rect 246798 218588 246804 218652
rect 246868 218650 246874 218652
rect 280797 218650 280863 218653
rect 293309 218650 293375 218653
rect 246868 218648 293375 218650
rect 246868 218592 280802 218648
rect 280858 218592 293314 218648
rect 293370 218592 293375 218648
rect 246868 218590 293375 218592
rect 246868 218588 246874 218590
rect 280797 218587 280863 218590
rect 293309 218587 293375 218590
rect 253105 218106 253171 218109
rect 253422 218106 253428 218108
rect 253105 218104 253428 218106
rect 253105 218048 253110 218104
rect 253166 218048 253428 218104
rect 253105 218046 253428 218048
rect 253105 218043 253171 218046
rect 253422 218044 253428 218046
rect 253492 218044 253498 218108
rect 166390 217908 166396 217972
rect 166460 217970 166466 217972
rect 224953 217970 225019 217973
rect 166460 217968 225019 217970
rect 166460 217912 224958 217968
rect 225014 217912 225019 217968
rect 166460 217910 225019 217912
rect 166460 217908 166466 217910
rect 224953 217907 225019 217910
rect 167862 217772 167868 217836
rect 167932 217834 167938 217836
rect 226793 217834 226859 217837
rect 167932 217832 226859 217834
rect 167932 217776 226798 217832
rect 226854 217776 226859 217832
rect 167932 217774 226859 217776
rect 167932 217772 167938 217774
rect 226793 217771 226859 217774
rect 170438 217636 170444 217700
rect 170508 217698 170514 217700
rect 230473 217698 230539 217701
rect 170508 217696 230539 217698
rect 170508 217640 230478 217696
rect 230534 217640 230539 217696
rect 170508 217638 230539 217640
rect 170508 217636 170514 217638
rect 230473 217635 230539 217638
rect 167678 217500 167684 217564
rect 167748 217562 167754 217564
rect 227897 217562 227963 217565
rect 167748 217560 227963 217562
rect 167748 217504 227902 217560
rect 227958 217504 227963 217560
rect 167748 217502 227963 217504
rect 167748 217500 167754 217502
rect 227897 217499 227963 217502
rect 169334 217364 169340 217428
rect 169404 217426 169410 217428
rect 229645 217426 229711 217429
rect 169404 217424 229711 217426
rect 169404 217368 229650 217424
rect 229706 217368 229711 217424
rect 169404 217366 229711 217368
rect 169404 217364 169410 217366
rect 229645 217363 229711 217366
rect 170254 217228 170260 217292
rect 170324 217290 170330 217292
rect 230565 217290 230631 217293
rect 170324 217288 230631 217290
rect 170324 217232 230570 217288
rect 230626 217232 230631 217288
rect 170324 217230 230631 217232
rect 170324 217228 170330 217230
rect 230565 217227 230631 217230
rect 172094 217092 172100 217156
rect 172164 217154 172170 217156
rect 231025 217154 231091 217157
rect 172164 217152 231091 217154
rect 172164 217096 231030 217152
rect 231086 217096 231091 217152
rect 172164 217094 231091 217096
rect 172164 217092 172170 217094
rect 231025 217091 231091 217094
rect 171910 215868 171916 215932
rect 171980 215930 171986 215932
rect 231669 215930 231735 215933
rect 171980 215928 231735 215930
rect 171980 215872 231674 215928
rect 231730 215872 231735 215928
rect 171980 215870 231735 215872
rect 171980 215868 171986 215870
rect 231669 215867 231735 215870
rect -960 214978 480 215068
rect 176142 215052 176148 215116
rect 176212 215114 176218 215116
rect 232405 215114 232471 215117
rect 176212 215112 232471 215114
rect 176212 215056 232410 215112
rect 232466 215056 232471 215112
rect 176212 215054 232471 215056
rect 176212 215052 176218 215054
rect 232405 215051 232471 215054
rect 3417 214978 3483 214981
rect -960 214976 3483 214978
rect -960 214920 3422 214976
rect 3478 214920 3483 214976
rect -960 214918 3483 214920
rect -960 214828 480 214918
rect 3417 214915 3483 214918
rect 195830 214916 195836 214980
rect 195900 214978 195906 214980
rect 255037 214978 255103 214981
rect 195900 214976 255103 214978
rect 195900 214920 255042 214976
rect 255098 214920 255103 214976
rect 195900 214918 255103 214920
rect 195900 214916 195906 214918
rect 255037 214915 255103 214918
rect 191230 214780 191236 214844
rect 191300 214842 191306 214844
rect 251173 214842 251239 214845
rect 191300 214840 251239 214842
rect 191300 214784 251178 214840
rect 251234 214784 251239 214840
rect 191300 214782 251239 214784
rect 191300 214780 191306 214782
rect 251173 214779 251239 214782
rect 195646 214644 195652 214708
rect 195716 214706 195722 214708
rect 256233 214706 256299 214709
rect 195716 214704 256299 214706
rect 195716 214648 256238 214704
rect 256294 214648 256299 214704
rect 195716 214646 256299 214648
rect 195716 214644 195722 214646
rect 256233 214643 256299 214646
rect 192886 214508 192892 214572
rect 192956 214570 192962 214572
rect 253105 214570 253171 214573
rect 192956 214568 253171 214570
rect 192956 214512 253110 214568
rect 253166 214512 253171 214568
rect 192956 214510 253171 214512
rect 192956 214508 192962 214510
rect 253105 214507 253171 214510
rect 180190 213828 180196 213892
rect 180260 213890 180266 213892
rect 238845 213890 238911 213893
rect 180260 213888 238911 213890
rect 180260 213832 238850 213888
rect 238906 213832 238911 213888
rect 180260 213830 238911 213832
rect 180260 213828 180266 213830
rect 238845 213827 238911 213830
rect 177614 213692 177620 213756
rect 177684 213754 177690 213756
rect 236361 213754 236427 213757
rect 177684 213752 236427 213754
rect 177684 213696 236366 213752
rect 236422 213696 236427 213752
rect 177684 213694 236427 213696
rect 177684 213692 177690 213694
rect 236361 213691 236427 213694
rect 173382 213556 173388 213620
rect 173452 213618 173458 213620
rect 231945 213618 232011 213621
rect 173452 213616 232011 213618
rect 173452 213560 231950 213616
rect 232006 213560 232011 213616
rect 173452 213558 232011 213560
rect 173452 213556 173458 213558
rect 231945 213555 232011 213558
rect 184606 213420 184612 213484
rect 184676 213482 184682 213484
rect 243905 213482 243971 213485
rect 184676 213480 243971 213482
rect 184676 213424 243910 213480
rect 243966 213424 243971 213480
rect 184676 213422 243971 213424
rect 184676 213420 184682 213422
rect 243905 213419 243971 213422
rect 173198 213284 173204 213348
rect 173268 213346 173274 213348
rect 232773 213346 232839 213349
rect 173268 213344 232839 213346
rect 173268 213288 232778 213344
rect 232834 213288 232839 213344
rect 173268 213286 232839 213288
rect 173268 213284 173274 213286
rect 232773 213283 232839 213286
rect 174486 213148 174492 213212
rect 174556 213210 174562 213212
rect 234797 213210 234863 213213
rect 174556 213208 234863 213210
rect 174556 213152 234802 213208
rect 234858 213152 234863 213208
rect 174556 213150 234863 213152
rect 174556 213148 174562 213150
rect 234797 213147 234863 213150
rect 177798 213012 177804 213076
rect 177868 213074 177874 213076
rect 236177 213074 236243 213077
rect 177868 213072 236243 213074
rect 177868 213016 236182 213072
rect 236238 213016 236243 213072
rect 177868 213014 236243 213016
rect 177868 213012 177874 213014
rect 236177 213011 236243 213014
rect 180885 212122 180951 212125
rect 215886 212122 215892 212124
rect 180885 212120 215892 212122
rect 180885 212064 180890 212120
rect 180946 212064 215892 212120
rect 180885 212062 215892 212064
rect 180885 212059 180951 212062
rect 215886 212060 215892 212062
rect 215956 212060 215962 212124
rect 169150 211924 169156 211988
rect 169220 211986 169226 211988
rect 227713 211986 227779 211989
rect 169220 211984 227779 211986
rect 169220 211928 227718 211984
rect 227774 211928 227779 211984
rect 169220 211926 227779 211928
rect 169220 211924 169226 211926
rect 227713 211923 227779 211926
rect 180006 211788 180012 211852
rect 180076 211850 180082 211852
rect 239438 211850 239444 211852
rect 180076 211790 239444 211850
rect 180076 211788 180082 211790
rect 239438 211788 239444 211790
rect 239508 211788 239514 211852
rect 164325 211306 164391 211309
rect 164325 211304 171150 211306
rect 164325 211248 164330 211304
rect 164386 211248 171150 211304
rect 164325 211246 171150 211248
rect 164325 211243 164391 211246
rect 157793 211170 157859 211173
rect 161974 211170 161980 211172
rect 157793 211168 161980 211170
rect 157793 211112 157798 211168
rect 157854 211112 161980 211168
rect 157793 211110 161980 211112
rect 157793 211107 157859 211110
rect 161974 211108 161980 211110
rect 162044 211170 162050 211172
rect 162577 211170 162643 211173
rect 162044 211168 162643 211170
rect 162044 211112 162582 211168
rect 162638 211112 162643 211168
rect 162044 211110 162643 211112
rect 162044 211108 162050 211110
rect 162577 211107 162643 211110
rect 162710 211108 162716 211172
rect 162780 211170 162786 211172
rect 164877 211170 164943 211173
rect 165429 211170 165495 211173
rect 162780 211168 165495 211170
rect 162780 211112 164882 211168
rect 164938 211112 165434 211168
rect 165490 211112 165495 211168
rect 162780 211110 165495 211112
rect 171090 211170 171150 211246
rect 203374 211170 203380 211172
rect 171090 211110 203380 211170
rect 162780 211108 162786 211110
rect 164877 211107 164943 211110
rect 165429 211107 165495 211110
rect 203374 211108 203380 211110
rect 203444 211108 203450 211172
rect 187325 210082 187391 210085
rect 196249 210082 196315 210085
rect 187325 210080 187434 210082
rect 187325 210024 187330 210080
rect 187386 210024 187434 210080
rect 187325 210019 187434 210024
rect 164734 209612 164740 209676
rect 164804 209674 164810 209676
rect 165337 209674 165403 209677
rect 164804 209672 165403 209674
rect 164804 209616 165342 209672
rect 165398 209616 165403 209672
rect 164804 209614 165403 209616
rect 164804 209612 164810 209614
rect 165337 209611 165403 209614
rect 166206 209612 166212 209676
rect 166276 209674 166282 209676
rect 166809 209674 166875 209677
rect 166276 209672 166875 209674
rect 166276 209616 166814 209672
rect 166870 209616 166875 209672
rect 166276 209614 166875 209616
rect 166276 209612 166282 209614
rect 166809 209611 166875 209614
rect 184054 209612 184060 209676
rect 184124 209674 184130 209676
rect 184841 209674 184907 209677
rect 184124 209672 184907 209674
rect 184124 209616 184846 209672
rect 184902 209616 184907 209672
rect 184124 209614 184907 209616
rect 184124 209612 184130 209614
rect 184841 209611 184907 209614
rect 171174 209476 171180 209540
rect 171244 209538 171250 209540
rect 171961 209538 172027 209541
rect 171244 209536 172027 209538
rect 171244 209480 171966 209536
rect 172022 209480 172027 209536
rect 171244 209478 172027 209480
rect 171244 209476 171250 209478
rect 171961 209475 172027 209478
rect 183870 209476 183876 209540
rect 183940 209538 183946 209540
rect 184749 209538 184815 209541
rect 183940 209536 184815 209538
rect 183940 209480 184754 209536
rect 184810 209480 184815 209536
rect 183940 209478 184815 209480
rect 183940 209476 183946 209478
rect 184749 209475 184815 209478
rect 187374 208994 187434 210019
rect 196206 210080 196315 210082
rect 196206 210024 196254 210080
rect 196310 210024 196315 210080
rect 196206 210019 196315 210024
rect 188797 209674 188863 209677
rect 188797 209672 190470 209674
rect 188797 209616 188802 209672
rect 188858 209616 190470 209672
rect 188797 209614 190470 209616
rect 188797 209611 188863 209614
rect 188286 209476 188292 209540
rect 188356 209538 188362 209540
rect 188889 209538 188955 209541
rect 188356 209536 188955 209538
rect 188356 209480 188894 209536
rect 188950 209480 188955 209536
rect 188356 209478 188955 209480
rect 188356 209476 188362 209478
rect 188889 209475 188955 209478
rect 190410 209130 190470 209614
rect 191046 209476 191052 209540
rect 191116 209538 191122 209540
rect 191741 209538 191807 209541
rect 191116 209536 191807 209538
rect 191116 209480 191746 209536
rect 191802 209480 191807 209536
rect 191116 209478 191807 209480
rect 191116 209476 191122 209478
rect 191741 209475 191807 209478
rect 192334 209476 192340 209540
rect 192404 209538 192410 209540
rect 192937 209538 193003 209541
rect 192404 209536 193003 209538
rect 192404 209480 192942 209536
rect 192998 209480 193003 209536
rect 192404 209478 193003 209480
rect 192404 209476 192410 209478
rect 192937 209475 193003 209478
rect 193990 209476 193996 209540
rect 194060 209538 194066 209540
rect 194409 209538 194475 209541
rect 194060 209536 194475 209538
rect 194060 209480 194414 209536
rect 194470 209480 194475 209536
rect 194060 209478 194475 209480
rect 194060 209476 194066 209478
rect 194409 209475 194475 209478
rect 195462 209476 195468 209540
rect 195532 209538 195538 209540
rect 195881 209538 195947 209541
rect 195532 209536 195947 209538
rect 195532 209480 195886 209536
rect 195942 209480 195947 209536
rect 195532 209478 195947 209480
rect 195532 209476 195538 209478
rect 195881 209475 195947 209478
rect 196206 209266 196266 210019
rect 196750 209612 196756 209676
rect 196820 209674 196826 209676
rect 196985 209674 197051 209677
rect 196820 209672 197051 209674
rect 196820 209616 196990 209672
rect 197046 209616 197051 209672
rect 196820 209614 197051 209616
rect 196820 209612 196826 209614
rect 196985 209611 197051 209614
rect 197854 209612 197860 209676
rect 197924 209674 197930 209676
rect 198457 209674 198523 209677
rect 197924 209672 198523 209674
rect 197924 209616 198462 209672
rect 198518 209616 198523 209672
rect 197924 209614 198523 209616
rect 197924 209612 197930 209614
rect 198457 209611 198523 209614
rect 199326 209612 199332 209676
rect 199396 209674 199402 209676
rect 199561 209674 199627 209677
rect 199396 209672 199627 209674
rect 199396 209616 199566 209672
rect 199622 209616 199627 209672
rect 199396 209614 199627 209616
rect 199396 209612 199402 209614
rect 199561 209611 199627 209614
rect 199694 209612 199700 209676
rect 199764 209674 199770 209676
rect 199837 209674 199903 209677
rect 199764 209672 199903 209674
rect 199764 209616 199842 209672
rect 199898 209616 199903 209672
rect 199764 209614 199903 209616
rect 199764 209612 199770 209614
rect 199837 209611 199903 209614
rect 196382 209476 196388 209540
rect 196452 209538 196458 209540
rect 196893 209538 196959 209541
rect 197261 209538 197327 209541
rect 196452 209536 196959 209538
rect 196452 209480 196898 209536
rect 196954 209480 196959 209536
rect 196452 209478 196959 209480
rect 196452 209476 196458 209478
rect 196893 209475 196959 209478
rect 197126 209536 197327 209538
rect 197126 209480 197266 209536
rect 197322 209480 197327 209536
rect 197126 209478 197327 209480
rect 196566 209340 196572 209404
rect 196636 209402 196642 209404
rect 197126 209402 197186 209478
rect 197261 209475 197327 209478
rect 199510 209476 199516 209540
rect 199580 209538 199586 209540
rect 199929 209538 199995 209541
rect 199580 209536 199995 209538
rect 199580 209480 199934 209536
rect 199990 209480 199995 209536
rect 199580 209478 199995 209480
rect 199580 209476 199586 209478
rect 199929 209475 199995 209478
rect 196636 209342 197186 209402
rect 196636 209340 196642 209342
rect 580533 209266 580599 209269
rect 196206 209264 580599 209266
rect 196206 209208 580538 209264
rect 580594 209208 580599 209264
rect 196206 209206 580599 209208
rect 580533 209203 580599 209206
rect 579613 209130 579679 209133
rect 190410 209128 579679 209130
rect 190410 209072 579618 209128
rect 579674 209072 579679 209128
rect 190410 209070 579679 209072
rect 579613 209067 579679 209070
rect 580717 208994 580783 208997
rect 187374 208992 580783 208994
rect 187374 208936 580722 208992
rect 580778 208936 580783 208992
rect 187374 208934 580783 208936
rect 580717 208931 580783 208934
rect 198590 207572 198596 207636
rect 198660 207634 198666 207636
rect 256734 207634 256740 207636
rect 198660 207574 256740 207634
rect 198660 207572 198666 207574
rect 256734 207572 256740 207574
rect 256804 207572 256810 207636
rect 579613 205730 579679 205733
rect 583520 205730 584960 205820
rect 579613 205728 584960 205730
rect 579613 205672 579618 205728
rect 579674 205672 584960 205728
rect 579613 205670 584960 205672
rect 579613 205667 579679 205670
rect 583520 205580 584960 205670
rect 207749 202194 207815 202197
rect 257521 202194 257587 202197
rect 207749 202192 257587 202194
rect 207749 202136 207754 202192
rect 207810 202136 257526 202192
rect 257582 202136 257587 202192
rect 207749 202134 257587 202136
rect 207749 202131 207815 202134
rect 257521 202131 257587 202134
rect -960 201922 480 202012
rect 3325 201922 3391 201925
rect -960 201920 3391 201922
rect -960 201864 3330 201920
rect 3386 201864 3391 201920
rect -960 201862 3391 201864
rect -960 201772 480 201862
rect 3325 201859 3391 201862
rect 203374 201316 203380 201380
rect 203444 201378 203450 201380
rect 218053 201378 218119 201381
rect 218513 201378 218579 201381
rect 203444 201376 218579 201378
rect 203444 201320 218058 201376
rect 218114 201320 218518 201376
rect 218574 201320 218579 201376
rect 203444 201318 218579 201320
rect 203444 201316 203450 201318
rect 218053 201315 218119 201318
rect 218513 201315 218579 201318
rect 218053 200698 218119 200701
rect 580349 200698 580415 200701
rect 218053 200696 580415 200698
rect 218053 200640 218058 200696
rect 218114 200640 580354 200696
rect 580410 200640 580415 200696
rect 218053 200638 580415 200640
rect 218053 200635 218119 200638
rect 580349 200635 580415 200638
rect 579613 192538 579679 192541
rect 583520 192538 584960 192628
rect 579613 192536 584960 192538
rect 579613 192480 579618 192536
rect 579674 192480 584960 192536
rect 579613 192478 584960 192480
rect 579613 192475 579679 192478
rect 583520 192388 584960 192478
rect 205950 190980 205956 191044
rect 206020 191042 206026 191044
rect 264973 191042 265039 191045
rect 206020 191040 265039 191042
rect 206020 190984 264978 191040
rect 265034 190984 265039 191040
rect 206020 190982 265039 190984
rect 206020 190980 206026 190982
rect 264973 190979 265039 190982
rect -960 188866 480 188956
rect 3141 188866 3207 188869
rect -960 188864 3207 188866
rect -960 188808 3146 188864
rect 3202 188808 3207 188864
rect -960 188806 3207 188808
rect -960 188716 480 188806
rect 3141 188803 3207 188806
rect 207841 188322 207907 188325
rect 230013 188322 230079 188325
rect 207841 188320 230079 188322
rect 207841 188264 207846 188320
rect 207902 188264 230018 188320
rect 230074 188264 230079 188320
rect 207841 188262 230079 188264
rect 207841 188259 207907 188262
rect 230013 188259 230079 188262
rect 207933 184242 207999 184245
rect 231577 184242 231643 184245
rect 207933 184240 231643 184242
rect 207933 184184 207938 184240
rect 207994 184184 231582 184240
rect 231638 184184 231643 184240
rect 207933 184182 231643 184184
rect 207933 184179 207999 184182
rect 231577 184179 231643 184182
rect 207606 182820 207612 182884
rect 207676 182882 207682 182884
rect 267457 182882 267523 182885
rect 207676 182880 267523 182882
rect 207676 182824 267462 182880
rect 267518 182824 267523 182880
rect 207676 182822 267523 182824
rect 207676 182820 207682 182822
rect 267457 182819 267523 182822
rect 204110 179964 204116 180028
rect 204180 180026 204186 180028
rect 264329 180026 264395 180029
rect 204180 180024 264395 180026
rect 204180 179968 264334 180024
rect 264390 179968 264395 180024
rect 204180 179966 264395 179968
rect 204180 179964 204186 179966
rect 264329 179963 264395 179966
rect 580441 179210 580507 179213
rect 583520 179210 584960 179300
rect 580441 179208 584960 179210
rect 580441 179152 580446 179208
rect 580502 179152 584960 179208
rect 580441 179150 584960 179152
rect 580441 179147 580507 179150
rect 583520 179060 584960 179150
rect 207974 178604 207980 178668
rect 208044 178666 208050 178668
rect 267641 178666 267707 178669
rect 208044 178664 267707 178666
rect 208044 178608 267646 178664
rect 267702 178608 267707 178664
rect 208044 178606 267707 178608
rect 208044 178604 208050 178606
rect 267641 178603 267707 178606
rect 205398 177244 205404 177308
rect 205468 177306 205474 177308
rect 265709 177306 265775 177309
rect 205468 177304 265775 177306
rect 205468 177248 265714 177304
rect 265770 177248 265775 177304
rect 205468 177246 265775 177248
rect 205468 177244 205474 177246
rect 265709 177243 265775 177246
rect -960 175796 480 176036
rect 208761 173634 208827 173637
rect 209221 173634 209287 173637
rect 208761 173632 209287 173634
rect 208761 173576 208766 173632
rect 208822 173576 209226 173632
rect 209282 173576 209287 173632
rect 208761 173574 209287 173576
rect 208761 173571 208827 173574
rect 209221 173571 209287 173574
rect 208025 173498 208091 173501
rect 231393 173498 231459 173501
rect 208025 173496 231459 173498
rect 208025 173440 208030 173496
rect 208086 173440 231398 173496
rect 231454 173440 231459 173496
rect 208025 173438 231459 173440
rect 208025 173435 208091 173438
rect 231393 173435 231459 173438
rect 209078 173300 209084 173364
rect 209148 173362 209154 173364
rect 267273 173362 267339 173365
rect 209148 173360 267339 173362
rect 209148 173304 267278 173360
rect 267334 173304 267339 173360
rect 209148 173302 267339 173304
rect 209148 173300 209154 173302
rect 267273 173299 267339 173302
rect 207790 173164 207796 173228
rect 207860 173226 207866 173228
rect 267089 173226 267155 173229
rect 207860 173224 267155 173226
rect 207860 173168 267094 173224
rect 267150 173168 267155 173224
rect 207860 173166 267155 173168
rect 207860 173164 207866 173166
rect 267089 173163 267155 173166
rect 206870 171668 206876 171732
rect 206940 171730 206946 171732
rect 266445 171730 266511 171733
rect 206940 171728 266511 171730
rect 206940 171672 266450 171728
rect 266506 171672 266511 171728
rect 206940 171670 266511 171672
rect 206940 171668 206946 171670
rect 266445 171667 266511 171670
rect 207565 170370 207631 170373
rect 224401 170370 224467 170373
rect 207565 170368 224467 170370
rect 207565 170312 207570 170368
rect 207626 170312 224406 170368
rect 224462 170312 224467 170368
rect 207565 170310 224467 170312
rect 207565 170307 207631 170310
rect 224401 170307 224467 170310
rect 209262 169084 209268 169148
rect 209332 169146 209338 169148
rect 266997 169146 267063 169149
rect 209332 169144 267063 169146
rect 209332 169088 267002 169144
rect 267058 169088 267063 169144
rect 209332 169086 267063 169088
rect 209332 169084 209338 169086
rect 266997 169083 267063 169086
rect 205214 168948 205220 169012
rect 205284 169010 205290 169012
rect 263910 169010 263916 169012
rect 205284 168950 263916 169010
rect 205284 168948 205290 168950
rect 263910 168948 263916 168950
rect 263980 168948 263986 169012
rect 207749 166426 207815 166429
rect 208117 166426 208183 166429
rect 265617 166426 265683 166429
rect 207749 166424 208183 166426
rect 207749 166368 207754 166424
rect 207810 166368 208122 166424
rect 208178 166368 208183 166424
rect 207749 166366 208183 166368
rect 207749 166363 207815 166366
rect 208117 166363 208183 166366
rect 208350 166424 265683 166426
rect 208350 166368 265622 166424
rect 265678 166368 265683 166424
rect 208350 166366 265683 166368
rect 207657 166154 207723 166157
rect 208350 166154 208410 166366
rect 265617 166363 265683 166366
rect 263685 166290 263751 166293
rect 207657 166152 208410 166154
rect 207657 166096 207662 166152
rect 207718 166096 208410 166152
rect 207657 166094 208410 166096
rect 209730 166288 263751 166290
rect 209730 166232 263690 166288
rect 263746 166232 263751 166288
rect 209730 166230 263751 166232
rect 207657 166091 207723 166094
rect 204662 165956 204668 166020
rect 204732 166018 204738 166020
rect 209730 166018 209790 166230
rect 263685 166227 263751 166230
rect 204732 165958 209790 166018
rect 204732 165956 204738 165958
rect 580717 165882 580783 165885
rect 583520 165882 584960 165972
rect 580717 165880 584960 165882
rect 580717 165824 580722 165880
rect 580778 165824 584960 165880
rect 580717 165822 584960 165824
rect 580717 165819 580783 165822
rect 583520 165732 584960 165822
rect 203926 165004 203932 165068
rect 203996 165066 204002 165068
rect 263593 165066 263659 165069
rect 203996 165064 263659 165066
rect 203996 165008 263598 165064
rect 263654 165008 263659 165064
rect 203996 165006 263659 165008
rect 203996 165004 204002 165006
rect 263593 165003 263659 165006
rect 206502 164868 206508 164932
rect 206572 164930 206578 164932
rect 267549 164930 267615 164933
rect 206572 164928 267615 164930
rect 206572 164872 267554 164928
rect 267610 164872 267615 164928
rect 206572 164870 267615 164872
rect 206572 164868 206578 164870
rect 267549 164867 267615 164870
rect 203558 163508 203564 163572
rect 203628 163570 203634 163572
rect 263041 163570 263107 163573
rect 203628 163568 263107 163570
rect 203628 163512 263046 163568
rect 263102 163512 263107 163568
rect 203628 163510 263107 163512
rect 203628 163508 203634 163510
rect 263041 163507 263107 163510
rect 204846 163372 204852 163436
rect 204916 163434 204922 163436
rect 266169 163434 266235 163437
rect 204916 163432 266235 163434
rect 204916 163376 266174 163432
rect 266230 163376 266235 163432
rect 204916 163374 266235 163376
rect 204916 163372 204922 163374
rect 266169 163371 266235 163374
rect -960 162890 480 162980
rect 3325 162890 3391 162893
rect -960 162888 3391 162890
rect -960 162832 3330 162888
rect 3386 162832 3391 162888
rect -960 162830 3391 162832
rect -960 162740 480 162830
rect 3325 162827 3391 162830
rect 206686 162148 206692 162212
rect 206756 162210 206762 162212
rect 223665 162210 223731 162213
rect 206756 162208 223731 162210
rect 206756 162152 223670 162208
rect 223726 162152 223731 162208
rect 206756 162150 223731 162152
rect 206756 162148 206762 162150
rect 223665 162147 223731 162150
rect 203190 162012 203196 162076
rect 203260 162074 203266 162076
rect 260281 162074 260347 162077
rect 203260 162072 260347 162074
rect 203260 162016 260286 162072
rect 260342 162016 260347 162072
rect 203260 162014 260347 162016
rect 203260 162012 203266 162014
rect 260281 162011 260347 162014
rect 161105 161938 161171 161941
rect 170990 161938 170996 161940
rect 161105 161936 170996 161938
rect 161105 161880 161110 161936
rect 161166 161880 170996 161936
rect 161105 161878 170996 161880
rect 161105 161875 161171 161878
rect 170990 161876 170996 161878
rect 171060 161876 171066 161940
rect 201350 161876 201356 161940
rect 201420 161938 201426 161940
rect 261845 161938 261911 161941
rect 201420 161936 261911 161938
rect 201420 161880 261850 161936
rect 261906 161880 261911 161936
rect 201420 161878 261911 161880
rect 201420 161876 201426 161878
rect 261845 161875 261911 161878
rect 169150 161740 169156 161804
rect 169220 161802 169226 161804
rect 228081 161802 228147 161805
rect 169220 161800 228147 161802
rect 169220 161744 228086 161800
rect 228142 161744 228147 161800
rect 169220 161742 228147 161744
rect 169220 161740 169226 161742
rect 228081 161739 228147 161742
rect 208209 161394 208275 161397
rect 260189 161394 260255 161397
rect 208209 161392 260255 161394
rect 208209 161336 208214 161392
rect 208270 161336 260194 161392
rect 260250 161336 260255 161392
rect 208209 161334 260255 161336
rect 208209 161331 208275 161334
rect 260189 161331 260255 161334
rect 197854 161196 197860 161260
rect 197924 161258 197930 161260
rect 257429 161258 257495 161261
rect 197924 161256 257495 161258
rect 197924 161200 257434 161256
rect 257490 161200 257495 161256
rect 197924 161198 257495 161200
rect 197924 161196 197930 161198
rect 257429 161195 257495 161198
rect 249425 161122 249491 161125
rect 195930 161120 249491 161122
rect 195930 161064 249430 161120
rect 249486 161064 249491 161120
rect 195930 161062 249491 161064
rect 164366 160788 164372 160852
rect 164436 160850 164442 160852
rect 165102 160850 165108 160852
rect 164436 160790 165108 160850
rect 164436 160788 164442 160790
rect 165102 160788 165108 160790
rect 165172 160788 165178 160852
rect 186814 160850 186820 160852
rect 176610 160790 186820 160850
rect 167126 160652 167132 160716
rect 167196 160714 167202 160716
rect 175958 160714 175964 160716
rect 167196 160654 175964 160714
rect 167196 160652 167202 160654
rect 175958 160652 175964 160654
rect 176028 160652 176034 160716
rect 159357 160578 159423 160581
rect 167310 160578 167316 160580
rect 159357 160576 167316 160578
rect 159357 160520 159362 160576
rect 159418 160520 167316 160576
rect 159357 160518 167316 160520
rect 159357 160515 159423 160518
rect 167310 160516 167316 160518
rect 167380 160516 167386 160580
rect 156965 160442 157031 160445
rect 166022 160442 166028 160444
rect 156965 160440 166028 160442
rect 156965 160384 156970 160440
rect 157026 160384 166028 160440
rect 156965 160382 166028 160384
rect 156965 160379 157031 160382
rect 166022 160380 166028 160382
rect 166092 160380 166098 160444
rect 158253 160306 158319 160309
rect 158253 160304 168298 160306
rect 158253 160248 158258 160304
rect 158314 160248 168298 160304
rect 158253 160246 168298 160248
rect 158253 160243 158319 160246
rect 155309 160170 155375 160173
rect 155309 160168 164756 160170
rect 155309 160112 155314 160168
rect 155370 160112 164756 160168
rect 155309 160110 164756 160112
rect 155309 160107 155375 160110
rect 156689 160034 156755 160037
rect 156689 160032 164112 160034
rect 156689 159976 156694 160032
rect 156750 159976 164112 160032
rect 156689 159974 164112 159976
rect 156689 159971 156755 159974
rect 155677 159898 155743 159901
rect 162117 159898 162183 159901
rect 163037 159898 163103 159901
rect 155677 159896 163103 159898
rect 155677 159840 155682 159896
rect 155738 159840 162122 159896
rect 162178 159840 163042 159896
rect 163098 159840 163103 159896
rect 155677 159838 163103 159840
rect 155677 159835 155743 159838
rect 162117 159835 162183 159838
rect 163037 159835 163103 159838
rect 163405 159898 163471 159901
rect 163589 159898 163655 159901
rect 163814 159898 163820 159900
rect 163405 159896 163514 159898
rect 163405 159840 163410 159896
rect 163466 159840 163514 159896
rect 163405 159835 163514 159840
rect 163589 159896 163820 159898
rect 163589 159840 163594 159896
rect 163650 159840 163820 159896
rect 163589 159838 163820 159840
rect 163589 159835 163655 159838
rect 163814 159836 163820 159838
rect 163884 159836 163890 159900
rect 160553 159762 160619 159765
rect 162945 159762 163011 159765
rect 160553 159760 163011 159762
rect 160553 159704 160558 159760
rect 160614 159704 162950 159760
rect 163006 159704 163011 159760
rect 160553 159702 163011 159704
rect 160553 159699 160619 159702
rect 162945 159699 163011 159702
rect 163262 159700 163268 159764
rect 163332 159762 163338 159764
rect 163454 159762 163514 159835
rect 163332 159702 163514 159762
rect 163332 159700 163338 159702
rect 152549 159626 152615 159629
rect 152917 159626 152983 159629
rect 163405 159626 163471 159629
rect 163630 159626 163636 159628
rect 152549 159624 157350 159626
rect 152549 159568 152554 159624
rect 152610 159568 152922 159624
rect 152978 159568 157350 159624
rect 152549 159566 157350 159568
rect 152549 159563 152615 159566
rect 152917 159563 152983 159566
rect 157290 159490 157350 159566
rect 163405 159624 163636 159626
rect 163405 159568 163410 159624
rect 163466 159568 163636 159624
rect 163405 159566 163636 159568
rect 163405 159563 163471 159566
rect 163630 159564 163636 159566
rect 163700 159564 163706 159628
rect 164052 159626 164112 159974
rect 164696 159935 164756 160110
rect 167126 160108 167132 160172
rect 167196 160108 167202 160172
rect 166758 160034 166764 160036
rect 165662 159974 166764 160034
rect 164693 159930 164759 159935
rect 164233 159898 164299 159901
rect 164366 159898 164372 159900
rect 164233 159896 164372 159898
rect 164233 159840 164238 159896
rect 164294 159840 164372 159896
rect 164233 159838 164372 159840
rect 164233 159835 164299 159838
rect 164366 159836 164372 159838
rect 164436 159836 164442 159900
rect 164693 159874 164698 159930
rect 164754 159874 164759 159930
rect 165662 159901 165722 159974
rect 166758 159972 166764 159974
rect 166828 159972 166834 160036
rect 167134 159901 167194 160108
rect 168238 159901 168298 160246
rect 176610 160170 176670 160790
rect 186814 160788 186820 160790
rect 186884 160788 186890 160852
rect 181478 160244 181484 160308
rect 181548 160244 181554 160308
rect 169710 160110 176670 160170
rect 169334 159972 169340 160036
rect 169404 160034 169410 160036
rect 169404 159974 169586 160034
rect 169404 159972 169410 159974
rect 169526 159901 169586 159974
rect 164693 159869 164759 159874
rect 164918 159836 164924 159900
rect 164988 159898 164994 159900
rect 165337 159898 165403 159901
rect 164988 159896 165403 159898
rect 164988 159840 165342 159896
rect 165398 159840 165403 159896
rect 164988 159838 165403 159840
rect 164988 159836 164994 159838
rect 165337 159835 165403 159838
rect 165613 159896 165722 159901
rect 165613 159840 165618 159896
rect 165674 159840 165722 159896
rect 165613 159838 165722 159840
rect 166257 159898 166323 159901
rect 166390 159898 166396 159900
rect 166257 159896 166396 159898
rect 166257 159840 166262 159896
rect 166318 159840 166396 159896
rect 166257 159838 166396 159840
rect 165613 159835 165679 159838
rect 166257 159835 166323 159838
rect 166390 159836 166396 159838
rect 166460 159836 166466 159900
rect 166574 159836 166580 159900
rect 166644 159898 166650 159900
rect 166717 159898 166783 159901
rect 166644 159896 166783 159898
rect 166644 159840 166722 159896
rect 166778 159840 166783 159896
rect 166644 159838 166783 159840
rect 167134 159896 167243 159901
rect 167134 159840 167182 159896
rect 167238 159840 167243 159896
rect 167134 159838 167243 159840
rect 166644 159836 166650 159838
rect 166717 159835 166783 159838
rect 167177 159835 167243 159838
rect 167310 159836 167316 159900
rect 167380 159898 167386 159900
rect 167453 159898 167519 159901
rect 167380 159896 167519 159898
rect 167380 159840 167458 159896
rect 167514 159840 167519 159896
rect 167380 159838 167519 159840
rect 167380 159836 167386 159838
rect 167453 159835 167519 159838
rect 167637 159898 167703 159901
rect 167862 159898 167868 159900
rect 167637 159896 167868 159898
rect 167637 159840 167642 159896
rect 167698 159840 167868 159896
rect 167637 159838 167868 159840
rect 167637 159835 167703 159838
rect 167862 159836 167868 159838
rect 167932 159836 167938 159900
rect 168238 159896 168347 159901
rect 168238 159840 168286 159896
rect 168342 159840 168347 159896
rect 168238 159838 168347 159840
rect 168281 159835 168347 159838
rect 168741 159898 168807 159901
rect 168966 159898 168972 159900
rect 168741 159896 168972 159898
rect 168741 159840 168746 159896
rect 168802 159840 168972 159896
rect 168741 159838 168972 159840
rect 168741 159835 168807 159838
rect 168966 159836 168972 159838
rect 169036 159836 169042 159900
rect 169201 159898 169267 159901
rect 169201 159896 169402 159898
rect 169201 159840 169206 159896
rect 169262 159840 169402 159896
rect 169201 159838 169402 159840
rect 169201 159835 169267 159838
rect 165153 159762 165219 159765
rect 165521 159764 165587 159765
rect 165286 159762 165292 159764
rect 165153 159760 165292 159762
rect 165153 159704 165158 159760
rect 165214 159704 165292 159760
rect 165153 159702 165292 159704
rect 165153 159699 165219 159702
rect 165286 159700 165292 159702
rect 165356 159700 165362 159764
rect 165470 159700 165476 159764
rect 165540 159762 165587 159764
rect 166165 159764 166231 159765
rect 166165 159762 166212 159764
rect 165540 159760 165632 159762
rect 165582 159704 165632 159760
rect 165540 159702 165632 159704
rect 166084 159760 166212 159762
rect 166276 159762 166282 159764
rect 166809 159762 166875 159765
rect 166276 159760 166875 159762
rect 166084 159704 166170 159760
rect 166276 159704 166814 159760
rect 166870 159704 166875 159760
rect 166084 159702 166212 159704
rect 165540 159700 165587 159702
rect 165521 159699 165587 159700
rect 166165 159700 166212 159702
rect 166276 159702 166875 159704
rect 166276 159700 166282 159702
rect 166165 159699 166231 159700
rect 166809 159699 166875 159702
rect 167678 159700 167684 159764
rect 167748 159762 167754 159764
rect 168189 159762 168255 159765
rect 167748 159760 168255 159762
rect 167748 159704 168194 159760
rect 168250 159704 168255 159760
rect 167748 159702 168255 159704
rect 167748 159700 167754 159702
rect 168189 159699 168255 159702
rect 168465 159762 168531 159765
rect 168598 159762 168604 159764
rect 168465 159760 168604 159762
rect 168465 159704 168470 159760
rect 168526 159704 168604 159760
rect 168465 159702 168604 159704
rect 168465 159699 168531 159702
rect 168598 159700 168604 159702
rect 168668 159700 168674 159764
rect 169017 159762 169083 159765
rect 169150 159762 169156 159764
rect 169017 159760 169156 159762
rect 169017 159704 169022 159760
rect 169078 159704 169156 159760
rect 169017 159702 169156 159704
rect 169017 159699 169083 159702
rect 169150 159700 169156 159702
rect 169220 159700 169226 159764
rect 169342 159762 169402 159838
rect 169477 159896 169586 159901
rect 169477 159840 169482 159896
rect 169538 159840 169586 159896
rect 169477 159838 169586 159840
rect 169477 159835 169543 159838
rect 169518 159762 169524 159764
rect 169342 159702 169524 159762
rect 169518 159700 169524 159702
rect 169588 159700 169594 159764
rect 165613 159626 165679 159629
rect 164052 159624 165679 159626
rect 164052 159568 165618 159624
rect 165674 159568 165679 159624
rect 164052 159566 165679 159568
rect 165613 159563 165679 159566
rect 166022 159564 166028 159628
rect 166092 159626 166098 159628
rect 166349 159626 166415 159629
rect 166092 159624 166415 159626
rect 166092 159568 166354 159624
rect 166410 159568 166415 159624
rect 166092 159566 166415 159568
rect 166092 159564 166098 159566
rect 166349 159563 166415 159566
rect 167913 159626 167979 159629
rect 168230 159626 168236 159628
rect 167913 159624 168236 159626
rect 167913 159568 167918 159624
rect 167974 159568 168236 159624
rect 167913 159566 168236 159568
rect 167913 159563 167979 159566
rect 168230 159564 168236 159566
rect 168300 159564 168306 159628
rect 169293 159626 169359 159629
rect 169710 159626 169770 160110
rect 172278 160034 172284 160036
rect 171366 159974 172284 160034
rect 170070 159836 170076 159900
rect 170140 159898 170146 159900
rect 170397 159898 170463 159901
rect 170140 159896 170463 159898
rect 170140 159840 170402 159896
rect 170458 159840 170463 159896
rect 170140 159838 170463 159840
rect 170140 159836 170146 159838
rect 170397 159835 170463 159838
rect 170622 159836 170628 159900
rect 170692 159898 170698 159900
rect 170949 159898 171015 159901
rect 170692 159896 171015 159898
rect 170692 159840 170954 159896
rect 171010 159840 171015 159896
rect 170692 159838 171015 159840
rect 170692 159836 170698 159838
rect 170949 159835 171015 159838
rect 171133 159898 171199 159901
rect 171366 159898 171426 159974
rect 172278 159972 172284 159974
rect 172348 159972 172354 160036
rect 173198 160034 173204 160036
rect 172470 159974 173204 160034
rect 171133 159896 171426 159898
rect 171133 159840 171138 159896
rect 171194 159840 171426 159896
rect 171133 159838 171426 159840
rect 171777 159898 171843 159901
rect 171910 159898 171916 159900
rect 171777 159896 171916 159898
rect 171777 159840 171782 159896
rect 171838 159840 171916 159896
rect 171777 159838 171916 159840
rect 171133 159835 171199 159838
rect 171777 159835 171843 159838
rect 171910 159836 171916 159838
rect 171980 159836 171986 159900
rect 172470 159898 172530 159974
rect 173198 159972 173204 159974
rect 173268 159972 173274 160036
rect 175038 160034 175044 160036
rect 174126 159974 175044 160034
rect 172605 159898 172671 159901
rect 172881 159900 172947 159901
rect 172830 159898 172836 159900
rect 172470 159896 172671 159898
rect 172470 159840 172610 159896
rect 172666 159840 172671 159896
rect 172470 159838 172671 159840
rect 172754 159838 172836 159898
rect 172900 159898 172947 159900
rect 173382 159898 173388 159900
rect 172900 159896 173388 159898
rect 172942 159840 173388 159896
rect 170581 159764 170647 159765
rect 170581 159762 170628 159764
rect 170536 159760 170628 159762
rect 170536 159704 170586 159760
rect 170536 159702 170628 159704
rect 170581 159700 170628 159702
rect 170692 159700 170698 159764
rect 170765 159762 170831 159765
rect 170949 159764 171015 159765
rect 170765 159760 170874 159762
rect 170765 159704 170770 159760
rect 170826 159704 170874 159760
rect 170581 159699 170647 159700
rect 170765 159699 170874 159704
rect 170949 159760 170996 159764
rect 171060 159762 171066 159764
rect 171409 159762 171475 159765
rect 172094 159762 172100 159764
rect 170949 159704 170954 159760
rect 170949 159700 170996 159704
rect 171060 159702 171106 159762
rect 171409 159760 172100 159762
rect 171409 159704 171414 159760
rect 171470 159704 172100 159760
rect 171409 159702 172100 159704
rect 171060 159700 171066 159702
rect 170949 159699 171015 159700
rect 171409 159699 171475 159702
rect 172094 159700 172100 159702
rect 172164 159700 172170 159764
rect 172470 159762 172530 159838
rect 172605 159835 172671 159838
rect 172830 159836 172836 159838
rect 172900 159838 173388 159840
rect 172900 159836 172947 159838
rect 173382 159836 173388 159838
rect 173452 159836 173458 159900
rect 173566 159836 173572 159900
rect 173636 159898 173642 159900
rect 173709 159898 173775 159901
rect 173636 159896 173775 159898
rect 173636 159840 173714 159896
rect 173770 159840 173775 159896
rect 173636 159838 173775 159840
rect 173636 159836 173642 159838
rect 172881 159835 172947 159836
rect 173709 159835 173775 159838
rect 173985 159898 174051 159901
rect 174126 159898 174186 159974
rect 175038 159972 175044 159974
rect 175108 159972 175114 160036
rect 180742 159972 180748 160036
rect 180812 160034 180818 160036
rect 181486 160034 181546 160244
rect 195930 160170 195990 161062
rect 249425 161059 249491 161062
rect 257613 160986 257679 160989
rect 201358 160984 257679 160986
rect 201358 160928 257618 160984
rect 257674 160928 257679 160984
rect 201358 160926 257679 160928
rect 201358 160442 201418 160926
rect 257613 160923 257679 160926
rect 203374 160788 203380 160852
rect 203444 160850 203450 160852
rect 273621 160850 273687 160853
rect 203444 160848 273687 160850
rect 203444 160792 273626 160848
rect 273682 160792 273687 160848
rect 203444 160790 273687 160792
rect 203444 160788 203450 160790
rect 273621 160787 273687 160790
rect 208393 160714 208459 160717
rect 277485 160714 277551 160717
rect 208393 160712 277551 160714
rect 208393 160656 208398 160712
rect 208454 160656 277490 160712
rect 277546 160656 277551 160712
rect 208393 160654 277551 160656
rect 208393 160651 208459 160654
rect 277485 160651 277551 160654
rect 202822 160516 202828 160580
rect 202892 160578 202898 160580
rect 245694 160578 245700 160580
rect 202892 160518 245700 160578
rect 202892 160516 202898 160518
rect 245694 160516 245700 160518
rect 245764 160516 245770 160580
rect 197678 160382 201418 160442
rect 197678 160170 197738 160382
rect 208209 160306 208275 160309
rect 202462 160304 208275 160306
rect 202462 160248 208214 160304
rect 208270 160248 208275 160304
rect 202462 160246 208275 160248
rect 189582 160110 195990 160170
rect 197126 160110 197738 160170
rect 182582 160034 182588 160036
rect 180812 159974 182098 160034
rect 180812 159972 180818 159974
rect 173985 159896 174186 159898
rect 173985 159840 173990 159896
rect 174046 159840 174186 159896
rect 173985 159838 174186 159840
rect 174537 159898 174603 159901
rect 174854 159898 174860 159900
rect 174537 159896 174860 159898
rect 174537 159840 174542 159896
rect 174598 159840 174860 159896
rect 174537 159838 174860 159840
rect 173985 159835 174051 159838
rect 174537 159835 174603 159838
rect 174854 159836 174860 159838
rect 174924 159836 174930 159900
rect 175917 159898 175983 159901
rect 176510 159898 176516 159900
rect 175917 159896 176516 159898
rect 175917 159840 175922 159896
rect 175978 159840 176516 159896
rect 175917 159838 176516 159840
rect 175917 159835 175983 159838
rect 176510 159836 176516 159838
rect 176580 159836 176586 159900
rect 177297 159898 177363 159901
rect 178953 159900 179019 159901
rect 180057 159900 180123 159901
rect 177614 159898 177620 159900
rect 177297 159896 177620 159898
rect 177297 159840 177302 159896
rect 177358 159840 177620 159896
rect 177297 159838 177620 159840
rect 177297 159835 177363 159838
rect 177614 159836 177620 159838
rect 177684 159836 177690 159900
rect 178902 159836 178908 159900
rect 178972 159898 179019 159900
rect 178972 159896 179064 159898
rect 179014 159840 179064 159896
rect 178972 159838 179064 159840
rect 178972 159836 179019 159838
rect 180006 159836 180012 159900
rect 180076 159898 180123 159900
rect 180333 159900 180399 159901
rect 180609 159900 180675 159901
rect 180333 159898 180380 159900
rect 180076 159896 180168 159898
rect 180118 159840 180168 159896
rect 180076 159838 180168 159840
rect 180288 159896 180380 159898
rect 180288 159840 180338 159896
rect 180288 159838 180380 159840
rect 180076 159836 180123 159838
rect 178953 159835 179019 159836
rect 180057 159835 180123 159836
rect 180333 159836 180380 159838
rect 180444 159836 180450 159900
rect 180558 159836 180564 159900
rect 180628 159898 180675 159900
rect 180628 159896 180720 159898
rect 180670 159840 180720 159896
rect 180628 159838 180720 159840
rect 180628 159836 180675 159838
rect 180926 159836 180932 159900
rect 180996 159898 181002 159900
rect 181161 159898 181227 159901
rect 180996 159896 181227 159898
rect 180996 159840 181166 159896
rect 181222 159840 181227 159896
rect 180996 159838 181227 159840
rect 180996 159836 181002 159838
rect 180333 159835 180399 159836
rect 180609 159835 180675 159836
rect 181161 159835 181227 159838
rect 181294 159836 181300 159900
rect 181364 159898 181370 159900
rect 181897 159898 181963 159901
rect 181364 159896 181963 159898
rect 181364 159840 181902 159896
rect 181958 159840 181963 159896
rect 181364 159838 181963 159840
rect 181364 159836 181370 159838
rect 181897 159835 181963 159838
rect 172697 159762 172763 159765
rect 172470 159760 172763 159762
rect 172470 159704 172702 159760
rect 172758 159704 172763 159760
rect 172470 159702 172763 159704
rect 172697 159699 172763 159702
rect 173014 159700 173020 159764
rect 173084 159762 173090 159764
rect 173249 159762 173315 159765
rect 173433 159764 173499 159765
rect 173084 159760 173315 159762
rect 173084 159704 173254 159760
rect 173310 159704 173315 159760
rect 173084 159702 173315 159704
rect 173084 159700 173090 159702
rect 173249 159699 173315 159702
rect 173382 159700 173388 159764
rect 173452 159762 173499 159764
rect 173750 159762 173756 159764
rect 173452 159760 173756 159762
rect 173494 159704 173756 159760
rect 173452 159702 173756 159704
rect 173452 159700 173499 159702
rect 173750 159700 173756 159702
rect 173820 159700 173826 159764
rect 174261 159762 174327 159765
rect 174670 159762 174676 159764
rect 173942 159760 174676 159762
rect 173942 159704 174266 159760
rect 174322 159704 174676 159760
rect 173942 159702 174676 159704
rect 173433 159699 173499 159700
rect 169293 159624 169770 159626
rect 169293 159568 169298 159624
rect 169354 159568 169770 159624
rect 169293 159566 169770 159568
rect 169293 159563 169359 159566
rect 170438 159564 170444 159628
rect 170508 159626 170514 159628
rect 170814 159626 170874 159699
rect 173942 159629 174002 159702
rect 174261 159699 174327 159702
rect 174670 159700 174676 159702
rect 174740 159700 174746 159764
rect 174813 159762 174879 159765
rect 176878 159762 176884 159764
rect 174813 159760 176884 159762
rect 174813 159704 174818 159760
rect 174874 159704 176884 159760
rect 174813 159702 176884 159704
rect 174813 159699 174879 159702
rect 176878 159700 176884 159702
rect 176948 159700 176954 159764
rect 177021 159762 177087 159765
rect 177798 159762 177804 159764
rect 177021 159760 177804 159762
rect 177021 159704 177026 159760
rect 177082 159704 177804 159760
rect 177021 159702 177804 159704
rect 177021 159699 177087 159702
rect 177798 159700 177804 159702
rect 177868 159700 177874 159764
rect 179086 159700 179092 159764
rect 179156 159762 179162 159764
rect 179229 159762 179295 159765
rect 179156 159760 179295 159762
rect 179156 159704 179234 159760
rect 179290 159704 179295 159760
rect 179156 159702 179295 159704
rect 179156 159700 179162 159702
rect 179229 159699 179295 159702
rect 179781 159762 179847 159765
rect 180190 159762 180196 159764
rect 179781 159760 180196 159762
rect 179781 159704 179786 159760
rect 179842 159704 180196 159760
rect 179781 159702 180196 159704
rect 179781 159699 179847 159702
rect 180190 159700 180196 159702
rect 180260 159762 180266 159764
rect 180333 159762 180399 159765
rect 180260 159760 180399 159762
rect 180260 159704 180338 159760
rect 180394 159704 180399 159760
rect 180260 159702 180399 159704
rect 180260 159700 180266 159702
rect 180333 159699 180399 159702
rect 180885 159762 180951 159765
rect 181478 159762 181484 159764
rect 180885 159760 181484 159762
rect 180885 159704 180890 159760
rect 180946 159704 181484 159760
rect 180885 159702 181484 159704
rect 180885 159699 180951 159702
rect 181478 159700 181484 159702
rect 181548 159700 181554 159764
rect 181713 159762 181779 159765
rect 182038 159762 182098 159974
rect 182406 159974 182588 160034
rect 182265 159898 182331 159901
rect 182406 159898 182466 159974
rect 182582 159972 182588 159974
rect 182652 160034 182658 160036
rect 183134 160034 183140 160036
rect 182652 159974 183140 160034
rect 182652 159972 182658 159974
rect 183134 159972 183140 159974
rect 183204 159972 183210 160036
rect 184606 160034 184612 160036
rect 184062 159974 184612 160034
rect 182817 159900 182883 159901
rect 182265 159896 182466 159898
rect 182265 159840 182270 159896
rect 182326 159840 182466 159896
rect 182265 159838 182466 159840
rect 182265 159835 182331 159838
rect 182766 159836 182772 159900
rect 182836 159898 182883 159900
rect 183277 159900 183343 159901
rect 183277 159898 183324 159900
rect 182836 159896 182928 159898
rect 182878 159840 182928 159896
rect 182836 159838 182928 159840
rect 183232 159896 183324 159898
rect 183232 159840 183282 159896
rect 183232 159838 183324 159840
rect 182836 159836 182883 159838
rect 182817 159835 182883 159836
rect 183277 159836 183324 159838
rect 183388 159836 183394 159900
rect 183921 159898 183987 159901
rect 184062 159898 184122 159974
rect 184606 159972 184612 159974
rect 184676 159972 184682 160036
rect 183921 159896 184122 159898
rect 183921 159840 183926 159896
rect 183982 159840 184122 159896
rect 183921 159838 184122 159840
rect 184197 159898 184263 159901
rect 188337 159900 188403 159901
rect 184422 159898 184428 159900
rect 184197 159896 184428 159898
rect 184197 159840 184202 159896
rect 184258 159840 184428 159896
rect 184197 159838 184428 159840
rect 183277 159835 183343 159836
rect 183921 159835 183987 159838
rect 184197 159835 184263 159838
rect 184422 159836 184428 159838
rect 184492 159836 184498 159900
rect 188286 159836 188292 159900
rect 188356 159898 188403 159900
rect 188356 159896 188448 159898
rect 188398 159840 188448 159896
rect 188356 159838 188448 159840
rect 188356 159836 188403 159838
rect 188337 159835 188403 159836
rect 189582 159765 189642 160110
rect 190862 159972 190868 160036
rect 190932 160034 190938 160036
rect 190932 159974 191298 160034
rect 190932 159972 190938 159974
rect 189717 159898 189783 159901
rect 190310 159898 190316 159900
rect 189717 159896 190316 159898
rect 189717 159840 189722 159896
rect 189778 159840 190316 159896
rect 189717 159838 190316 159840
rect 189717 159835 189783 159838
rect 190310 159836 190316 159838
rect 190380 159836 190386 159900
rect 190821 159898 190887 159901
rect 191046 159898 191052 159900
rect 190821 159896 191052 159898
rect 190821 159840 190826 159896
rect 190882 159840 191052 159896
rect 190821 159838 191052 159840
rect 190821 159835 190887 159838
rect 191046 159836 191052 159838
rect 191116 159836 191122 159900
rect 191238 159898 191298 159974
rect 196382 159972 196388 160036
rect 196452 160034 196458 160036
rect 196452 159974 196818 160034
rect 196452 159972 196458 159974
rect 191373 159898 191439 159901
rect 191238 159896 191439 159898
rect 191238 159840 191378 159896
rect 191434 159840 191439 159896
rect 191238 159838 191439 159840
rect 191373 159835 191439 159838
rect 192334 159836 192340 159900
rect 192404 159898 192410 159900
rect 192477 159898 192543 159901
rect 192404 159896 192543 159898
rect 192404 159840 192482 159896
rect 192538 159840 192543 159896
rect 192404 159838 192543 159840
rect 192404 159836 192410 159838
rect 192477 159835 192543 159838
rect 192753 159898 192819 159901
rect 192886 159898 192892 159900
rect 192753 159896 192892 159898
rect 192753 159840 192758 159896
rect 192814 159840 192892 159896
rect 192753 159838 192892 159840
rect 192753 159835 192819 159838
rect 192886 159836 192892 159838
rect 192956 159836 192962 159900
rect 193581 159898 193647 159901
rect 193806 159898 193812 159900
rect 193581 159896 193812 159898
rect 193581 159840 193586 159896
rect 193642 159840 193812 159896
rect 193581 159838 193812 159840
rect 193581 159835 193647 159838
rect 193806 159836 193812 159838
rect 193876 159836 193882 159900
rect 194174 159836 194180 159900
rect 194244 159898 194250 159900
rect 194409 159898 194475 159901
rect 194244 159896 194475 159898
rect 194244 159840 194414 159896
rect 194470 159840 194475 159896
rect 194244 159838 194475 159840
rect 194244 159836 194250 159838
rect 194409 159835 194475 159838
rect 194961 159898 195027 159901
rect 195094 159898 195100 159900
rect 194961 159896 195100 159898
rect 194961 159840 194966 159896
rect 195022 159840 195100 159896
rect 194961 159838 195100 159840
rect 194961 159835 195027 159838
rect 195094 159836 195100 159838
rect 195164 159898 195170 159900
rect 195462 159898 195468 159900
rect 195164 159838 195468 159898
rect 195164 159836 195170 159838
rect 195462 159836 195468 159838
rect 195532 159836 195538 159900
rect 195646 159836 195652 159900
rect 195716 159898 195722 159900
rect 195789 159898 195855 159901
rect 195716 159896 195855 159898
rect 195716 159840 195794 159896
rect 195850 159840 195855 159896
rect 195716 159838 195855 159840
rect 195716 159836 195722 159838
rect 195789 159835 195855 159838
rect 196341 159898 196407 159901
rect 196566 159898 196572 159900
rect 196341 159896 196572 159898
rect 196341 159840 196346 159896
rect 196402 159840 196572 159896
rect 196341 159838 196572 159840
rect 196341 159835 196407 159838
rect 196566 159836 196572 159838
rect 196636 159836 196642 159900
rect 196758 159898 196818 159974
rect 197126 159901 197186 160110
rect 197854 160108 197860 160172
rect 197924 160108 197930 160172
rect 199694 160170 199700 160172
rect 198966 160110 199700 160170
rect 197862 159901 197922 160108
rect 196893 159898 196959 159901
rect 196758 159896 196959 159898
rect 196758 159840 196898 159896
rect 196954 159840 196959 159896
rect 196758 159838 196959 159840
rect 197126 159896 197235 159901
rect 197126 159840 197174 159896
rect 197230 159840 197235 159896
rect 197126 159838 197235 159840
rect 197862 159896 197971 159901
rect 197862 159840 197910 159896
rect 197966 159840 197971 159896
rect 197862 159838 197971 159840
rect 196893 159835 196959 159838
rect 197169 159835 197235 159838
rect 197905 159835 197971 159838
rect 198406 159836 198412 159900
rect 198476 159898 198482 159900
rect 198549 159898 198615 159901
rect 198476 159896 198615 159898
rect 198476 159840 198554 159896
rect 198610 159840 198615 159896
rect 198476 159838 198615 159840
rect 198476 159836 198482 159838
rect 198549 159835 198615 159838
rect 198825 159898 198891 159901
rect 198966 159898 199026 160110
rect 199694 160108 199700 160110
rect 199764 160108 199770 160172
rect 199510 160034 199516 160036
rect 199150 159974 199516 160034
rect 199150 159901 199210 159974
rect 199510 159972 199516 159974
rect 199580 159972 199586 160036
rect 198825 159896 199026 159898
rect 198825 159840 198830 159896
rect 198886 159840 199026 159896
rect 198825 159838 199026 159840
rect 199101 159896 199210 159901
rect 199377 159900 199443 159901
rect 199101 159840 199106 159896
rect 199162 159840 199210 159896
rect 199101 159838 199210 159840
rect 198825 159835 198891 159838
rect 199101 159835 199167 159838
rect 199326 159836 199332 159900
rect 199396 159898 199443 159900
rect 201309 159900 201375 159901
rect 201309 159898 201356 159900
rect 199396 159896 199488 159898
rect 199438 159840 199488 159896
rect 199396 159838 199488 159840
rect 201264 159896 201356 159898
rect 201264 159840 201314 159896
rect 201264 159838 201356 159840
rect 199396 159836 199443 159838
rect 199377 159835 199443 159836
rect 201309 159836 201356 159838
rect 201420 159836 201426 159900
rect 202321 159898 202387 159901
rect 202462 159898 202522 160246
rect 208209 160243 208275 160246
rect 208393 160170 208459 160173
rect 205774 160168 208459 160170
rect 205774 160112 208398 160168
rect 208454 160112 208459 160168
rect 205774 160110 208459 160112
rect 203517 159900 203583 159901
rect 203517 159898 203564 159900
rect 202321 159896 202522 159898
rect 202321 159840 202326 159896
rect 202382 159840 202522 159896
rect 202321 159838 202522 159840
rect 203472 159896 203564 159898
rect 203472 159840 203522 159896
rect 203472 159838 203564 159840
rect 201309 159835 201375 159836
rect 202321 159835 202387 159838
rect 203517 159836 203564 159838
rect 203628 159836 203634 159900
rect 203793 159898 203859 159901
rect 204110 159898 204116 159900
rect 203793 159896 204116 159898
rect 203793 159840 203798 159896
rect 203854 159840 204116 159896
rect 203793 159838 204116 159840
rect 203517 159835 203583 159836
rect 203793 159835 203859 159838
rect 204110 159836 204116 159838
rect 204180 159836 204186 159900
rect 204621 159898 204687 159901
rect 205030 159898 205036 159900
rect 204621 159896 205036 159898
rect 204621 159840 204626 159896
rect 204682 159840 205036 159896
rect 204621 159838 205036 159840
rect 204621 159835 204687 159838
rect 205030 159836 205036 159838
rect 205100 159836 205106 159900
rect 205173 159898 205239 159901
rect 205398 159898 205404 159900
rect 205173 159896 205404 159898
rect 205173 159840 205178 159896
rect 205234 159840 205404 159896
rect 205173 159838 205404 159840
rect 205173 159835 205239 159838
rect 205398 159836 205404 159838
rect 205468 159836 205474 159900
rect 183369 159764 183435 159765
rect 181713 159760 182098 159762
rect 181713 159704 181718 159760
rect 181774 159704 182098 159760
rect 181713 159702 182098 159704
rect 181713 159699 181779 159702
rect 182950 159700 182956 159764
rect 183020 159762 183026 159764
rect 183318 159762 183324 159764
rect 183020 159702 183324 159762
rect 183388 159760 183435 159764
rect 183430 159704 183435 159760
rect 183020 159700 183026 159702
rect 183318 159700 183324 159702
rect 183388 159700 183435 159704
rect 184054 159700 184060 159764
rect 184124 159762 184130 159764
rect 184473 159762 184539 159765
rect 184124 159760 184539 159762
rect 184124 159704 184478 159760
rect 184534 159704 184539 159760
rect 184124 159702 184539 159704
rect 189582 159760 189691 159765
rect 189582 159704 189630 159760
rect 189686 159704 189691 159760
rect 189582 159702 189691 159704
rect 184124 159700 184130 159702
rect 183369 159699 183435 159700
rect 184473 159699 184539 159702
rect 189625 159699 189691 159702
rect 191097 159762 191163 159765
rect 191414 159762 191420 159764
rect 191097 159760 191420 159762
rect 191097 159704 191102 159760
rect 191158 159704 191420 159760
rect 191097 159702 191420 159704
rect 191097 159699 191163 159702
rect 191414 159700 191420 159702
rect 191484 159700 191490 159764
rect 192201 159762 192267 159765
rect 192702 159762 192708 159764
rect 192201 159760 192708 159762
rect 192201 159704 192206 159760
rect 192262 159704 192708 159760
rect 192201 159702 192708 159704
rect 192201 159699 192267 159702
rect 192702 159700 192708 159702
rect 192772 159700 192778 159764
rect 195237 159762 195303 159765
rect 195830 159762 195836 159764
rect 195237 159760 195836 159762
rect 195237 159704 195242 159760
rect 195298 159704 195836 159760
rect 195237 159702 195836 159704
rect 195237 159699 195303 159702
rect 195830 159700 195836 159702
rect 195900 159700 195906 159764
rect 196617 159762 196683 159765
rect 196934 159762 196940 159764
rect 196617 159760 196940 159762
rect 196617 159704 196622 159760
rect 196678 159704 196940 159760
rect 196617 159702 196940 159704
rect 196617 159699 196683 159702
rect 196934 159700 196940 159702
rect 197004 159700 197010 159764
rect 197997 159762 198063 159765
rect 198590 159762 198596 159764
rect 197997 159760 198596 159762
rect 197997 159704 198002 159760
rect 198058 159704 198596 159760
rect 197997 159702 198596 159704
rect 197997 159699 198063 159702
rect 198590 159700 198596 159702
rect 198660 159700 198666 159764
rect 199377 159762 199443 159765
rect 203425 159764 203491 159765
rect 203190 159762 203196 159764
rect 199377 159760 203196 159762
rect 199377 159704 199382 159760
rect 199438 159704 203196 159760
rect 199377 159702 203196 159704
rect 199377 159699 199443 159702
rect 203190 159700 203196 159702
rect 203260 159700 203266 159764
rect 203374 159700 203380 159764
rect 203444 159762 203491 159764
rect 203444 159760 203536 159762
rect 203486 159704 203536 159760
rect 203444 159702 203536 159704
rect 203444 159700 203491 159702
rect 203926 159700 203932 159764
rect 203996 159762 204002 159764
rect 204069 159762 204135 159765
rect 203996 159760 204135 159762
rect 203996 159704 204074 159760
rect 204130 159704 204135 159760
rect 203996 159702 204135 159704
rect 203996 159700 204002 159702
rect 203425 159699 203491 159700
rect 204069 159699 204135 159702
rect 204846 159700 204852 159764
rect 204916 159762 204922 159764
rect 205449 159762 205515 159765
rect 204916 159760 205515 159762
rect 204916 159704 205454 159760
rect 205510 159704 205515 159760
rect 204916 159702 205515 159704
rect 204916 159700 204922 159702
rect 205449 159699 205515 159702
rect 205633 159762 205699 159765
rect 205774 159762 205834 160110
rect 208393 160107 208459 160110
rect 205950 159836 205956 159900
rect 206020 159898 206026 159900
rect 206277 159898 206343 159901
rect 206553 159900 206619 159901
rect 206020 159896 206343 159898
rect 206020 159840 206282 159896
rect 206338 159840 206343 159896
rect 206020 159838 206343 159840
rect 206020 159836 206026 159838
rect 206277 159835 206343 159838
rect 206502 159836 206508 159900
rect 206572 159898 206619 159900
rect 206829 159900 206895 159901
rect 206572 159896 206664 159898
rect 206614 159840 206664 159896
rect 206572 159838 206664 159840
rect 206829 159896 206876 159900
rect 206940 159898 206946 159900
rect 207289 159898 207355 159901
rect 207790 159898 207796 159900
rect 206829 159840 206834 159896
rect 206572 159836 206619 159838
rect 206553 159835 206619 159836
rect 206829 159836 206876 159840
rect 206940 159838 206986 159898
rect 207289 159896 207796 159898
rect 207289 159840 207294 159896
rect 207350 159840 207796 159896
rect 207289 159838 207796 159840
rect 206940 159836 206946 159838
rect 206829 159835 206895 159836
rect 207289 159835 207355 159838
rect 207790 159836 207796 159838
rect 207860 159836 207866 159900
rect 205633 159760 205834 159762
rect 205633 159704 205638 159760
rect 205694 159704 205834 159760
rect 205633 159702 205834 159704
rect 207381 159762 207447 159765
rect 207606 159762 207612 159764
rect 207381 159760 207612 159762
rect 207381 159704 207386 159760
rect 207442 159704 207612 159760
rect 207381 159702 207612 159704
rect 205633 159699 205699 159702
rect 207381 159699 207447 159702
rect 207606 159700 207612 159702
rect 207676 159700 207682 159764
rect 170508 159566 170874 159626
rect 171225 159626 171291 159629
rect 171501 159626 171567 159629
rect 171225 159624 171567 159626
rect 171225 159568 171230 159624
rect 171286 159568 171506 159624
rect 171562 159568 171567 159624
rect 171225 159566 171567 159568
rect 170508 159564 170514 159566
rect 171225 159563 171291 159566
rect 171501 159563 171567 159566
rect 172513 159626 172579 159629
rect 172646 159626 172652 159628
rect 172513 159624 172652 159626
rect 172513 159568 172518 159624
rect 172574 159568 172652 159624
rect 172513 159566 172652 159568
rect 172513 159563 172579 159566
rect 172646 159564 172652 159566
rect 172716 159626 172722 159628
rect 173433 159626 173499 159629
rect 172716 159624 173499 159626
rect 172716 159568 173438 159624
rect 173494 159568 173499 159624
rect 172716 159566 173499 159568
rect 172716 159564 172722 159566
rect 173433 159563 173499 159566
rect 173893 159624 174002 159629
rect 173893 159568 173898 159624
rect 173954 159568 174002 159624
rect 173893 159566 174002 159568
rect 173893 159563 173959 159566
rect 174486 159564 174492 159628
rect 174556 159626 174562 159628
rect 175089 159626 175155 159629
rect 209129 159626 209195 159629
rect 174556 159624 175155 159626
rect 174556 159568 175094 159624
rect 175150 159568 175155 159624
rect 174556 159566 175155 159568
rect 174556 159564 174562 159566
rect 175089 159563 175155 159566
rect 176610 159624 209195 159626
rect 176610 159568 209134 159624
rect 209190 159568 209195 159624
rect 176610 159566 209195 159568
rect 169385 159490 169451 159493
rect 157290 159488 169451 159490
rect 157290 159432 169390 159488
rect 169446 159432 169451 159488
rect 157290 159430 169451 159432
rect 169385 159427 169451 159430
rect 169845 159490 169911 159493
rect 175774 159490 175780 159492
rect 169845 159488 175780 159490
rect 169845 159432 169850 159488
rect 169906 159432 175780 159488
rect 169845 159430 175780 159432
rect 169845 159427 169911 159430
rect 175774 159428 175780 159430
rect 175844 159428 175850 159492
rect 156873 159354 156939 159357
rect 167177 159354 167243 159357
rect 156873 159352 167243 159354
rect 156873 159296 156878 159352
rect 156934 159296 167182 159352
rect 167238 159296 167243 159352
rect 156873 159294 167243 159296
rect 156873 159291 156939 159294
rect 167177 159291 167243 159294
rect 168598 159292 168604 159356
rect 168668 159354 168674 159356
rect 176610 159354 176670 159566
rect 209129 159563 209195 159566
rect 183870 159428 183876 159492
rect 183940 159490 183946 159492
rect 184749 159490 184815 159493
rect 183940 159488 184815 159490
rect 183940 159432 184754 159488
rect 184810 159432 184815 159488
rect 183940 159430 184815 159432
rect 183940 159428 183946 159430
rect 184749 159427 184815 159430
rect 191230 159428 191236 159492
rect 191300 159490 191306 159492
rect 191649 159490 191715 159493
rect 191300 159488 191715 159490
rect 191300 159432 191654 159488
rect 191710 159432 191715 159488
rect 191300 159430 191715 159432
rect 191300 159428 191306 159430
rect 191649 159427 191715 159430
rect 197905 159490 197971 159493
rect 202321 159490 202387 159493
rect 197905 159488 202387 159490
rect 197905 159432 197910 159488
rect 197966 159432 202326 159488
rect 202382 159432 202387 159488
rect 197905 159430 202387 159432
rect 197905 159427 197971 159430
rect 202321 159427 202387 159430
rect 202873 159490 202939 159493
rect 238569 159490 238635 159493
rect 202873 159488 238635 159490
rect 202873 159432 202878 159488
rect 202934 159432 238574 159488
rect 238630 159432 238635 159488
rect 202873 159430 238635 159432
rect 202873 159427 202939 159430
rect 238569 159427 238635 159430
rect 168668 159294 176670 159354
rect 168668 159292 168674 159294
rect 176878 159292 176884 159356
rect 176948 159354 176954 159356
rect 185158 159354 185164 159356
rect 176948 159294 185164 159354
rect 176948 159292 176954 159294
rect 185158 159292 185164 159294
rect 185228 159292 185234 159356
rect 200113 159354 200179 159357
rect 239765 159354 239831 159357
rect 200113 159352 239831 159354
rect 200113 159296 200118 159352
rect 200174 159296 239770 159352
rect 239826 159296 239831 159352
rect 200113 159294 239831 159296
rect 200113 159291 200179 159294
rect 239765 159291 239831 159294
rect 158713 159218 158779 159221
rect 166441 159218 166507 159221
rect 224033 159218 224099 159221
rect 158713 159216 166274 159218
rect 158713 159160 158718 159216
rect 158774 159160 166274 159216
rect 158713 159158 166274 159160
rect 158713 159155 158779 159158
rect 162945 159082 163011 159085
rect 165889 159084 165955 159085
rect 162945 159080 165354 159082
rect 162945 159024 162950 159080
rect 163006 159024 165354 159080
rect 162945 159022 165354 159024
rect 162945 159019 163011 159022
rect 151261 158946 151327 158949
rect 151537 158946 151603 158949
rect 165153 158946 165219 158949
rect 151261 158944 165219 158946
rect 151261 158888 151266 158944
rect 151322 158888 151542 158944
rect 151598 158888 165158 158944
rect 165214 158888 165219 158944
rect 151261 158886 165219 158888
rect 151261 158883 151327 158886
rect 151537 158883 151603 158886
rect 165153 158883 165219 158886
rect 156781 158810 156847 158813
rect 164325 158810 164391 158813
rect 156781 158808 164391 158810
rect 156781 158752 156786 158808
rect 156842 158752 164330 158808
rect 164386 158752 164391 158808
rect 156781 158750 164391 158752
rect 165294 158810 165354 159022
rect 165838 159020 165844 159084
rect 165908 159082 165955 159084
rect 166214 159082 166274 159158
rect 166441 159216 224099 159218
rect 166441 159160 166446 159216
rect 166502 159160 224038 159216
rect 224094 159160 224099 159216
rect 166441 159158 224099 159160
rect 166441 159155 166507 159158
rect 224033 159155 224099 159158
rect 174721 159082 174787 159085
rect 165908 159080 166000 159082
rect 165950 159024 166000 159080
rect 165908 159022 166000 159024
rect 166214 159080 174787 159082
rect 166214 159024 174726 159080
rect 174782 159024 174787 159080
rect 166214 159022 174787 159024
rect 165908 159020 165955 159022
rect 165889 159019 165955 159020
rect 174721 159019 174787 159022
rect 188429 159082 188495 159085
rect 201401 159084 201467 159085
rect 201350 159082 201356 159084
rect 188429 159080 188538 159082
rect 188429 159024 188434 159080
rect 188490 159024 188538 159080
rect 188429 159019 188538 159024
rect 201310 159022 201356 159082
rect 201420 159080 201467 159084
rect 201462 159024 201467 159080
rect 201350 159020 201356 159022
rect 201420 159020 201467 159024
rect 204662 159020 204668 159084
rect 204732 159082 204738 159084
rect 204897 159082 204963 159085
rect 204732 159080 204963 159082
rect 204732 159024 204902 159080
rect 204958 159024 204963 159080
rect 204732 159022 204963 159024
rect 204732 159020 204738 159022
rect 201401 159019 201467 159020
rect 204897 159019 204963 159022
rect 206185 159082 206251 159085
rect 278957 159082 279023 159085
rect 206185 159080 279023 159082
rect 206185 159024 206190 159080
rect 206246 159024 278962 159080
rect 279018 159024 279023 159080
rect 206185 159022 279023 159024
rect 206185 159019 206251 159022
rect 278957 159019 279023 159022
rect 165613 158946 165679 158949
rect 166349 158946 166415 158949
rect 168557 158948 168623 158949
rect 168557 158946 168604 158948
rect 165613 158944 166415 158946
rect 165613 158888 165618 158944
rect 165674 158888 166354 158944
rect 166410 158888 166415 158944
rect 165613 158886 166415 158888
rect 168512 158944 168604 158946
rect 168512 158888 168562 158944
rect 168512 158886 168604 158888
rect 165613 158883 165679 158886
rect 166349 158883 166415 158886
rect 168557 158884 168604 158886
rect 168668 158884 168674 158948
rect 170581 158946 170647 158949
rect 173014 158946 173020 158948
rect 170581 158944 173020 158946
rect 170581 158888 170586 158944
rect 170642 158888 173020 158944
rect 170581 158886 173020 158888
rect 168557 158883 168623 158884
rect 170581 158883 170647 158886
rect 173014 158884 173020 158886
rect 173084 158884 173090 158948
rect 173433 158946 173499 158949
rect 181897 158946 181963 158949
rect 173433 158944 181963 158946
rect 173433 158888 173438 158944
rect 173494 158888 181902 158944
rect 181958 158888 181963 158944
rect 173433 158886 181963 158888
rect 173433 158883 173499 158886
rect 181897 158883 181963 158886
rect 188478 158813 188538 159019
rect 190545 158946 190611 158949
rect 200389 158946 200455 158949
rect 273529 158946 273595 158949
rect 190545 158944 190746 158946
rect 190545 158888 190550 158944
rect 190606 158888 190746 158944
rect 190545 158886 190746 158888
rect 190545 158883 190611 158886
rect 174813 158810 174879 158813
rect 165294 158808 174879 158810
rect 165294 158752 174818 158808
rect 174874 158752 174879 158808
rect 165294 158750 174879 158752
rect 156781 158747 156847 158750
rect 164325 158747 164391 158750
rect 174813 158747 174879 158750
rect 176377 158810 176443 158813
rect 176510 158810 176516 158812
rect 176377 158808 176516 158810
rect 176377 158752 176382 158808
rect 176438 158752 176516 158808
rect 176377 158750 176516 158752
rect 176377 158747 176443 158750
rect 176510 158748 176516 158750
rect 176580 158748 176586 158812
rect 186313 158810 186379 158813
rect 186446 158810 186452 158812
rect 186313 158808 186452 158810
rect 186313 158752 186318 158808
rect 186374 158752 186452 158808
rect 186313 158750 186452 158752
rect 186313 158747 186379 158750
rect 186446 158748 186452 158750
rect 186516 158748 186522 158812
rect 188429 158808 188538 158813
rect 188429 158752 188434 158808
rect 188490 158752 188538 158808
rect 188429 158750 188538 158752
rect 188429 158747 188495 158750
rect 159449 158674 159515 158677
rect 160001 158674 160067 158677
rect 159449 158672 160067 158674
rect 159449 158616 159454 158672
rect 159510 158616 160006 158672
rect 160062 158616 160067 158672
rect 159449 158614 160067 158616
rect 159449 158611 159515 158614
rect 160001 158611 160067 158614
rect 163037 158676 163103 158677
rect 163037 158672 163084 158676
rect 163148 158674 163154 158676
rect 164693 158674 164759 158677
rect 164918 158674 164924 158676
rect 163037 158616 163042 158672
rect 163037 158612 163084 158616
rect 163148 158614 163194 158674
rect 164693 158672 164924 158674
rect 164693 158616 164698 158672
rect 164754 158616 164924 158672
rect 164693 158614 164924 158616
rect 163148 158612 163154 158614
rect 163037 158611 163103 158612
rect 164693 158611 164759 158614
rect 164918 158612 164924 158614
rect 164988 158612 164994 158676
rect 165705 158674 165771 158677
rect 166257 158674 166323 158677
rect 166809 158676 166875 158677
rect 165705 158672 166323 158674
rect 165705 158616 165710 158672
rect 165766 158616 166262 158672
rect 166318 158616 166323 158672
rect 165705 158614 166323 158616
rect 165705 158611 165771 158614
rect 166257 158611 166323 158614
rect 166758 158612 166764 158676
rect 166828 158674 166875 158676
rect 167085 158674 167151 158677
rect 168046 158674 168052 158676
rect 166828 158672 166920 158674
rect 166870 158616 166920 158672
rect 166828 158614 166920 158616
rect 167085 158672 168052 158674
rect 167085 158616 167090 158672
rect 167146 158616 168052 158672
rect 167085 158614 168052 158616
rect 166828 158612 166875 158614
rect 166809 158611 166875 158612
rect 167085 158611 167151 158614
rect 168046 158612 168052 158614
rect 168116 158612 168122 158676
rect 168414 158612 168420 158676
rect 168484 158674 168490 158676
rect 168649 158674 168715 158677
rect 168484 158672 168715 158674
rect 168484 158616 168654 158672
rect 168710 158616 168715 158672
rect 168484 158614 168715 158616
rect 168484 158612 168490 158614
rect 168649 158611 168715 158614
rect 169385 158674 169451 158677
rect 169518 158674 169524 158676
rect 169385 158672 169524 158674
rect 169385 158616 169390 158672
rect 169446 158616 169524 158672
rect 169385 158614 169524 158616
rect 169385 158611 169451 158614
rect 169518 158612 169524 158614
rect 169588 158612 169594 158676
rect 170070 158612 170076 158676
rect 170140 158674 170146 158676
rect 171041 158674 171107 158677
rect 170140 158672 171107 158674
rect 170140 158616 171046 158672
rect 171102 158616 171107 158672
rect 170140 158614 171107 158616
rect 170140 158612 170146 158614
rect 171041 158611 171107 158614
rect 171317 158674 171383 158677
rect 171542 158674 171548 158676
rect 171317 158672 171548 158674
rect 171317 158616 171322 158672
rect 171378 158616 171548 158672
rect 171317 158614 171548 158616
rect 171317 158611 171383 158614
rect 171542 158612 171548 158614
rect 171612 158612 171618 158676
rect 171910 158612 171916 158676
rect 171980 158674 171986 158676
rect 172145 158674 172211 158677
rect 171980 158672 172211 158674
rect 171980 158616 172150 158672
rect 172206 158616 172211 158672
rect 171980 158614 172211 158616
rect 171980 158612 171986 158614
rect 172145 158611 172211 158614
rect 173065 158674 173131 158677
rect 174629 158676 174695 158677
rect 173566 158674 173572 158676
rect 173065 158672 173572 158674
rect 173065 158616 173070 158672
rect 173126 158616 173572 158672
rect 173065 158614 173572 158616
rect 173065 158611 173131 158614
rect 173566 158612 173572 158614
rect 173636 158612 173642 158676
rect 174629 158672 174676 158676
rect 174740 158674 174746 158676
rect 175641 158674 175707 158677
rect 176142 158674 176148 158676
rect 174629 158616 174634 158672
rect 174629 158612 174676 158616
rect 174740 158614 174786 158674
rect 175641 158672 176148 158674
rect 175641 158616 175646 158672
rect 175702 158616 176148 158672
rect 175641 158614 176148 158616
rect 174740 158612 174746 158614
rect 174629 158611 174695 158612
rect 175641 158611 175707 158614
rect 176142 158612 176148 158614
rect 176212 158612 176218 158676
rect 176377 158674 176443 158677
rect 177573 158676 177639 158677
rect 176377 158672 177498 158674
rect 176377 158616 176382 158672
rect 176438 158616 177498 158672
rect 176377 158614 177498 158616
rect 176377 158611 176443 158614
rect 157885 158538 157951 158541
rect 163446 158538 163452 158540
rect 157885 158536 163452 158538
rect 157885 158480 157890 158536
rect 157946 158480 163452 158536
rect 157885 158478 163452 158480
rect 157885 158475 157951 158478
rect 163446 158476 163452 158478
rect 163516 158538 163522 158540
rect 163865 158538 163931 158541
rect 163516 158536 163931 158538
rect 163516 158480 163870 158536
rect 163926 158480 163931 158536
rect 163516 158478 163931 158480
rect 163516 158476 163522 158478
rect 163865 158475 163931 158478
rect 164601 158538 164667 158541
rect 164877 158538 164943 158541
rect 164601 158536 164943 158538
rect 164601 158480 164606 158536
rect 164662 158480 164882 158536
rect 164938 158480 164943 158536
rect 164601 158478 164943 158480
rect 164601 158475 164667 158478
rect 164877 158475 164943 158478
rect 165153 158538 165219 158541
rect 165286 158538 165292 158540
rect 165153 158536 165292 158538
rect 165153 158480 165158 158536
rect 165214 158480 165292 158536
rect 165153 158478 165292 158480
rect 165153 158475 165219 158478
rect 165286 158476 165292 158478
rect 165356 158476 165362 158540
rect 165654 158476 165660 158540
rect 165724 158538 165730 158540
rect 166717 158538 166783 158541
rect 177438 158538 177498 158614
rect 177573 158672 177620 158676
rect 177684 158674 177690 158676
rect 177573 158616 177578 158672
rect 177573 158612 177620 158616
rect 177684 158614 177730 158674
rect 177684 158612 177690 158614
rect 178718 158612 178724 158676
rect 178788 158674 178794 158676
rect 179137 158674 179203 158677
rect 178788 158672 179203 158674
rect 178788 158616 179142 158672
rect 179198 158616 179203 158672
rect 178788 158614 179203 158616
rect 178788 158612 178794 158614
rect 177573 158611 177639 158612
rect 179137 158611 179203 158614
rect 179822 158612 179828 158676
rect 179892 158674 179898 158676
rect 180558 158674 180564 158676
rect 179892 158614 180564 158674
rect 179892 158612 179898 158614
rect 180558 158612 180564 158614
rect 180628 158612 180634 158676
rect 181110 158612 181116 158676
rect 181180 158674 181186 158676
rect 181437 158674 181503 158677
rect 181180 158672 181503 158674
rect 181180 158616 181442 158672
rect 181498 158616 181503 158672
rect 181180 158614 181503 158616
rect 181180 158612 181186 158614
rect 181437 158611 181503 158614
rect 182541 158674 182607 158677
rect 183093 158676 183159 158677
rect 185025 158676 185091 158677
rect 182950 158674 182956 158676
rect 182541 158672 182956 158674
rect 182541 158616 182546 158672
rect 182602 158616 182956 158672
rect 182541 158614 182956 158616
rect 182541 158611 182607 158614
rect 182950 158612 182956 158614
rect 183020 158612 183026 158676
rect 183093 158672 183140 158676
rect 183204 158674 183210 158676
rect 184974 158674 184980 158676
rect 183093 158616 183098 158672
rect 183093 158612 183140 158616
rect 183204 158614 183250 158674
rect 184934 158614 184980 158674
rect 185044 158672 185091 158676
rect 185086 158616 185091 158672
rect 183204 158612 183210 158614
rect 184974 158612 184980 158614
rect 185044 158612 185091 158616
rect 185158 158612 185164 158676
rect 185228 158674 185234 158676
rect 185853 158674 185919 158677
rect 185228 158672 185919 158674
rect 185228 158616 185858 158672
rect 185914 158616 185919 158672
rect 185228 158614 185919 158616
rect 185228 158612 185234 158614
rect 183093 158611 183159 158612
rect 185025 158611 185091 158612
rect 185853 158611 185919 158614
rect 186681 158674 186747 158677
rect 186998 158674 187004 158676
rect 186681 158672 187004 158674
rect 186681 158616 186686 158672
rect 186742 158616 187004 158672
rect 186681 158614 187004 158616
rect 186681 158611 186747 158614
rect 186998 158612 187004 158614
rect 187068 158612 187074 158676
rect 187233 158674 187299 158677
rect 187509 158676 187575 158677
rect 187366 158674 187372 158676
rect 187233 158672 187372 158674
rect 187233 158616 187238 158672
rect 187294 158616 187372 158672
rect 187233 158614 187372 158616
rect 187233 158611 187299 158614
rect 187366 158612 187372 158614
rect 187436 158612 187442 158676
rect 187509 158672 187556 158676
rect 187620 158674 187626 158676
rect 188061 158674 188127 158677
rect 188613 158676 188679 158677
rect 188470 158674 188476 158676
rect 187509 158616 187514 158672
rect 187509 158612 187556 158616
rect 187620 158614 187666 158674
rect 188061 158672 188476 158674
rect 188061 158616 188066 158672
rect 188122 158616 188476 158672
rect 188061 158614 188476 158616
rect 187620 158612 187626 158614
rect 187509 158611 187575 158612
rect 188061 158611 188127 158614
rect 188470 158612 188476 158614
rect 188540 158612 188546 158676
rect 188613 158672 188660 158676
rect 188724 158674 188730 158676
rect 189165 158674 189231 158677
rect 189993 158676 190059 158677
rect 189758 158674 189764 158676
rect 188613 158616 188618 158672
rect 188613 158612 188660 158616
rect 188724 158614 188770 158674
rect 189165 158672 189764 158674
rect 189165 158616 189170 158672
rect 189226 158616 189764 158672
rect 189165 158614 189764 158616
rect 188724 158612 188730 158614
rect 188613 158611 188679 158612
rect 189165 158611 189231 158614
rect 189758 158612 189764 158614
rect 189828 158612 189834 158676
rect 189942 158674 189948 158676
rect 189902 158614 189948 158674
rect 190012 158672 190059 158676
rect 190054 158616 190059 158672
rect 189942 158612 189948 158614
rect 190012 158612 190059 158616
rect 190126 158612 190132 158676
rect 190196 158674 190202 158676
rect 190269 158674 190335 158677
rect 190196 158672 190335 158674
rect 190196 158616 190274 158672
rect 190330 158616 190335 158672
rect 190196 158614 190335 158616
rect 190686 158674 190746 158886
rect 200389 158944 273595 158946
rect 200389 158888 200394 158944
rect 200450 158888 273534 158944
rect 273590 158888 273595 158944
rect 200389 158886 273595 158888
rect 200389 158883 200455 158886
rect 273529 158883 273595 158886
rect 201493 158810 201559 158813
rect 276197 158810 276263 158813
rect 201493 158808 276263 158810
rect 201493 158752 201498 158808
rect 201554 158752 276202 158808
rect 276258 158752 276263 158808
rect 201493 158750 276263 158752
rect 201493 158747 201559 158750
rect 276197 158747 276263 158750
rect 191230 158674 191236 158676
rect 190686 158614 191236 158674
rect 190196 158612 190202 158614
rect 189993 158611 190059 158612
rect 190269 158611 190335 158614
rect 191230 158612 191236 158614
rect 191300 158612 191306 158676
rect 191925 158674 191991 158677
rect 192702 158674 192708 158676
rect 191925 158672 192708 158674
rect 191925 158616 191930 158672
rect 191986 158616 192708 158672
rect 191925 158614 192708 158616
rect 191925 158611 191991 158614
rect 192702 158612 192708 158614
rect 192772 158612 192778 158676
rect 192886 158612 192892 158676
rect 192956 158674 192962 158676
rect 193029 158674 193095 158677
rect 192956 158672 193095 158674
rect 192956 158616 193034 158672
rect 193090 158616 193095 158672
rect 192956 158614 193095 158616
rect 192956 158612 192962 158614
rect 193029 158611 193095 158614
rect 193990 158612 193996 158676
rect 194060 158674 194066 158676
rect 194133 158674 194199 158677
rect 194060 158672 194199 158674
rect 194060 158616 194138 158672
rect 194194 158616 194199 158672
rect 194060 158614 194199 158616
rect 194060 158612 194066 158614
rect 194133 158611 194199 158614
rect 195278 158612 195284 158676
rect 195348 158674 195354 158676
rect 195605 158674 195671 158677
rect 195881 158676 195947 158677
rect 195830 158674 195836 158676
rect 195348 158672 195671 158674
rect 195348 158616 195610 158672
rect 195666 158616 195671 158672
rect 195348 158614 195671 158616
rect 195790 158614 195836 158674
rect 195900 158672 195947 158676
rect 195942 158616 195947 158672
rect 195348 158612 195354 158614
rect 195605 158611 195671 158614
rect 195830 158612 195836 158614
rect 195900 158612 195947 158616
rect 195881 158611 195947 158612
rect 196065 158674 196131 158677
rect 196198 158674 196204 158676
rect 196065 158672 196204 158674
rect 196065 158616 196070 158672
rect 196126 158616 196204 158672
rect 196065 158614 196204 158616
rect 196065 158611 196131 158614
rect 196198 158612 196204 158614
rect 196268 158612 196274 158676
rect 196750 158612 196756 158676
rect 196820 158674 196826 158676
rect 197261 158674 197327 158677
rect 198273 158676 198339 158677
rect 198222 158674 198228 158676
rect 196820 158672 197327 158674
rect 196820 158616 197266 158672
rect 197322 158616 197327 158672
rect 196820 158614 197327 158616
rect 198182 158614 198228 158674
rect 198292 158672 198339 158676
rect 198334 158616 198339 158672
rect 196820 158612 196826 158614
rect 197261 158611 197327 158614
rect 198222 158612 198228 158614
rect 198292 158612 198339 158616
rect 198273 158611 198339 158612
rect 199193 158674 199259 158677
rect 199837 158676 199903 158677
rect 199326 158674 199332 158676
rect 199193 158672 199332 158674
rect 199193 158616 199198 158672
rect 199254 158616 199332 158672
rect 199193 158614 199332 158616
rect 199193 158611 199259 158614
rect 199326 158612 199332 158614
rect 199396 158612 199402 158676
rect 199837 158672 199884 158676
rect 199948 158674 199954 158676
rect 200205 158674 200271 158677
rect 200941 158676 201007 158677
rect 200614 158674 200620 158676
rect 199837 158616 199842 158672
rect 199837 158612 199884 158616
rect 199948 158614 199994 158674
rect 200205 158672 200620 158674
rect 200205 158616 200210 158672
rect 200266 158616 200620 158672
rect 200205 158614 200620 158616
rect 199948 158612 199954 158614
rect 199837 158611 199903 158612
rect 200205 158611 200271 158614
rect 200614 158612 200620 158614
rect 200684 158612 200690 158676
rect 200941 158672 200988 158676
rect 201052 158674 201058 158676
rect 202413 158674 202479 158677
rect 202638 158674 202644 158676
rect 200941 158616 200946 158672
rect 200941 158612 200988 158616
rect 201052 158614 201098 158674
rect 202413 158672 202644 158674
rect 202413 158616 202418 158672
rect 202474 158616 202644 158672
rect 202413 158614 202644 158616
rect 201052 158612 201058 158614
rect 200941 158611 201007 158612
rect 202413 158611 202479 158614
rect 202638 158612 202644 158614
rect 202708 158612 202714 158676
rect 202965 158674 203031 158677
rect 203977 158676 204043 158677
rect 203742 158674 203748 158676
rect 202965 158672 203748 158674
rect 202965 158616 202970 158672
rect 203026 158616 203748 158672
rect 202965 158614 203748 158616
rect 202965 158611 203031 158614
rect 203742 158612 203748 158614
rect 203812 158612 203818 158676
rect 203926 158674 203932 158676
rect 203886 158614 203932 158674
rect 203996 158672 204043 158676
rect 204038 158616 204043 158672
rect 203926 158612 203932 158614
rect 203996 158612 204043 158616
rect 203977 158611 204043 158612
rect 204345 158674 204411 158677
rect 205030 158674 205036 158676
rect 204345 158672 205036 158674
rect 204345 158616 204350 158672
rect 204406 158616 205036 158672
rect 204345 158614 205036 158616
rect 204345 158611 204411 158614
rect 205030 158612 205036 158614
rect 205100 158612 205106 158676
rect 207013 158674 207079 158677
rect 209078 158674 209084 158676
rect 207013 158672 209084 158674
rect 207013 158616 207018 158672
rect 207074 158616 209084 158672
rect 207013 158614 209084 158616
rect 207013 158611 207079 158614
rect 209078 158612 209084 158614
rect 209148 158612 209154 158676
rect 165724 158536 166783 158538
rect 165724 158480 166722 158536
rect 166778 158480 166783 158536
rect 165724 158478 166783 158480
rect 165724 158476 165730 158478
rect 166717 158475 166783 158478
rect 166950 158478 176670 158538
rect 177438 158478 209790 158538
rect 162894 158340 162900 158404
rect 162964 158402 162970 158404
rect 163957 158402 164023 158405
rect 162964 158400 164023 158402
rect 162964 158344 163962 158400
rect 164018 158344 164023 158400
rect 162964 158342 164023 158344
rect 162964 158340 162970 158342
rect 163957 158339 164023 158342
rect 164233 158402 164299 158405
rect 164877 158402 164943 158405
rect 166950 158402 167010 158478
rect 164233 158400 164943 158402
rect 164233 158344 164238 158400
rect 164294 158344 164882 158400
rect 164938 158344 164943 158400
rect 164233 158342 164943 158344
rect 164233 158339 164299 158342
rect 164877 158339 164943 158342
rect 166766 158342 167010 158402
rect 167453 158402 167519 158405
rect 168230 158402 168236 158404
rect 167453 158400 168236 158402
rect 167453 158344 167458 158400
rect 167514 158344 168236 158400
rect 167453 158342 168236 158344
rect 164325 158266 164391 158269
rect 166766 158266 166826 158342
rect 167453 158339 167519 158342
rect 168230 158340 168236 158342
rect 168300 158340 168306 158404
rect 168373 158402 168439 158405
rect 169477 158402 169543 158405
rect 170990 158402 170996 158404
rect 168373 158400 169543 158402
rect 168373 158344 168378 158400
rect 168434 158344 169482 158400
rect 169538 158344 169543 158400
rect 168373 158342 169543 158344
rect 168373 158339 168439 158342
rect 169477 158339 169543 158342
rect 169710 158342 170996 158402
rect 164325 158264 166826 158266
rect 164325 158208 164330 158264
rect 164386 158208 166826 158264
rect 164325 158206 166826 158208
rect 164325 158203 164391 158206
rect 166942 158204 166948 158268
rect 167012 158266 167018 158268
rect 168281 158266 168347 158269
rect 167012 158264 168347 158266
rect 167012 158208 168286 158264
rect 168342 158208 168347 158264
rect 167012 158206 168347 158208
rect 167012 158204 167018 158206
rect 168281 158203 168347 158206
rect 168465 158266 168531 158269
rect 168966 158266 168972 158268
rect 168465 158264 168972 158266
rect 168465 158208 168470 158264
rect 168526 158208 168972 158264
rect 168465 158206 168972 158208
rect 168465 158203 168531 158206
rect 168966 158204 168972 158206
rect 169036 158266 169042 158268
rect 169710 158266 169770 158342
rect 170990 158340 170996 158342
rect 171060 158340 171066 158404
rect 171174 158340 171180 158404
rect 171244 158402 171250 158404
rect 171593 158402 171659 158405
rect 171244 158400 171659 158402
rect 171244 158344 171598 158400
rect 171654 158344 171659 158400
rect 171244 158342 171659 158344
rect 171244 158340 171250 158342
rect 171593 158339 171659 158342
rect 173985 158402 174051 158405
rect 175038 158402 175044 158404
rect 173985 158400 175044 158402
rect 173985 158344 173990 158400
rect 174046 158344 175044 158400
rect 173985 158342 175044 158344
rect 173985 158339 174051 158342
rect 175038 158340 175044 158342
rect 175108 158340 175114 158404
rect 175273 158402 175339 158405
rect 175958 158402 175964 158404
rect 175273 158400 175964 158402
rect 175273 158344 175278 158400
rect 175334 158344 175964 158400
rect 175273 158342 175964 158344
rect 175273 158339 175339 158342
rect 175958 158340 175964 158342
rect 176028 158340 176034 158404
rect 176610 158402 176670 158478
rect 197905 158402 197971 158405
rect 176610 158400 197971 158402
rect 176610 158344 197910 158400
rect 197966 158344 197971 158400
rect 176610 158342 197971 158344
rect 197905 158339 197971 158342
rect 198038 158340 198044 158404
rect 198108 158402 198114 158404
rect 198365 158402 198431 158405
rect 198108 158400 198431 158402
rect 198108 158344 198370 158400
rect 198426 158344 198431 158400
rect 198108 158342 198431 158344
rect 198108 158340 198114 158342
rect 198365 158339 198431 158342
rect 199510 158340 199516 158404
rect 199580 158402 199586 158404
rect 199929 158402 199995 158405
rect 199580 158400 199995 158402
rect 199580 158344 199934 158400
rect 199990 158344 199995 158400
rect 199580 158342 199995 158344
rect 199580 158340 199586 158342
rect 199929 158339 199995 158342
rect 201033 158402 201099 158405
rect 201401 158404 201467 158405
rect 201166 158402 201172 158404
rect 201033 158400 201172 158402
rect 201033 158344 201038 158400
rect 201094 158344 201172 158400
rect 201033 158342 201172 158344
rect 201033 158339 201099 158342
rect 201166 158340 201172 158342
rect 201236 158340 201242 158404
rect 201350 158340 201356 158404
rect 201420 158402 201467 158404
rect 202137 158402 202203 158405
rect 202454 158402 202460 158404
rect 201420 158400 201512 158402
rect 201462 158344 201512 158400
rect 201420 158342 201512 158344
rect 202137 158400 202460 158402
rect 202137 158344 202142 158400
rect 202198 158344 202460 158400
rect 202137 158342 202460 158344
rect 201420 158340 201467 158342
rect 201401 158339 201467 158340
rect 202137 158339 202203 158342
rect 202454 158340 202460 158342
rect 202524 158340 202530 158404
rect 204253 158402 204319 158405
rect 204662 158402 204668 158404
rect 204253 158400 204668 158402
rect 204253 158344 204258 158400
rect 204314 158344 204668 158400
rect 204253 158342 204668 158344
rect 204253 158339 204319 158342
rect 204662 158340 204668 158342
rect 204732 158340 204738 158404
rect 205173 158402 205239 158405
rect 209405 158402 209471 158405
rect 205173 158400 209471 158402
rect 205173 158344 205178 158400
rect 205234 158344 209410 158400
rect 209466 158344 209471 158400
rect 205173 158342 209471 158344
rect 205173 158339 205239 158342
rect 209405 158339 209471 158342
rect 169036 158206 169770 158266
rect 169036 158204 169042 158206
rect 169886 158204 169892 158268
rect 169956 158266 169962 158268
rect 170489 158266 170555 158269
rect 169956 158264 170555 158266
rect 169956 158208 170494 158264
rect 170550 158208 170555 158264
rect 169956 158206 170555 158208
rect 169956 158204 169962 158206
rect 170489 158203 170555 158206
rect 170622 158204 170628 158268
rect 170692 158266 170698 158268
rect 170857 158266 170923 158269
rect 170692 158264 170923 158266
rect 170692 158208 170862 158264
rect 170918 158208 170923 158264
rect 170692 158206 170923 158208
rect 170692 158204 170698 158206
rect 170857 158203 170923 158206
rect 172697 158266 172763 158269
rect 173382 158266 173388 158268
rect 172697 158264 173388 158266
rect 172697 158208 172702 158264
rect 172758 158208 173388 158264
rect 172697 158206 173388 158208
rect 172697 158203 172763 158206
rect 173382 158204 173388 158206
rect 173452 158204 173458 158268
rect 173985 158266 174051 158269
rect 174486 158266 174492 158268
rect 173985 158264 174492 158266
rect 173985 158208 173990 158264
rect 174046 158208 174492 158264
rect 173985 158206 174492 158208
rect 173985 158203 174051 158206
rect 174486 158204 174492 158206
rect 174556 158204 174562 158268
rect 175273 158266 175339 158269
rect 175917 158266 175983 158269
rect 206686 158266 206692 158268
rect 175273 158264 175983 158266
rect 175273 158208 175278 158264
rect 175334 158208 175922 158264
rect 175978 158208 175983 158264
rect 175273 158206 175983 158208
rect 175273 158203 175339 158206
rect 175917 158203 175983 158206
rect 176610 158206 206692 158266
rect 158621 158130 158687 158133
rect 165838 158130 165844 158132
rect 158621 158128 165844 158130
rect 158621 158072 158626 158128
rect 158682 158072 165844 158128
rect 158621 158070 165844 158072
rect 158621 158067 158687 158070
rect 165838 158068 165844 158070
rect 165908 158068 165914 158132
rect 166257 158130 166323 158133
rect 168465 158130 168531 158133
rect 166257 158128 168531 158130
rect 166257 158072 166262 158128
rect 166318 158072 168470 158128
rect 168526 158072 168531 158128
rect 166257 158070 168531 158072
rect 166257 158067 166323 158070
rect 168465 158067 168531 158070
rect 168598 158068 168604 158132
rect 168668 158130 168674 158132
rect 168925 158130 168991 158133
rect 168668 158128 168991 158130
rect 168668 158072 168930 158128
rect 168986 158072 168991 158128
rect 168668 158070 168991 158072
rect 168668 158068 168674 158070
rect 168925 158067 168991 158070
rect 170254 158068 170260 158132
rect 170324 158130 170330 158132
rect 170673 158130 170739 158133
rect 170324 158128 170739 158130
rect 170324 158072 170678 158128
rect 170734 158072 170739 158128
rect 170324 158070 170739 158072
rect 170324 158068 170330 158070
rect 170673 158067 170739 158070
rect 170806 158068 170812 158132
rect 170876 158130 170882 158132
rect 170949 158130 171015 158133
rect 170876 158128 171015 158130
rect 170876 158072 170954 158128
rect 171010 158072 171015 158128
rect 170876 158070 171015 158072
rect 170876 158068 170882 158070
rect 170949 158067 171015 158070
rect 171961 158130 172027 158133
rect 176326 158130 176332 158132
rect 171961 158128 176332 158130
rect 171961 158072 171966 158128
rect 172022 158072 176332 158128
rect 171961 158070 176332 158072
rect 171961 158067 172027 158070
rect 176326 158068 176332 158070
rect 176396 158068 176402 158132
rect 159725 157994 159791 157997
rect 163497 157994 163563 157997
rect 159725 157992 163563 157994
rect 159725 157936 159730 157992
rect 159786 157936 163502 157992
rect 163558 157936 163563 157992
rect 159725 157934 163563 157936
rect 159725 157931 159791 157934
rect 163497 157931 163563 157934
rect 164601 157994 164667 157997
rect 176610 157994 176670 158206
rect 206686 158204 206692 158206
rect 206756 158204 206762 158268
rect 207657 158266 207723 158269
rect 206878 158264 207723 158266
rect 206878 158208 207662 158264
rect 207718 158208 207723 158264
rect 206878 158206 207723 158208
rect 177430 158068 177436 158132
rect 177500 158130 177506 158132
rect 177757 158130 177823 158133
rect 177500 158128 177823 158130
rect 177500 158072 177762 158128
rect 177818 158072 177823 158128
rect 177500 158070 177823 158072
rect 177500 158068 177506 158070
rect 177757 158067 177823 158070
rect 181478 158068 181484 158132
rect 181548 158130 181554 158132
rect 181989 158130 182055 158133
rect 181548 158128 182055 158130
rect 181548 158072 181994 158128
rect 182050 158072 182055 158128
rect 181548 158070 182055 158072
rect 181548 158068 181554 158070
rect 181989 158067 182055 158070
rect 182817 158130 182883 158133
rect 183461 158130 183527 158133
rect 182817 158128 183527 158130
rect 182817 158072 182822 158128
rect 182878 158072 183466 158128
rect 183522 158072 183527 158128
rect 182817 158070 183527 158072
rect 182817 158067 182883 158070
rect 183461 158067 183527 158070
rect 186957 158130 187023 158133
rect 187182 158130 187188 158132
rect 186957 158128 187188 158130
rect 186957 158072 186962 158128
rect 187018 158072 187188 158128
rect 186957 158070 187188 158072
rect 186957 158067 187023 158070
rect 187182 158068 187188 158070
rect 187252 158068 187258 158132
rect 190453 158130 190519 158133
rect 191649 158130 191715 158133
rect 190453 158128 191715 158130
rect 190453 158072 190458 158128
rect 190514 158072 191654 158128
rect 191710 158072 191715 158128
rect 190453 158070 191715 158072
rect 190453 158067 190519 158070
rect 191649 158067 191715 158070
rect 193305 158130 193371 158133
rect 194358 158130 194364 158132
rect 193305 158128 194364 158130
rect 193305 158072 193310 158128
rect 193366 158072 194364 158128
rect 193305 158070 194364 158072
rect 193305 158067 193371 158070
rect 194358 158068 194364 158070
rect 194428 158068 194434 158132
rect 194685 158130 194751 158133
rect 195462 158130 195468 158132
rect 194685 158128 195468 158130
rect 194685 158072 194690 158128
rect 194746 158072 195468 158128
rect 194685 158070 195468 158072
rect 194685 158067 194751 158070
rect 195462 158068 195468 158070
rect 195532 158068 195538 158132
rect 196065 158130 196131 158133
rect 196382 158130 196388 158132
rect 196065 158128 196388 158130
rect 196065 158072 196070 158128
rect 196126 158072 196388 158128
rect 196065 158070 196388 158072
rect 196065 158067 196131 158070
rect 196382 158068 196388 158070
rect 196452 158068 196458 158132
rect 197905 158130 197971 158133
rect 206878 158130 206938 158206
rect 207657 158203 207723 158206
rect 197905 158128 206938 158130
rect 197905 158072 197910 158128
rect 197966 158072 206938 158128
rect 197905 158070 206938 158072
rect 207105 158130 207171 158133
rect 207974 158130 207980 158132
rect 207105 158128 207980 158130
rect 207105 158072 207110 158128
rect 207166 158072 207980 158128
rect 207105 158070 207980 158072
rect 197905 158067 197971 158070
rect 207105 158067 207171 158070
rect 207974 158068 207980 158070
rect 208044 158130 208050 158132
rect 208209 158130 208275 158133
rect 208044 158128 208275 158130
rect 208044 158072 208214 158128
rect 208270 158072 208275 158128
rect 208044 158070 208275 158072
rect 209730 158130 209790 158478
rect 210509 158130 210575 158133
rect 209730 158128 210575 158130
rect 209730 158072 210514 158128
rect 210570 158072 210575 158128
rect 209730 158070 210575 158072
rect 208044 158068 208050 158070
rect 208209 158067 208275 158070
rect 210509 158067 210575 158070
rect 164601 157992 176670 157994
rect 164601 157936 164606 157992
rect 164662 157936 176670 157992
rect 164601 157934 176670 157936
rect 164601 157931 164667 157934
rect 177246 157932 177252 157996
rect 177316 157994 177322 157996
rect 177849 157994 177915 157997
rect 177316 157992 177915 157994
rect 177316 157936 177854 157992
rect 177910 157936 177915 157992
rect 177316 157934 177915 157936
rect 177316 157932 177322 157934
rect 177849 157931 177915 157934
rect 199101 157994 199167 157997
rect 200021 157994 200087 157997
rect 199101 157992 200087 157994
rect 199101 157936 199106 157992
rect 199162 157936 200026 157992
rect 200082 157936 200087 157992
rect 199101 157934 200087 157936
rect 199101 157931 199167 157934
rect 200021 157931 200087 157934
rect 200297 157994 200363 157997
rect 201350 157994 201356 157996
rect 200297 157992 201356 157994
rect 200297 157936 200302 157992
rect 200358 157936 201356 157992
rect 200297 157934 201356 157936
rect 200297 157931 200363 157934
rect 201350 157932 201356 157934
rect 201420 157932 201426 157996
rect 202086 157932 202092 157996
rect 202156 157994 202162 157996
rect 202689 157994 202755 157997
rect 202156 157992 202755 157994
rect 202156 157936 202694 157992
rect 202750 157936 202755 157992
rect 202156 157934 202755 157936
rect 202156 157932 202162 157934
rect 202689 157931 202755 157934
rect 208485 157994 208551 157997
rect 244774 157994 244780 157996
rect 208485 157992 244780 157994
rect 208485 157936 208490 157992
rect 208546 157936 244780 157992
rect 208485 157934 244780 157936
rect 208485 157931 208551 157934
rect 244774 157932 244780 157934
rect 244844 157932 244850 157996
rect 157333 157858 157399 157861
rect 157793 157858 157859 157861
rect 163681 157858 163747 157861
rect 164325 157860 164391 157861
rect 164325 157858 164372 157860
rect 157333 157856 163747 157858
rect 157333 157800 157338 157856
rect 157394 157800 157798 157856
rect 157854 157800 163686 157856
rect 163742 157800 163747 157856
rect 157333 157798 163747 157800
rect 164280 157856 164372 157858
rect 164280 157800 164330 157856
rect 164280 157798 164372 157800
rect 157333 157795 157399 157798
rect 157793 157795 157859 157798
rect 163681 157795 163747 157798
rect 164325 157796 164372 157798
rect 164436 157796 164442 157860
rect 165245 157858 165311 157861
rect 176377 157858 176443 157861
rect 165245 157856 176443 157858
rect 165245 157800 165250 157856
rect 165306 157800 176382 157856
rect 176438 157800 176443 157856
rect 165245 157798 176443 157800
rect 164325 157795 164391 157796
rect 165245 157795 165311 157798
rect 176377 157795 176443 157798
rect 177205 157858 177271 157861
rect 177982 157858 177988 157860
rect 177205 157856 177988 157858
rect 177205 157800 177210 157856
rect 177266 157800 177988 157856
rect 177205 157798 177988 157800
rect 177205 157795 177271 157798
rect 177982 157796 177988 157798
rect 178052 157796 178058 157860
rect 186446 157796 186452 157860
rect 186516 157858 186522 157860
rect 198825 157858 198891 157861
rect 199929 157858 199995 157861
rect 186516 157798 195990 157858
rect 186516 157796 186522 157798
rect 160001 157722 160067 157725
rect 166758 157722 166764 157724
rect 160001 157720 166764 157722
rect 160001 157664 160006 157720
rect 160062 157664 166764 157720
rect 160001 157662 166764 157664
rect 160001 157659 160067 157662
rect 166758 157660 166764 157662
rect 166828 157660 166834 157724
rect 166993 157722 167059 157725
rect 168230 157722 168236 157724
rect 166993 157720 168236 157722
rect 166993 157664 166998 157720
rect 167054 157664 168236 157720
rect 166993 157662 168236 157664
rect 166993 157659 167059 157662
rect 168230 157660 168236 157662
rect 168300 157660 168306 157724
rect 168465 157722 168531 157725
rect 174445 157722 174511 157725
rect 168465 157720 174511 157722
rect 168465 157664 168470 157720
rect 168526 157664 174450 157720
rect 174506 157664 174511 157720
rect 168465 157662 174511 157664
rect 195930 157722 195990 157798
rect 198825 157856 199995 157858
rect 198825 157800 198830 157856
rect 198886 157800 199934 157856
rect 199990 157800 199995 157856
rect 198825 157798 199995 157800
rect 198825 157795 198891 157798
rect 199929 157795 199995 157798
rect 207381 157858 207447 157861
rect 208301 157858 208367 157861
rect 207381 157856 208367 157858
rect 207381 157800 207386 157856
rect 207442 157800 208306 157856
rect 208362 157800 208367 157856
rect 207381 157798 208367 157800
rect 207381 157795 207447 157798
rect 208301 157795 208367 157798
rect 202822 157722 202828 157724
rect 195930 157662 202828 157722
rect 168465 157659 168531 157662
rect 174445 157659 174511 157662
rect 202822 157660 202828 157662
rect 202892 157660 202898 157724
rect 207289 157722 207355 157725
rect 208117 157722 208183 157725
rect 209262 157722 209268 157724
rect 207289 157720 209268 157722
rect 207289 157664 207294 157720
rect 207350 157664 208122 157720
rect 208178 157664 209268 157720
rect 207289 157662 209268 157664
rect 207289 157659 207355 157662
rect 208117 157659 208183 157662
rect 209262 157660 209268 157662
rect 209332 157660 209338 157724
rect 158161 157586 158227 157589
rect 166257 157586 166323 157589
rect 158161 157584 166323 157586
rect 158161 157528 158166 157584
rect 158222 157528 166262 157584
rect 166318 157528 166323 157584
rect 158161 157526 166323 157528
rect 158161 157523 158227 157526
rect 166257 157523 166323 157526
rect 169702 157524 169708 157588
rect 169772 157586 169778 157588
rect 170765 157586 170831 157589
rect 192385 157588 192451 157589
rect 192334 157586 192340 157588
rect 169772 157584 170831 157586
rect 169772 157528 170770 157584
rect 170826 157528 170831 157584
rect 169772 157526 170831 157528
rect 192294 157526 192340 157586
rect 192404 157584 192451 157588
rect 210325 157586 210391 157589
rect 192446 157528 192451 157584
rect 169772 157524 169778 157526
rect 170765 157523 170831 157526
rect 192334 157524 192340 157526
rect 192404 157524 192451 157528
rect 192385 157523 192451 157524
rect 195930 157584 210391 157586
rect 195930 157528 210330 157584
rect 210386 157528 210391 157584
rect 195930 157526 210391 157528
rect 157425 157450 157491 157453
rect 158345 157450 158411 157453
rect 163497 157450 163563 157453
rect 157425 157448 163563 157450
rect 157425 157392 157430 157448
rect 157486 157392 158350 157448
rect 158406 157392 163502 157448
rect 163558 157392 163563 157448
rect 157425 157390 163563 157392
rect 157425 157387 157491 157390
rect 158345 157387 158411 157390
rect 163497 157387 163563 157390
rect 164141 157450 164207 157453
rect 195930 157450 195990 157526
rect 210325 157523 210391 157526
rect 164141 157448 195990 157450
rect 164141 157392 164146 157448
rect 164202 157392 195990 157448
rect 164141 157390 195990 157392
rect 164141 157387 164207 157390
rect 200798 157388 200804 157452
rect 200868 157450 200874 157452
rect 201309 157450 201375 157453
rect 200868 157448 201375 157450
rect 200868 157392 201314 157448
rect 201370 157392 201375 157448
rect 200868 157390 201375 157392
rect 200868 157388 200874 157390
rect 201309 157387 201375 157390
rect 157241 157314 157307 157317
rect 158069 157314 158135 157317
rect 164366 157314 164372 157316
rect 157241 157312 157350 157314
rect 157241 157256 157246 157312
rect 157302 157256 157350 157312
rect 157241 157251 157350 157256
rect 158069 157312 164372 157314
rect 158069 157256 158074 157312
rect 158130 157256 164372 157312
rect 158069 157254 164372 157256
rect 158069 157251 158135 157254
rect 164366 157252 164372 157254
rect 164436 157314 164442 157316
rect 164785 157314 164851 157317
rect 164436 157312 164851 157314
rect 164436 157256 164790 157312
rect 164846 157256 164851 157312
rect 164436 157254 164851 157256
rect 164436 157252 164442 157254
rect 164785 157251 164851 157254
rect 170121 157314 170187 157317
rect 170438 157314 170444 157316
rect 170121 157312 170444 157314
rect 170121 157256 170126 157312
rect 170182 157256 170444 157312
rect 170121 157254 170444 157256
rect 170121 157251 170187 157254
rect 170438 157252 170444 157254
rect 170508 157252 170514 157316
rect 173341 157314 173407 157317
rect 173750 157314 173756 157316
rect 173341 157312 173756 157314
rect 173341 157256 173346 157312
rect 173402 157256 173756 157312
rect 173341 157254 173756 157256
rect 173341 157251 173407 157254
rect 173750 157252 173756 157254
rect 173820 157252 173826 157316
rect 188286 157252 188292 157316
rect 188356 157314 188362 157316
rect 188981 157314 189047 157317
rect 192385 157316 192451 157317
rect 192334 157314 192340 157316
rect 188356 157312 191114 157314
rect 188356 157256 188986 157312
rect 189042 157256 191114 157312
rect 188356 157254 191114 157256
rect 192294 157254 192340 157314
rect 192404 157312 192451 157316
rect 192446 157256 192451 157312
rect 188356 157252 188362 157254
rect 188981 157251 189047 157254
rect 157290 157178 157350 157251
rect 162894 157178 162900 157180
rect 157290 157118 162900 157178
rect 162894 157116 162900 157118
rect 162964 157178 162970 157180
rect 164049 157178 164115 157181
rect 162964 157176 164115 157178
rect 162964 157120 164054 157176
rect 164110 157120 164115 157176
rect 162964 157118 164115 157120
rect 162964 157116 162970 157118
rect 164049 157115 164115 157118
rect 155585 157042 155651 157045
rect 165981 157042 166047 157045
rect 155585 157040 166047 157042
rect 155585 156984 155590 157040
rect 155646 156984 165986 157040
rect 166042 156984 166047 157040
rect 155585 156982 166047 156984
rect 191054 157042 191114 157254
rect 192334 157252 192340 157254
rect 192404 157252 192451 157256
rect 192385 157251 192451 157252
rect 200665 157314 200731 157317
rect 270585 157314 270651 157317
rect 200665 157312 270651 157314
rect 200665 157256 200670 157312
rect 200726 157256 270590 157312
rect 270646 157256 270651 157312
rect 200665 157254 270651 157256
rect 200665 157251 200731 157254
rect 270585 157251 270651 157254
rect 199878 157116 199884 157180
rect 199948 157178 199954 157180
rect 239673 157178 239739 157181
rect 199948 157176 239739 157178
rect 199948 157120 239678 157176
rect 239734 157120 239739 157176
rect 199948 157118 239739 157120
rect 199948 157116 199954 157118
rect 239673 157115 239739 157118
rect 217685 157042 217751 157045
rect 191054 157040 217751 157042
rect 191054 156984 217690 157040
rect 217746 156984 217751 157040
rect 191054 156982 217751 156984
rect 155585 156979 155651 156982
rect 165981 156979 166047 156982
rect 217685 156979 217751 156982
rect 159817 156906 159883 156909
rect 168414 156906 168420 156908
rect 159817 156904 168420 156906
rect 159817 156848 159822 156904
rect 159878 156848 168420 156904
rect 159817 156846 168420 156848
rect 159817 156843 159883 156846
rect 168414 156844 168420 156846
rect 168484 156844 168490 156908
rect 200849 156906 200915 156909
rect 201033 156906 201099 156909
rect 200849 156904 201099 156906
rect 200849 156848 200854 156904
rect 200910 156848 201038 156904
rect 201094 156848 201099 156904
rect 200849 156846 201099 156848
rect 200849 156843 200915 156846
rect 201033 156843 201099 156846
rect 152825 156770 152891 156773
rect 168833 156770 168899 156773
rect 152825 156768 168899 156770
rect 152825 156712 152830 156768
rect 152886 156712 168838 156768
rect 168894 156712 168899 156768
rect 152825 156710 168899 156712
rect 152825 156707 152891 156710
rect 168833 156707 168899 156710
rect 194501 156770 194567 156773
rect 213085 156770 213151 156773
rect 194501 156768 213151 156770
rect 194501 156712 194506 156768
rect 194562 156712 213090 156768
rect 213146 156712 213151 156768
rect 194501 156710 213151 156712
rect 194501 156707 194567 156710
rect 213085 156707 213151 156710
rect 156505 156634 156571 156637
rect 156873 156634 156939 156637
rect 168005 156634 168071 156637
rect 156505 156632 168071 156634
rect 156505 156576 156510 156632
rect 156566 156576 156878 156632
rect 156934 156576 168010 156632
rect 168066 156576 168071 156632
rect 156505 156574 168071 156576
rect 156505 156571 156571 156574
rect 156873 156571 156939 156574
rect 168005 156571 168071 156574
rect 179045 156634 179111 156637
rect 213913 156634 213979 156637
rect 179045 156632 213979 156634
rect 179045 156576 179050 156632
rect 179106 156576 213918 156632
rect 213974 156576 213979 156632
rect 179045 156574 213979 156576
rect 179045 156571 179111 156574
rect 213913 156571 213979 156574
rect 163262 156436 163268 156500
rect 163332 156498 163338 156500
rect 163497 156498 163563 156501
rect 163332 156496 163563 156498
rect 163332 156440 163502 156496
rect 163558 156440 163563 156496
rect 163332 156438 163563 156440
rect 163332 156436 163338 156438
rect 163497 156435 163563 156438
rect 198457 156498 198523 156501
rect 210785 156498 210851 156501
rect 198457 156496 210851 156498
rect 198457 156440 198462 156496
rect 198518 156440 210790 156496
rect 210846 156440 210851 156496
rect 198457 156438 210851 156440
rect 198457 156435 198523 156438
rect 210785 156435 210851 156438
rect 192477 156090 192543 156093
rect 193121 156090 193187 156093
rect 192477 156088 193187 156090
rect 192477 156032 192482 156088
rect 192538 156032 193126 156088
rect 193182 156032 193187 156088
rect 192477 156030 193187 156032
rect 192477 156027 192543 156030
rect 193121 156027 193187 156030
rect 201861 156090 201927 156093
rect 202270 156090 202276 156092
rect 201861 156088 202276 156090
rect 201861 156032 201866 156088
rect 201922 156032 202276 156088
rect 201861 156030 202276 156032
rect 201861 156027 201927 156030
rect 202270 156028 202276 156030
rect 202340 156028 202346 156092
rect 196801 155954 196867 155957
rect 208393 155954 208459 155957
rect 196801 155952 208459 155954
rect 196801 155896 196806 155952
rect 196862 155896 208398 155952
rect 208454 155896 208459 155952
rect 196801 155894 208459 155896
rect 196801 155891 196867 155894
rect 208393 155891 208459 155894
rect 190821 155818 190887 155821
rect 207473 155818 207539 155821
rect 190821 155816 207539 155818
rect 190821 155760 190826 155816
rect 190882 155760 207478 155816
rect 207534 155760 207539 155816
rect 190821 155758 207539 155760
rect 190821 155755 190887 155758
rect 207473 155755 207539 155758
rect 210417 155682 210483 155685
rect 267917 155682 267983 155685
rect 210417 155680 267983 155682
rect 210417 155624 210422 155680
rect 210478 155624 267922 155680
rect 267978 155624 267983 155680
rect 210417 155622 267983 155624
rect 210417 155619 210483 155622
rect 267917 155619 267983 155622
rect 202873 155546 202939 155549
rect 204161 155546 204227 155549
rect 267825 155546 267891 155549
rect 202873 155544 267891 155546
rect 202873 155488 202878 155544
rect 202934 155488 204166 155544
rect 204222 155488 267830 155544
rect 267886 155488 267891 155544
rect 202873 155486 267891 155488
rect 202873 155483 202939 155486
rect 204161 155483 204227 155486
rect 267825 155483 267891 155486
rect 195278 155348 195284 155412
rect 195348 155410 195354 155412
rect 197905 155410 197971 155413
rect 195348 155408 197971 155410
rect 195348 155352 197910 155408
rect 197966 155352 197971 155408
rect 195348 155350 197971 155352
rect 195348 155348 195354 155350
rect 197905 155347 197971 155350
rect 100753 155274 100819 155277
rect 157333 155274 157399 155277
rect 100753 155272 157399 155274
rect 100753 155216 100758 155272
rect 100814 155216 157338 155272
rect 157394 155216 157399 155272
rect 100753 155214 157399 155216
rect 100753 155211 100819 155214
rect 157333 155211 157399 155214
rect 193397 155274 193463 155277
rect 204529 155274 204595 155277
rect 205449 155274 205515 155277
rect 270677 155274 270743 155277
rect 384297 155274 384363 155277
rect 193397 155272 195990 155274
rect 193397 155216 193402 155272
rect 193458 155216 195990 155272
rect 193397 155214 195990 155216
rect 193397 155211 193463 155214
rect 195930 155138 195990 155214
rect 204529 155272 270743 155274
rect 204529 155216 204534 155272
rect 204590 155216 205454 155272
rect 205510 155216 270682 155272
rect 270738 155216 270743 155272
rect 204529 155214 270743 155216
rect 204529 155211 204595 155214
rect 205449 155211 205515 155214
rect 270677 155211 270743 155214
rect 277350 155272 384363 155274
rect 277350 155216 384302 155272
rect 384358 155216 384363 155272
rect 277350 155214 384363 155216
rect 277025 155138 277091 155141
rect 277350 155138 277410 155214
rect 384297 155211 384363 155214
rect 195930 155136 277410 155138
rect 195930 155080 277030 155136
rect 277086 155080 277410 155136
rect 195930 155078 277410 155080
rect 277025 155075 277091 155078
rect 197905 155002 197971 155005
rect 211705 155002 211771 155005
rect 197905 155000 211771 155002
rect 197905 154944 197910 155000
rect 197966 154944 211710 155000
rect 211766 154944 211771 155000
rect 197905 154942 211771 154944
rect 197905 154939 197971 154942
rect 211705 154939 211771 154942
rect 201677 154866 201743 154869
rect 202689 154866 202755 154869
rect 210417 154866 210483 154869
rect 201677 154864 210483 154866
rect 201677 154808 201682 154864
rect 201738 154808 202694 154864
rect 202750 154808 210422 154864
rect 210478 154808 210483 154864
rect 201677 154806 210483 154808
rect 201677 154803 201743 154806
rect 202689 154803 202755 154806
rect 210417 154803 210483 154806
rect 199653 154730 199719 154733
rect 203609 154730 203675 154733
rect 199653 154728 203675 154730
rect 199653 154672 199658 154728
rect 199714 154672 203614 154728
rect 203670 154672 203675 154728
rect 199653 154670 203675 154672
rect 199653 154667 199719 154670
rect 203609 154667 203675 154670
rect 199694 154532 199700 154596
rect 199764 154594 199770 154596
rect 199837 154594 199903 154597
rect 199764 154592 199903 154594
rect 199764 154536 199842 154592
rect 199898 154536 199903 154592
rect 199764 154534 199903 154536
rect 199764 154532 199770 154534
rect 199837 154531 199903 154534
rect 203149 154458 203215 154461
rect 262949 154458 263015 154461
rect 203149 154456 263015 154458
rect 203149 154400 203154 154456
rect 203210 154400 262954 154456
rect 263010 154400 263015 154456
rect 203149 154398 263015 154400
rect 203149 154395 203215 154398
rect 262949 154395 263015 154398
rect 205357 154322 205423 154325
rect 238477 154322 238543 154325
rect 205357 154320 238543 154322
rect 205357 154264 205362 154320
rect 205418 154264 238482 154320
rect 238538 154264 238543 154320
rect 205357 154262 238543 154264
rect 205357 154259 205423 154262
rect 238477 154259 238543 154262
rect 200982 154124 200988 154188
rect 201052 154186 201058 154188
rect 240869 154186 240935 154189
rect 201052 154184 240935 154186
rect 201052 154128 240874 154184
rect 240930 154128 240935 154184
rect 201052 154126 240935 154128
rect 201052 154124 201058 154126
rect 240869 154123 240935 154126
rect 126973 154050 127039 154053
rect 157425 154050 157491 154053
rect 126973 154048 157491 154050
rect 126973 153992 126978 154048
rect 127034 153992 157430 154048
rect 157486 153992 157491 154048
rect 126973 153990 157491 153992
rect 126973 153987 127039 153990
rect 157425 153987 157491 153990
rect 177982 153988 177988 154052
rect 178052 154050 178058 154052
rect 212165 154050 212231 154053
rect 178052 154048 212231 154050
rect 178052 153992 212170 154048
rect 212226 153992 212231 154048
rect 178052 153990 212231 153992
rect 178052 153988 178058 153990
rect 212165 153987 212231 153990
rect 71037 153914 71103 153917
rect 155493 153914 155559 153917
rect 71037 153912 155559 153914
rect 71037 153856 71042 153912
rect 71098 153856 155498 153912
rect 155554 153856 155559 153912
rect 71037 153854 155559 153856
rect 71037 153851 71103 153854
rect 155493 153851 155559 153854
rect 203926 153852 203932 153916
rect 203996 153914 204002 153916
rect 236821 153914 236887 153917
rect 203996 153912 236887 153914
rect 203996 153856 236826 153912
rect 236882 153856 236887 153912
rect 203996 153854 236887 153856
rect 203996 153852 204002 153854
rect 236821 153851 236887 153854
rect 28993 153778 29059 153781
rect 155309 153778 155375 153781
rect 28993 153776 155375 153778
rect 28993 153720 28998 153776
rect 29054 153720 155314 153776
rect 155370 153720 155375 153776
rect 28993 153718 155375 153720
rect 28993 153715 29059 153718
rect 155309 153715 155375 153718
rect 157333 153778 157399 153781
rect 174670 153778 174676 153780
rect 157333 153776 174676 153778
rect 157333 153720 157338 153776
rect 157394 153720 174676 153776
rect 157333 153718 174676 153720
rect 157333 153715 157399 153718
rect 174670 153716 174676 153718
rect 174740 153778 174746 153780
rect 215017 153778 215083 153781
rect 174740 153776 215083 153778
rect 174740 153720 215022 153776
rect 215078 153720 215083 153776
rect 174740 153718 215083 153720
rect 174740 153716 174746 153718
rect 215017 153715 215083 153718
rect 197077 153642 197143 153645
rect 208485 153642 208551 153645
rect 197077 153640 208551 153642
rect 197077 153584 197082 153640
rect 197138 153584 208490 153640
rect 208546 153584 208551 153640
rect 197077 153582 208551 153584
rect 197077 153579 197143 153582
rect 208485 153579 208551 153582
rect 154573 153098 154639 153101
rect 158161 153098 158227 153101
rect 154573 153096 158227 153098
rect 154573 153040 154578 153096
rect 154634 153040 158166 153096
rect 158222 153040 158227 153096
rect 154573 153038 158227 153040
rect 154573 153035 154639 153038
rect 158161 153035 158227 153038
rect 171726 153036 171732 153100
rect 171796 153098 171802 153100
rect 172237 153098 172303 153101
rect 176193 153100 176259 153101
rect 171796 153096 174922 153098
rect 171796 153040 172242 153096
rect 172298 153040 174922 153096
rect 171796 153038 174922 153040
rect 171796 153036 171802 153038
rect 172237 153035 172303 153038
rect 174862 152826 174922 153038
rect 176142 153036 176148 153100
rect 176212 153098 176259 153100
rect 235533 153098 235599 153101
rect 176212 153096 176304 153098
rect 176254 153040 176304 153096
rect 176212 153038 176304 153040
rect 176610 153096 235599 153098
rect 176610 153040 235538 153096
rect 235594 153040 235599 153096
rect 176610 153038 235599 153040
rect 176212 153036 176259 153038
rect 176193 153035 176259 153036
rect 175958 152900 175964 152964
rect 176028 152962 176034 152964
rect 176610 152962 176670 153038
rect 235533 153035 235599 153038
rect 176028 152902 176670 152962
rect 176028 152900 176034 152902
rect 199326 152900 199332 152964
rect 199396 152962 199402 152964
rect 258574 152962 258580 152964
rect 199396 152902 258580 152962
rect 199396 152900 199402 152902
rect 258574 152900 258580 152902
rect 258644 152900 258650 152964
rect 217593 152826 217659 152829
rect 174862 152824 217659 152826
rect 174862 152768 217598 152824
rect 217654 152768 217659 152824
rect 174862 152766 217659 152768
rect 217593 152763 217659 152766
rect 192017 152690 192083 152693
rect 236494 152690 236500 152692
rect 192017 152688 236500 152690
rect 192017 152632 192022 152688
rect 192078 152632 236500 152688
rect 192017 152630 236500 152632
rect 192017 152627 192083 152630
rect 236494 152628 236500 152630
rect 236564 152628 236570 152692
rect 579889 152690 579955 152693
rect 583520 152690 584960 152780
rect 579889 152688 584960 152690
rect 579889 152632 579894 152688
rect 579950 152632 584960 152688
rect 579889 152630 584960 152632
rect 579889 152627 579955 152630
rect 199326 152492 199332 152556
rect 199396 152554 199402 152556
rect 199694 152554 199700 152556
rect 199396 152494 199700 152554
rect 199396 152492 199402 152494
rect 199694 152492 199700 152494
rect 199764 152492 199770 152556
rect 200297 152554 200363 152557
rect 220169 152554 220235 152557
rect 200297 152552 220235 152554
rect 200297 152496 200302 152552
rect 200358 152496 220174 152552
rect 220230 152496 220235 152552
rect 583520 152540 584960 152630
rect 200297 152494 220235 152496
rect 200297 152491 200363 152494
rect 220169 152491 220235 152494
rect 89713 152418 89779 152421
rect 152549 152418 152615 152421
rect 89713 152416 152615 152418
rect 89713 152360 89718 152416
rect 89774 152360 152554 152416
rect 152610 152360 152615 152416
rect 89713 152358 152615 152360
rect 89713 152355 89779 152358
rect 152549 152355 152615 152358
rect 198038 152356 198044 152420
rect 198108 152418 198114 152420
rect 213453 152418 213519 152421
rect 198108 152416 213519 152418
rect 198108 152360 213458 152416
rect 213514 152360 213519 152416
rect 198108 152358 213519 152360
rect 198108 152356 198114 152358
rect 213453 152355 213519 152358
rect 196750 152220 196756 152284
rect 196820 152282 196826 152284
rect 200297 152282 200363 152285
rect 196820 152280 200363 152282
rect 196820 152224 200302 152280
rect 200358 152224 200363 152280
rect 196820 152222 200363 152224
rect 196820 152220 196826 152222
rect 200297 152219 200363 152222
rect 193305 152146 193371 152149
rect 193581 152146 193647 152149
rect 193305 152144 193647 152146
rect 193305 152088 193310 152144
rect 193366 152088 193586 152144
rect 193642 152088 193647 152144
rect 193305 152086 193647 152088
rect 193305 152083 193371 152086
rect 193581 152083 193647 152086
rect 203793 151738 203859 151741
rect 273161 151738 273227 151741
rect 203793 151736 273227 151738
rect 203793 151680 203798 151736
rect 203854 151680 273166 151736
rect 273222 151680 273227 151736
rect 203793 151678 273227 151680
rect 203793 151675 203859 151678
rect 273161 151675 273227 151678
rect 201125 151602 201191 151605
rect 269757 151602 269823 151605
rect 201125 151600 269823 151602
rect 201125 151544 201130 151600
rect 201186 151544 269762 151600
rect 269818 151544 269823 151600
rect 201125 151542 269823 151544
rect 201125 151539 201191 151542
rect 269757 151539 269823 151542
rect 196617 151466 196683 151469
rect 254761 151466 254827 151469
rect 196617 151464 254827 151466
rect 196617 151408 196622 151464
rect 196678 151408 254766 151464
rect 254822 151408 254827 151464
rect 196617 151406 254827 151408
rect 196617 151403 196683 151406
rect 254761 151403 254827 151406
rect 64873 151330 64939 151333
rect 159357 151330 159423 151333
rect 64873 151328 159423 151330
rect 64873 151272 64878 151328
rect 64934 151272 159362 151328
rect 159418 151272 159423 151328
rect 64873 151270 159423 151272
rect 64873 151267 64939 151270
rect 159357 151267 159423 151270
rect 205173 151330 205239 151333
rect 253289 151330 253355 151333
rect 205173 151328 253355 151330
rect 205173 151272 205178 151328
rect 205234 151272 253294 151328
rect 253350 151272 253355 151328
rect 205173 151270 253355 151272
rect 205173 151267 205239 151270
rect 253289 151267 253355 151270
rect 51073 151194 51139 151197
rect 156965 151194 157031 151197
rect 51073 151192 157031 151194
rect 51073 151136 51078 151192
rect 51134 151136 156970 151192
rect 157026 151136 157031 151192
rect 51073 151134 157031 151136
rect 51073 151131 51139 151134
rect 156965 151131 157031 151134
rect 199561 151194 199627 151197
rect 226926 151194 226932 151196
rect 199561 151192 226932 151194
rect 199561 151136 199566 151192
rect 199622 151136 226932 151192
rect 199561 151134 226932 151136
rect 199561 151131 199627 151134
rect 226926 151132 226932 151134
rect 226996 151132 227002 151196
rect 269757 151194 269823 151197
rect 498285 151194 498351 151197
rect 269757 151192 498351 151194
rect 269757 151136 269762 151192
rect 269818 151136 498290 151192
rect 498346 151136 498351 151192
rect 269757 151134 498351 151136
rect 269757 151131 269823 151134
rect 498285 151131 498351 151134
rect 34513 151058 34579 151061
rect 149697 151058 149763 151061
rect 34513 151056 149763 151058
rect 34513 151000 34518 151056
rect 34574 151000 149702 151056
rect 149758 151000 149763 151056
rect 34513 150998 149763 151000
rect 34513 150995 34579 150998
rect 149697 150995 149763 150998
rect 178902 150996 178908 151060
rect 178972 151058 178978 151060
rect 212533 151058 212599 151061
rect 178972 151056 212599 151058
rect 178972 151000 212538 151056
rect 212594 151000 212599 151056
rect 178972 150998 212599 151000
rect 178972 150996 178978 150998
rect 212533 150995 212599 150998
rect 273161 151058 273227 151061
rect 536833 151058 536899 151061
rect 273161 151056 536899 151058
rect 273161 151000 273166 151056
rect 273222 151000 536838 151056
rect 536894 151000 536899 151056
rect 273161 150998 536899 151000
rect 273161 150995 273227 150998
rect 536833 150995 536899 150998
rect 204069 150378 204135 150381
rect 298185 150378 298251 150381
rect 299381 150378 299447 150381
rect 204069 150376 299447 150378
rect 204069 150320 204074 150376
rect 204130 150320 298190 150376
rect 298246 150320 299386 150376
rect 299442 150320 299447 150376
rect 204069 150318 299447 150320
rect 204069 150315 204135 150318
rect 298185 150315 298251 150318
rect 299381 150315 299447 150318
rect 201033 150242 201099 150245
rect 275645 150242 275711 150245
rect 201033 150240 275711 150242
rect 201033 150184 201038 150240
rect 201094 150184 275650 150240
rect 275706 150184 275711 150240
rect 201033 150182 275711 150184
rect 201033 150179 201099 150182
rect 275645 150179 275711 150182
rect 197905 150106 197971 150109
rect 257521 150106 257587 150109
rect 197905 150104 257587 150106
rect 197905 150048 197910 150104
rect 197966 150048 257526 150104
rect 257582 150048 257587 150104
rect 197905 150046 257587 150048
rect 197905 150043 197971 150046
rect 257521 150043 257587 150046
rect 135345 149970 135411 149973
rect 172830 149970 172836 149972
rect 135345 149968 172836 149970
rect -960 149834 480 149924
rect 135345 149912 135350 149968
rect 135406 149912 172836 149968
rect 135345 149910 172836 149912
rect 135345 149907 135411 149910
rect 172830 149908 172836 149910
rect 172900 149908 172906 149972
rect 194961 149970 195027 149973
rect 250529 149970 250595 149973
rect 194961 149968 250595 149970
rect 194961 149912 194966 149968
rect 195022 149912 250534 149968
rect 250590 149912 250595 149968
rect 194961 149910 250595 149912
rect 194961 149907 195027 149910
rect 250529 149907 250595 149910
rect 3693 149834 3759 149837
rect -960 149832 3759 149834
rect -960 149776 3698 149832
rect 3754 149776 3759 149832
rect -960 149774 3759 149776
rect -960 149684 480 149774
rect 3693 149771 3759 149774
rect 110413 149834 110479 149837
rect 170070 149834 170076 149836
rect 110413 149832 170076 149834
rect 110413 149776 110418 149832
rect 110474 149776 170076 149832
rect 110413 149774 170076 149776
rect 110413 149771 110479 149774
rect 170070 149772 170076 149774
rect 170140 149772 170146 149836
rect 177430 149772 177436 149836
rect 177500 149834 177506 149836
rect 232681 149834 232747 149837
rect 177500 149832 232747 149834
rect 177500 149776 232686 149832
rect 232742 149776 232747 149832
rect 177500 149774 232747 149776
rect 177500 149772 177506 149774
rect 232681 149771 232747 149774
rect 53833 149698 53899 149701
rect 155769 149698 155835 149701
rect 53833 149696 155835 149698
rect 53833 149640 53838 149696
rect 53894 149640 155774 149696
rect 155830 149640 155835 149696
rect 53833 149638 155835 149640
rect 53833 149635 53899 149638
rect 155769 149635 155835 149638
rect 299381 149698 299447 149701
rect 529933 149698 529999 149701
rect 299381 149696 529999 149698
rect 299381 149640 299386 149696
rect 299442 149640 529938 149696
rect 529994 149640 529999 149696
rect 299381 149638 529999 149640
rect 299381 149635 299447 149638
rect 529933 149635 529999 149638
rect 173566 149500 173572 149564
rect 173636 149562 173642 149564
rect 211153 149562 211219 149565
rect 173636 149560 211219 149562
rect 173636 149504 211158 149560
rect 211214 149504 211219 149560
rect 173636 149502 211219 149504
rect 173636 149500 173642 149502
rect 211153 149499 211219 149502
rect 173157 149154 173223 149157
rect 175958 149154 175964 149156
rect 173157 149152 175964 149154
rect 173157 149096 173162 149152
rect 173218 149096 175964 149152
rect 173157 149094 175964 149096
rect 173157 149091 173223 149094
rect 175958 149092 175964 149094
rect 176028 149092 176034 149156
rect 204713 149018 204779 149021
rect 275185 149018 275251 149021
rect 204713 149016 275251 149018
rect 204713 148960 204718 149016
rect 204774 148960 275190 149016
rect 275246 148960 275251 149016
rect 204713 148958 275251 148960
rect 204713 148955 204779 148958
rect 275185 148955 275251 148958
rect 199009 148882 199075 148885
rect 258809 148882 258875 148885
rect 199009 148880 258875 148882
rect 199009 148824 199014 148880
rect 199070 148824 258814 148880
rect 258870 148824 258875 148880
rect 199009 148822 258875 148824
rect 199009 148819 199075 148822
rect 258809 148819 258875 148822
rect 199469 148746 199535 148749
rect 256049 148746 256115 148749
rect 199469 148744 256115 148746
rect 199469 148688 199474 148744
rect 199530 148688 256054 148744
rect 256110 148688 256115 148744
rect 199469 148686 256115 148688
rect 199469 148683 199535 148686
rect 256049 148683 256115 148686
rect 178718 148548 178724 148612
rect 178788 148610 178794 148612
rect 215845 148610 215911 148613
rect 178788 148608 215911 148610
rect 178788 148552 215850 148608
rect 215906 148552 215911 148608
rect 178788 148550 215911 148552
rect 178788 148548 178794 148550
rect 215845 148547 215911 148550
rect 136633 148474 136699 148477
rect 173566 148474 173572 148476
rect 136633 148472 173572 148474
rect 136633 148416 136638 148472
rect 136694 148416 173572 148472
rect 136633 148414 173572 148416
rect 136633 148411 136699 148414
rect 173566 148412 173572 148414
rect 173636 148412 173642 148476
rect 75913 148338 75979 148341
rect 158253 148338 158319 148341
rect 75913 148336 158319 148338
rect 75913 148280 75918 148336
rect 75974 148280 158258 148336
rect 158314 148280 158319 148336
rect 75913 148278 158319 148280
rect 75913 148275 75979 148278
rect 158253 148275 158319 148278
rect 275185 148338 275251 148341
rect 543733 148338 543799 148341
rect 275185 148336 543799 148338
rect 275185 148280 275190 148336
rect 275246 148280 543738 148336
rect 543794 148280 543799 148336
rect 275185 148278 543799 148280
rect 275185 148275 275251 148278
rect 543733 148275 543799 148278
rect 215293 147794 215359 147797
rect 215845 147794 215911 147797
rect 215293 147792 215911 147794
rect 215293 147736 215298 147792
rect 215354 147736 215850 147792
rect 215906 147736 215911 147792
rect 215293 147734 215911 147736
rect 215293 147731 215359 147734
rect 215845 147731 215911 147734
rect 154113 147658 154179 147661
rect 171174 147658 171180 147660
rect 142110 147656 171180 147658
rect 142110 147600 154118 147656
rect 154174 147600 171180 147656
rect 142110 147598 171180 147600
rect 120717 147114 120783 147117
rect 142110 147114 142170 147598
rect 154113 147595 154179 147598
rect 171174 147596 171180 147598
rect 171244 147596 171250 147660
rect 206553 147658 206619 147661
rect 265566 147658 265572 147660
rect 206553 147656 265572 147658
rect 206553 147600 206558 147656
rect 206614 147600 265572 147656
rect 206553 147598 265572 147600
rect 206553 147595 206619 147598
rect 265566 147596 265572 147598
rect 265636 147596 265642 147660
rect 153101 147522 153167 147525
rect 169886 147522 169892 147524
rect 120717 147112 142170 147114
rect 120717 147056 120722 147112
rect 120778 147056 142170 147112
rect 120717 147054 142170 147056
rect 151770 147520 169892 147522
rect 151770 147464 153106 147520
rect 153162 147464 169892 147520
rect 151770 147462 169892 147464
rect 120717 147051 120783 147054
rect 103513 146978 103579 146981
rect 151770 146978 151830 147462
rect 153101 147459 153167 147462
rect 169886 147460 169892 147462
rect 169956 147460 169962 147524
rect 174486 147460 174492 147524
rect 174556 147522 174562 147524
rect 233734 147522 233740 147524
rect 174556 147462 233740 147522
rect 174556 147460 174562 147462
rect 233734 147460 233740 147462
rect 233804 147460 233810 147524
rect 173750 147324 173756 147388
rect 173820 147386 173826 147388
rect 213361 147386 213427 147389
rect 173820 147384 213427 147386
rect 173820 147328 213366 147384
rect 213422 147328 213427 147384
rect 173820 147326 213427 147328
rect 173820 147324 173826 147326
rect 213361 147323 213427 147326
rect 177614 147188 177620 147252
rect 177684 147250 177690 147252
rect 214741 147250 214807 147253
rect 177684 147248 214807 147250
rect 177684 147192 214746 147248
rect 214802 147192 214807 147248
rect 177684 147190 214807 147192
rect 177684 147188 177690 147190
rect 214741 147187 214807 147190
rect 196341 147114 196407 147117
rect 232446 147114 232452 147116
rect 196341 147112 232452 147114
rect 196341 147056 196346 147112
rect 196402 147056 232452 147112
rect 196341 147054 232452 147056
rect 196341 147051 196407 147054
rect 232446 147052 232452 147054
rect 232516 147052 232522 147116
rect 103513 146976 151830 146978
rect 103513 146920 103518 146976
rect 103574 146920 151830 146976
rect 103513 146918 151830 146920
rect 103513 146915 103579 146918
rect 202638 146236 202644 146300
rect 202708 146298 202714 146300
rect 262806 146298 262812 146300
rect 202708 146238 262812 146298
rect 202708 146236 202714 146238
rect 262806 146236 262812 146238
rect 262876 146236 262882 146300
rect 201350 146100 201356 146164
rect 201420 146162 201426 146164
rect 260925 146162 260991 146165
rect 201420 146160 260991 146162
rect 201420 146104 260930 146160
rect 260986 146104 260991 146160
rect 201420 146102 260991 146104
rect 201420 146100 201426 146102
rect 260925 146099 260991 146102
rect 203742 145964 203748 146028
rect 203812 146026 203818 146028
rect 262254 146026 262260 146028
rect 203812 145966 262260 146026
rect 203812 145964 203818 145966
rect 262254 145964 262260 145966
rect 262324 145964 262330 146028
rect 202454 145828 202460 145892
rect 202524 145890 202530 145892
rect 261150 145890 261156 145892
rect 202524 145830 261156 145890
rect 202524 145828 202530 145830
rect 261150 145828 261156 145830
rect 261220 145828 261226 145892
rect 205030 145692 205036 145756
rect 205100 145754 205106 145756
rect 231301 145754 231367 145757
rect 205100 145752 231367 145754
rect 205100 145696 231306 145752
rect 231362 145696 231367 145752
rect 205100 145694 231367 145696
rect 205100 145692 205106 145694
rect 231301 145691 231367 145694
rect 18597 145618 18663 145621
rect 163078 145618 163084 145620
rect 18597 145616 163084 145618
rect 18597 145560 18602 145616
rect 18658 145560 163084 145616
rect 18597 145558 163084 145560
rect 18597 145555 18663 145558
rect 163078 145556 163084 145558
rect 163148 145556 163154 145620
rect 160093 144802 160159 144805
rect 161381 144802 161447 144805
rect 235206 144802 235212 144804
rect 160093 144800 235212 144802
rect 160093 144744 160098 144800
rect 160154 144744 161386 144800
rect 161442 144744 235212 144800
rect 160093 144742 235212 144744
rect 160093 144739 160159 144742
rect 161381 144739 161447 144742
rect 235206 144740 235212 144742
rect 235276 144740 235282 144804
rect 186998 144604 187004 144668
rect 187068 144666 187074 144668
rect 211889 144666 211955 144669
rect 187068 144664 211955 144666
rect 187068 144608 211894 144664
rect 211950 144608 211955 144664
rect 187068 144606 211955 144608
rect 187068 144604 187074 144606
rect 211889 144603 211955 144606
rect 171542 144530 171548 144532
rect 161430 144470 171548 144530
rect 117957 144122 118023 144125
rect 161430 144122 161490 144470
rect 171542 144468 171548 144470
rect 171612 144530 171618 144532
rect 230974 144530 230980 144532
rect 171612 144470 230980 144530
rect 171612 144468 171618 144470
rect 230974 144468 230980 144470
rect 231044 144468 231050 144532
rect 196198 144332 196204 144396
rect 196268 144394 196274 144396
rect 197077 144394 197143 144397
rect 196268 144392 197143 144394
rect 196268 144336 197082 144392
rect 197138 144336 197143 144392
rect 196268 144334 197143 144336
rect 196268 144332 196274 144334
rect 197077 144331 197143 144334
rect 200614 144332 200620 144396
rect 200684 144394 200690 144396
rect 201217 144394 201283 144397
rect 200684 144392 201283 144394
rect 200684 144336 201222 144392
rect 201278 144336 201283 144392
rect 200684 144334 201283 144336
rect 200684 144332 200690 144334
rect 201217 144331 201283 144334
rect 202086 144332 202092 144396
rect 202156 144394 202162 144396
rect 202689 144394 202755 144397
rect 202156 144392 202755 144394
rect 202156 144336 202694 144392
rect 202750 144336 202755 144392
rect 202156 144334 202755 144336
rect 202156 144332 202162 144334
rect 202689 144331 202755 144334
rect 203701 144394 203767 144397
rect 259678 144394 259684 144396
rect 203701 144392 259684 144394
rect 203701 144336 203706 144392
rect 203762 144336 259684 144392
rect 203701 144334 259684 144336
rect 203701 144331 203767 144334
rect 259678 144332 259684 144334
rect 259748 144332 259754 144396
rect 238109 144258 238175 144261
rect 117957 144120 161490 144122
rect 117957 144064 117962 144120
rect 118018 144064 161490 144120
rect 117957 144062 161490 144064
rect 200070 144256 238175 144258
rect 200070 144200 238114 144256
rect 238170 144200 238175 144256
rect 200070 144198 238175 144200
rect 117957 144059 118023 144062
rect 199510 143924 199516 143988
rect 199580 143986 199586 143988
rect 199878 143986 199884 143988
rect 199580 143926 199884 143986
rect 199580 143924 199586 143926
rect 199878 143924 199884 143926
rect 199948 143986 199954 143988
rect 200070 143986 200130 144198
rect 238109 144195 238175 144198
rect 200205 144122 200271 144125
rect 201125 144122 201191 144125
rect 200205 144120 202154 144122
rect 200205 144064 200210 144120
rect 200266 144064 201130 144120
rect 201186 144064 202154 144120
rect 200205 144062 202154 144064
rect 200205 144059 200271 144062
rect 201125 144059 201191 144062
rect 199948 143926 200130 143986
rect 202094 143986 202154 144062
rect 202270 144060 202276 144124
rect 202340 144122 202346 144124
rect 238293 144122 238359 144125
rect 202340 144120 238359 144122
rect 202340 144064 238298 144120
rect 238354 144064 238359 144120
rect 202340 144062 238359 144064
rect 202340 144060 202346 144062
rect 238293 144059 238359 144062
rect 203701 143986 203767 143989
rect 202094 143984 203767 143986
rect 202094 143928 203706 143984
rect 203762 143928 203767 143984
rect 202094 143926 203767 143928
rect 199948 143924 199954 143926
rect 203701 143923 203767 143926
rect 201166 143788 201172 143852
rect 201236 143850 201242 143852
rect 261334 143850 261340 143852
rect 201236 143790 261340 143850
rect 201236 143788 201242 143790
rect 261334 143788 261340 143790
rect 261404 143788 261410 143852
rect 189758 143380 189764 143444
rect 189828 143442 189834 143444
rect 248454 143442 248460 143444
rect 189828 143382 248460 143442
rect 189828 143380 189834 143382
rect 248454 143380 248460 143382
rect 248524 143380 248530 143444
rect 189942 143244 189948 143308
rect 190012 143306 190018 143308
rect 246389 143306 246455 143309
rect 190012 143304 246455 143306
rect 190012 143248 246394 143304
rect 246450 143248 246455 143304
rect 190012 143246 246455 143248
rect 190012 143244 190018 143246
rect 246389 143243 246455 143246
rect 187182 143108 187188 143172
rect 187252 143170 187258 143172
rect 242014 143170 242020 143172
rect 187252 143110 242020 143170
rect 187252 143108 187258 143110
rect 242014 143108 242020 143110
rect 242084 143108 242090 143172
rect 187366 142972 187372 143036
rect 187436 143034 187442 143036
rect 236729 143034 236795 143037
rect 187436 143032 236795 143034
rect 187436 142976 236734 143032
rect 236790 142976 236795 143032
rect 187436 142974 236795 142976
rect 187436 142972 187442 142974
rect 236729 142971 236795 142974
rect 188654 142836 188660 142900
rect 188724 142898 188730 142900
rect 228449 142898 228515 142901
rect 188724 142896 228515 142898
rect 188724 142840 228454 142896
rect 228510 142840 228515 142896
rect 188724 142838 228515 142840
rect 188724 142836 188730 142838
rect 228449 142835 228515 142838
rect 255313 142898 255379 142901
rect 255814 142898 255820 142900
rect 255313 142896 255820 142898
rect 255313 142840 255318 142896
rect 255374 142840 255820 142896
rect 255313 142838 255820 142840
rect 255313 142835 255379 142838
rect 255814 142836 255820 142838
rect 255884 142836 255890 142900
rect 185158 142700 185164 142764
rect 185228 142762 185234 142764
rect 224217 142762 224283 142765
rect 185228 142760 224283 142762
rect 185228 142704 224222 142760
rect 224278 142704 224283 142760
rect 185228 142702 224283 142704
rect 185228 142700 185234 142702
rect 224217 142699 224283 142702
rect 187550 142564 187556 142628
rect 187620 142626 187626 142628
rect 225781 142626 225847 142629
rect 187620 142624 225847 142626
rect 187620 142568 225786 142624
rect 225842 142568 225847 142624
rect 187620 142566 225847 142568
rect 187620 142564 187626 142566
rect 225781 142563 225847 142566
rect 181478 142020 181484 142084
rect 181548 142082 181554 142084
rect 242249 142082 242315 142085
rect 181548 142080 242315 142082
rect 181548 142024 242254 142080
rect 242310 142024 242315 142080
rect 181548 142022 242315 142024
rect 181548 142020 181554 142022
rect 242249 142019 242315 142022
rect 181110 141884 181116 141948
rect 181180 141946 181186 141948
rect 240726 141946 240732 141948
rect 181180 141886 240732 141946
rect 181180 141884 181186 141886
rect 240726 141884 240732 141886
rect 240796 141884 240802 141948
rect 183134 141748 183140 141812
rect 183204 141810 183210 141812
rect 238702 141810 238708 141812
rect 183204 141750 238708 141810
rect 183204 141748 183210 141750
rect 238702 141748 238708 141750
rect 238772 141748 238778 141812
rect 267917 141810 267983 141813
rect 268326 141810 268332 141812
rect 267917 141808 268332 141810
rect 267917 141752 267922 141808
rect 267978 141752 268332 141808
rect 267917 141750 268332 141752
rect 267917 141747 267983 141750
rect 268326 141748 268332 141750
rect 268396 141748 268402 141812
rect 188470 141612 188476 141676
rect 188540 141674 188546 141676
rect 239489 141674 239555 141677
rect 188540 141672 239555 141674
rect 188540 141616 239494 141672
rect 239550 141616 239555 141672
rect 188540 141614 239555 141616
rect 188540 141612 188546 141614
rect 239489 141611 239555 141614
rect 177798 141476 177804 141540
rect 177868 141538 177874 141540
rect 189717 141538 189783 141541
rect 177868 141536 189783 141538
rect 177868 141480 189722 141536
rect 189778 141480 189783 141536
rect 177868 141478 189783 141480
rect 177868 141476 177874 141478
rect 189717 141475 189783 141478
rect 192886 141476 192892 141540
rect 192956 141538 192962 141540
rect 236637 141538 236703 141541
rect 192956 141536 236703 141538
rect 192956 141480 236642 141536
rect 236698 141480 236703 141536
rect 192956 141478 236703 141480
rect 192956 141476 192962 141478
rect 236637 141475 236703 141478
rect 147673 141402 147739 141405
rect 174486 141402 174492 141404
rect 147673 141400 174492 141402
rect 147673 141344 147678 141400
rect 147734 141344 174492 141400
rect 147673 141342 174492 141344
rect 147673 141339 147739 141342
rect 174486 141340 174492 141342
rect 174556 141340 174562 141404
rect 177798 141340 177804 141404
rect 177868 141402 177874 141404
rect 217409 141402 217475 141405
rect 177868 141400 217475 141402
rect 177868 141344 217414 141400
rect 217470 141344 217475 141400
rect 177868 141342 217475 141344
rect 177868 141340 177874 141342
rect 217409 141339 217475 141342
rect 186129 141266 186195 141269
rect 220077 141266 220143 141269
rect 186129 141264 220143 141266
rect 186129 141208 186134 141264
rect 186190 141208 220082 141264
rect 220138 141208 220143 141264
rect 186129 141206 220143 141208
rect 186129 141203 186195 141206
rect 220077 141203 220143 141206
rect 177246 140796 177252 140860
rect 177316 140858 177322 140860
rect 177798 140858 177804 140860
rect 177316 140798 177804 140858
rect 177316 140796 177322 140798
rect 177798 140796 177804 140798
rect 177868 140796 177874 140860
rect 184974 140796 184980 140860
rect 185044 140858 185050 140860
rect 186129 140858 186195 140861
rect 185044 140856 186195 140858
rect 185044 140800 186134 140856
rect 186190 140800 186195 140856
rect 185044 140798 186195 140800
rect 185044 140796 185050 140798
rect 186129 140795 186195 140798
rect 198222 140660 198228 140724
rect 198292 140722 198298 140724
rect 258533 140722 258599 140725
rect 198292 140720 258599 140722
rect 198292 140664 258538 140720
rect 258594 140664 258599 140720
rect 198292 140662 258599 140664
rect 198292 140660 198298 140662
rect 258533 140659 258599 140662
rect 168230 140524 168236 140588
rect 168300 140586 168306 140588
rect 225873 140586 225939 140589
rect 168300 140584 225939 140586
rect 168300 140528 225878 140584
rect 225934 140528 225939 140584
rect 168300 140526 225939 140528
rect 168300 140524 168306 140526
rect 225873 140523 225939 140526
rect 140773 140042 140839 140045
rect 173014 140042 173020 140044
rect 140773 140040 173020 140042
rect 140773 139984 140778 140040
rect 140834 139984 173020 140040
rect 140773 139982 173020 139984
rect 140773 139979 140839 139982
rect 173014 139980 173020 139982
rect 173084 139980 173090 140044
rect 179086 139980 179092 140044
rect 179156 140042 179162 140044
rect 216673 140042 216739 140045
rect 179156 140040 216739 140042
rect 179156 139984 216678 140040
rect 216734 139984 216739 140040
rect 179156 139982 216739 139984
rect 179156 139980 179162 139982
rect 216673 139979 216739 139982
rect 197537 139362 197603 139365
rect 198641 139362 198707 139365
rect 204713 139362 204779 139365
rect 262857 139362 262923 139365
rect 197537 139360 204779 139362
rect 197537 139304 197542 139360
rect 197598 139304 198646 139360
rect 198702 139304 204718 139360
rect 204774 139304 204779 139360
rect 197537 139302 204779 139304
rect 197537 139299 197603 139302
rect 198641 139299 198707 139302
rect 204713 139299 204779 139302
rect 204854 139360 262923 139362
rect 204854 139304 262862 139360
rect 262918 139304 262923 139360
rect 204854 139302 262923 139304
rect 194358 139164 194364 139228
rect 194428 139226 194434 139228
rect 204854 139226 204914 139302
rect 262857 139299 262923 139302
rect 580257 139362 580323 139365
rect 583520 139362 584960 139452
rect 580257 139360 584960 139362
rect 580257 139304 580262 139360
rect 580318 139304 584960 139360
rect 580257 139302 584960 139304
rect 580257 139299 580323 139302
rect 194428 139166 204914 139226
rect 204989 139226 205055 139229
rect 257102 139226 257108 139228
rect 204989 139224 257108 139226
rect 204989 139168 204994 139224
rect 205050 139168 257108 139224
rect 204989 139166 257108 139168
rect 194428 139164 194434 139166
rect 204989 139163 205055 139166
rect 257102 139164 257108 139166
rect 257172 139164 257178 139228
rect 583520 139212 584960 139302
rect 195462 139028 195468 139092
rect 195532 139090 195538 139092
rect 254894 139090 254900 139092
rect 195532 139030 254900 139090
rect 195532 139028 195538 139030
rect 254894 139028 254900 139030
rect 254964 139028 254970 139092
rect 191230 138892 191236 138956
rect 191300 138954 191306 138956
rect 231209 138954 231275 138957
rect 191300 138952 231275 138954
rect 191300 138896 231214 138952
rect 231270 138896 231275 138952
rect 191300 138894 231275 138896
rect 191300 138892 191306 138894
rect 231209 138891 231275 138894
rect 190126 138756 190132 138820
rect 190196 138818 190202 138820
rect 229737 138818 229803 138821
rect 190196 138816 229803 138818
rect 190196 138760 229742 138816
rect 229798 138760 229803 138816
rect 190196 138758 229803 138760
rect 190196 138756 190202 138758
rect 229737 138755 229803 138758
rect 193990 138620 193996 138684
rect 194060 138682 194066 138684
rect 232589 138682 232655 138685
rect 194060 138680 232655 138682
rect 194060 138624 232594 138680
rect 232650 138624 232655 138680
rect 194060 138622 232655 138624
rect 194060 138620 194066 138622
rect 232589 138619 232655 138622
rect 192702 138484 192708 138548
rect 192772 138546 192778 138548
rect 223021 138546 223087 138549
rect 192772 138544 223087 138546
rect 192772 138488 223026 138544
rect 223082 138488 223087 138544
rect 192772 138486 223087 138488
rect 192772 138484 192778 138486
rect 223021 138483 223087 138486
rect 271822 137940 271828 138004
rect 271892 138002 271898 138004
rect 272241 138002 272307 138005
rect 271892 138000 272307 138002
rect 271892 137944 272246 138000
rect 272302 137944 272307 138000
rect 271892 137942 272307 137944
rect 271892 137940 271898 137942
rect 272241 137939 272307 137942
rect 59353 137322 59419 137325
rect 168230 137322 168236 137324
rect 59353 137320 168236 137322
rect 59353 137264 59358 137320
rect 59414 137264 168236 137320
rect 59353 137262 168236 137264
rect 59353 137259 59419 137262
rect 168230 137260 168236 137262
rect 168300 137260 168306 137324
rect -960 136778 480 136868
rect 3601 136778 3667 136781
rect -960 136776 3667 136778
rect -960 136720 3606 136776
rect 3662 136720 3667 136776
rect -960 136718 3667 136720
rect -960 136628 480 136718
rect 3601 136715 3667 136718
rect 128997 136098 129063 136101
rect 171726 136098 171732 136100
rect 128997 136096 171732 136098
rect 128997 136040 129002 136096
rect 129058 136040 171732 136096
rect 128997 136038 171732 136040
rect 128997 136035 129063 136038
rect 171726 136036 171732 136038
rect 171796 136036 171802 136100
rect 80697 135962 80763 135965
rect 168966 135962 168972 135964
rect 80697 135960 168972 135962
rect 80697 135904 80702 135960
rect 80758 135904 168972 135960
rect 80697 135902 168972 135904
rect 80697 135899 80763 135902
rect 168966 135900 168972 135902
rect 169036 135900 169042 135964
rect 55213 131746 55279 131749
rect 165654 131746 165660 131748
rect 55213 131744 165660 131746
rect 55213 131688 55218 131744
rect 55274 131688 165660 131744
rect 55213 131686 165660 131688
rect 55213 131683 55279 131686
rect 165654 131684 165660 131686
rect 165724 131684 165730 131748
rect 84193 130522 84259 130525
rect 168598 130522 168604 130524
rect 84193 130520 168604 130522
rect 84193 130464 84198 130520
rect 84254 130464 168604 130520
rect 84193 130462 168604 130464
rect 84193 130459 84259 130462
rect 168598 130460 168604 130462
rect 168668 130460 168674 130524
rect 36537 130386 36603 130389
rect 164366 130386 164372 130388
rect 36537 130384 164372 130386
rect 36537 130328 36542 130384
rect 36598 130328 164372 130384
rect 36537 130326 164372 130328
rect 36537 130323 36603 130326
rect 164366 130324 164372 130326
rect 164436 130324 164442 130388
rect 182950 130324 182956 130388
rect 183020 130386 183026 130388
rect 259545 130386 259611 130389
rect 183020 130384 259611 130386
rect 183020 130328 259550 130384
rect 259606 130328 259611 130384
rect 183020 130326 259611 130328
rect 183020 130324 183026 130326
rect 259545 130323 259611 130326
rect 182582 127604 182588 127668
rect 182652 127666 182658 127668
rect 255313 127666 255379 127669
rect 182652 127664 255379 127666
rect 182652 127608 255318 127664
rect 255374 127608 255379 127664
rect 182652 127606 255379 127608
rect 182652 127604 182658 127606
rect 255313 127603 255379 127606
rect 129733 126442 129799 126445
rect 172462 126442 172468 126444
rect 129733 126440 172468 126442
rect 129733 126384 129738 126440
rect 129794 126384 172468 126440
rect 129733 126382 172468 126384
rect 129733 126379 129799 126382
rect 172462 126380 172468 126382
rect 172532 126380 172538 126444
rect 80053 126306 80119 126309
rect 168414 126306 168420 126308
rect 80053 126304 168420 126306
rect 80053 126248 80058 126304
rect 80114 126248 168420 126304
rect 80053 126246 168420 126248
rect 80053 126243 80119 126246
rect 168414 126244 168420 126246
rect 168484 126244 168490 126308
rect 580533 126034 580599 126037
rect 583520 126034 584960 126124
rect 580533 126032 584960 126034
rect 580533 125976 580538 126032
rect 580594 125976 584960 126032
rect 580533 125974 584960 125976
rect 580533 125971 580599 125974
rect 583520 125884 584960 125974
rect 180374 124748 180380 124812
rect 180444 124810 180450 124812
rect 230473 124810 230539 124813
rect 180444 124808 230539 124810
rect 180444 124752 230478 124808
rect 230534 124752 230539 124808
rect 180444 124750 230539 124752
rect 180444 124748 180450 124750
rect 230473 124747 230539 124750
rect -960 123572 480 123812
rect 112437 122226 112503 122229
rect 169702 122226 169708 122228
rect 112437 122224 169708 122226
rect 112437 122168 112442 122224
rect 112498 122168 169708 122224
rect 112437 122166 169708 122168
rect 112437 122163 112503 122166
rect 169702 122164 169708 122166
rect 169772 122164 169778 122228
rect 181110 122164 181116 122228
rect 181180 122226 181186 122228
rect 244273 122226 244339 122229
rect 181180 122224 244339 122226
rect 181180 122168 244278 122224
rect 244334 122168 244339 122224
rect 181180 122166 244339 122168
rect 181180 122164 181186 122166
rect 244273 122163 244339 122166
rect 20713 122090 20779 122093
rect 162894 122090 162900 122092
rect 20713 122088 162900 122090
rect 20713 122032 20718 122088
rect 20774 122032 162900 122088
rect 20713 122030 162900 122032
rect 20713 122027 20779 122030
rect 162894 122028 162900 122030
rect 162964 122028 162970 122092
rect 203742 122028 203748 122092
rect 203812 122090 203818 122092
rect 520917 122090 520983 122093
rect 203812 122088 520983 122090
rect 203812 122032 520922 122088
rect 520978 122032 520983 122088
rect 203812 122030 520983 122032
rect 203812 122028 203818 122030
rect 520917 122027 520983 122030
rect 180006 120940 180012 121004
rect 180076 121002 180082 121004
rect 226425 121002 226491 121005
rect 180076 121000 226491 121002
rect 180076 120944 226430 121000
rect 226486 120944 226491 121000
rect 180076 120942 226491 120944
rect 180076 120940 180082 120942
rect 226425 120939 226491 120942
rect 195278 120804 195284 120868
rect 195348 120866 195354 120868
rect 426433 120866 426499 120869
rect 195348 120864 426499 120866
rect 195348 120808 426438 120864
rect 426494 120808 426499 120864
rect 195348 120806 426499 120808
rect 195348 120804 195354 120806
rect 426433 120803 426499 120806
rect 205030 120668 205036 120732
rect 205100 120730 205106 120732
rect 539593 120730 539659 120733
rect 205100 120728 539659 120730
rect 205100 120672 539598 120728
rect 539654 120672 539659 120728
rect 205100 120670 539659 120672
rect 205100 120668 205106 120670
rect 539593 120667 539659 120670
rect 196750 117948 196756 118012
rect 196820 118010 196826 118012
rect 448605 118010 448671 118013
rect 196820 118008 448671 118010
rect 196820 117952 448610 118008
rect 448666 117952 448671 118008
rect 196820 117950 448671 117952
rect 196820 117948 196826 117950
rect 448605 117947 448671 117950
rect 177430 116452 177436 116516
rect 177500 116514 177506 116516
rect 197353 116514 197419 116517
rect 177500 116512 197419 116514
rect 177500 116456 197358 116512
rect 197414 116456 197419 116512
rect 177500 116454 197419 116456
rect 177500 116452 177506 116454
rect 197353 116451 197419 116454
rect 198038 116452 198044 116516
rect 198108 116514 198114 116516
rect 462313 116514 462379 116517
rect 198108 116512 462379 116514
rect 198108 116456 462318 116512
rect 462374 116456 462379 116512
rect 198108 116454 462379 116456
rect 198108 116452 198114 116454
rect 462313 116451 462379 116454
rect 199694 115092 199700 115156
rect 199764 115154 199770 115156
rect 472617 115154 472683 115157
rect 199764 115152 472683 115154
rect 199764 115096 472622 115152
rect 472678 115096 472683 115152
rect 199764 115094 472683 115096
rect 199764 115092 199770 115094
rect 472617 115091 472683 115094
rect 44265 113794 44331 113797
rect 165838 113794 165844 113796
rect 44265 113792 165844 113794
rect 44265 113736 44270 113792
rect 44326 113736 165844 113792
rect 44265 113734 165844 113736
rect 44265 113731 44331 113734
rect 165838 113732 165844 113734
rect 165908 113732 165914 113796
rect 189758 113732 189764 113796
rect 189828 113794 189834 113796
rect 343633 113794 343699 113797
rect 189828 113792 343699 113794
rect 189828 113736 343638 113792
rect 343694 113736 343699 113792
rect 189828 113734 343699 113736
rect 189828 113732 189834 113734
rect 343633 113731 343699 113734
rect 580165 112842 580231 112845
rect 583520 112842 584960 112932
rect 580165 112840 584960 112842
rect 580165 112784 580170 112840
rect 580226 112784 584960 112840
rect 580165 112782 584960 112784
rect 580165 112779 580231 112782
rect 583520 112692 584960 112782
rect 180742 112372 180748 112436
rect 180812 112434 180818 112436
rect 247677 112434 247743 112437
rect 180812 112432 247743 112434
rect 180812 112376 247682 112432
rect 247738 112376 247743 112432
rect 180812 112374 247743 112376
rect 180812 112372 180818 112374
rect 247677 112371 247743 112374
rect 200982 111012 200988 111076
rect 201052 111074 201058 111076
rect 485773 111074 485839 111077
rect 201052 111072 485839 111074
rect 201052 111016 485778 111072
rect 485834 111016 485839 111072
rect 201052 111014 485839 111016
rect 201052 111012 201058 111014
rect 485773 111011 485839 111014
rect -960 110666 480 110756
rect 3141 110666 3207 110669
rect -960 110664 3207 110666
rect -960 110608 3146 110664
rect 3202 110608 3207 110664
rect -960 110606 3207 110608
rect -960 110516 480 110606
rect 3141 110603 3207 110606
rect 184606 109652 184612 109716
rect 184676 109714 184682 109716
rect 276105 109714 276171 109717
rect 184676 109712 276171 109714
rect 184676 109656 276110 109712
rect 276166 109656 276171 109712
rect 184676 109654 276171 109656
rect 184676 109652 184682 109654
rect 276105 109651 276171 109654
rect 184422 108292 184428 108356
rect 184492 108354 184498 108356
rect 280153 108354 280219 108357
rect 184492 108352 280219 108354
rect 184492 108296 280158 108352
rect 280214 108296 280219 108352
rect 184492 108294 280219 108296
rect 184492 108292 184498 108294
rect 280153 108291 280219 108294
rect 186998 106932 187004 106996
rect 187068 106994 187074 106996
rect 311893 106994 311959 106997
rect 187068 106992 311959 106994
rect 187068 106936 311898 106992
rect 311954 106936 311959 106992
rect 187068 106934 311959 106936
rect 187068 106932 187074 106934
rect 311893 106931 311959 106934
rect 201166 106796 201172 106860
rect 201236 106858 201242 106860
rect 496813 106858 496879 106861
rect 201236 106856 496879 106858
rect 201236 106800 496818 106856
rect 496874 106800 496879 106856
rect 201236 106798 496879 106800
rect 201236 106796 201242 106798
rect 496813 106795 496879 106798
rect 202270 105436 202276 105500
rect 202340 105498 202346 105500
rect 506565 105498 506631 105501
rect 202340 105496 506631 105498
rect 202340 105440 506570 105496
rect 506626 105440 506631 105496
rect 202340 105438 506631 105440
rect 202340 105436 202346 105438
rect 506565 105435 506631 105438
rect 202454 104076 202460 104140
rect 202524 104138 202530 104140
rect 510613 104138 510679 104141
rect 202524 104136 510679 104138
rect 202524 104080 510618 104136
rect 510674 104080 510679 104136
rect 202524 104078 510679 104080
rect 202524 104076 202530 104078
rect 510613 104075 510679 104078
rect 191046 102852 191052 102916
rect 191116 102914 191122 102916
rect 365805 102914 365871 102917
rect 191116 102912 365871 102914
rect 191116 102856 365810 102912
rect 365866 102856 365871 102912
rect 191116 102854 365871 102856
rect 191116 102852 191122 102854
rect 365805 102851 365871 102854
rect 202638 102716 202644 102780
rect 202708 102778 202714 102780
rect 514845 102778 514911 102781
rect 202708 102776 514911 102778
rect 202708 102720 514850 102776
rect 514906 102720 514911 102776
rect 202708 102718 514911 102720
rect 202708 102716 202714 102718
rect 514845 102715 514911 102718
rect 187182 100132 187188 100196
rect 187252 100194 187258 100196
rect 315297 100194 315363 100197
rect 187252 100192 315363 100194
rect 187252 100136 315302 100192
rect 315358 100136 315363 100192
rect 187252 100134 315363 100136
rect 187252 100132 187258 100134
rect 315297 100131 315363 100134
rect 161974 99996 161980 100060
rect 162044 100058 162050 100060
rect 580257 100058 580323 100061
rect 162044 100056 580323 100058
rect 162044 100000 580262 100056
rect 580318 100000 580323 100056
rect 162044 99998 580323 100000
rect 162044 99996 162050 99998
rect 580257 99995 580323 99998
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect 179822 98772 179828 98836
rect 179892 98834 179898 98836
rect 234705 98834 234771 98837
rect 179892 98832 234771 98834
rect 179892 98776 234710 98832
rect 234766 98776 234771 98832
rect 179892 98774 234771 98776
rect 179892 98772 179898 98774
rect 234705 98771 234771 98774
rect 176510 98636 176516 98700
rect 176580 98698 176586 98700
rect 179413 98698 179479 98701
rect 176580 98696 179479 98698
rect 176580 98640 179418 98696
rect 179474 98640 179479 98696
rect 176580 98638 179479 98640
rect 176580 98636 176586 98638
rect 179413 98635 179479 98638
rect 203190 98636 203196 98700
rect 203260 98698 203266 98700
rect 528553 98698 528619 98701
rect 203260 98696 528619 98698
rect 203260 98640 528558 98696
rect 528614 98640 528619 98696
rect 203260 98638 528619 98640
rect 203260 98636 203266 98638
rect 528553 98635 528619 98638
rect -960 97610 480 97700
rect 3509 97610 3575 97613
rect -960 97608 3575 97610
rect -960 97552 3514 97608
rect 3570 97552 3575 97608
rect -960 97550 3575 97552
rect -960 97460 480 97550
rect 3509 97547 3575 97550
rect 183134 97276 183140 97340
rect 183204 97338 183210 97340
rect 265617 97338 265683 97341
rect 183204 97336 265683 97338
rect 183204 97280 265622 97336
rect 265678 97280 265683 97336
rect 183204 97278 265683 97280
rect 183204 97276 183210 97278
rect 265617 97275 265683 97278
rect 204110 97140 204116 97204
rect 204180 97202 204186 97204
rect 531405 97202 531471 97205
rect 204180 97200 531471 97202
rect 204180 97144 531410 97200
rect 531466 97144 531471 97200
rect 204180 97142 531471 97144
rect 204180 97140 204186 97142
rect 531405 97139 531471 97142
rect 181478 95916 181484 95980
rect 181548 95978 181554 95980
rect 251265 95978 251331 95981
rect 181548 95976 251331 95978
rect 181548 95920 251270 95976
rect 251326 95920 251331 95976
rect 181548 95918 251331 95920
rect 181548 95916 181554 95918
rect 251265 95915 251331 95918
rect 205214 95780 205220 95844
rect 205284 95842 205290 95844
rect 542353 95842 542419 95845
rect 205284 95840 542419 95842
rect 205284 95784 542358 95840
rect 542414 95784 542419 95840
rect 205284 95782 542419 95784
rect 205284 95780 205290 95782
rect 542353 95779 542419 95782
rect 184054 94420 184060 94484
rect 184124 94482 184130 94484
rect 284385 94482 284451 94485
rect 184124 94480 284451 94482
rect 184124 94424 284390 94480
rect 284446 94424 284451 94480
rect 184124 94422 284451 94424
rect 184124 94420 184130 94422
rect 284385 94419 284451 94422
rect 205398 93060 205404 93124
rect 205468 93122 205474 93124
rect 549253 93122 549319 93125
rect 205468 93120 549319 93122
rect 205468 93064 549258 93120
rect 549314 93064 549319 93120
rect 205468 93062 549319 93064
rect 205468 93060 205474 93062
rect 549253 93059 549319 93062
rect 580257 86186 580323 86189
rect 583520 86186 584960 86276
rect 580257 86184 584960 86186
rect 580257 86128 580262 86184
rect 580318 86128 584960 86184
rect 580257 86126 584960 86128
rect 580257 86123 580323 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3509 84690 3575 84693
rect -960 84688 3575 84690
rect -960 84632 3514 84688
rect 3570 84632 3575 84688
rect -960 84630 3575 84632
rect -960 84540 480 84630
rect 3509 84627 3575 84630
rect 193806 82044 193812 82108
rect 193876 82106 193882 82108
rect 400213 82106 400279 82109
rect 193876 82104 400279 82106
rect 193876 82048 400218 82104
rect 400274 82048 400279 82104
rect 193876 82046 400279 82048
rect 193876 82044 193882 82046
rect 400213 82043 400279 82046
rect 198222 76468 198228 76532
rect 198292 76530 198298 76532
rect 460933 76530 460999 76533
rect 198292 76528 460999 76530
rect 198292 76472 460938 76528
rect 460994 76472 460999 76528
rect 198292 76470 460999 76472
rect 198292 76468 198298 76470
rect 460933 76467 460999 76470
rect 583520 72994 584960 73084
rect 583342 72934 584960 72994
rect 583342 72858 583402 72934
rect 583520 72858 584960 72934
rect 583342 72844 584960 72858
rect 583342 72798 583586 72844
rect 188286 72388 188292 72452
rect 188356 72450 188362 72452
rect 340965 72450 341031 72453
rect 188356 72448 341031 72450
rect 188356 72392 340970 72448
rect 341026 72392 341031 72448
rect 188356 72390 341031 72392
rect 188356 72388 188362 72390
rect 340965 72387 341031 72390
rect 281390 71844 281396 71908
rect 281460 71906 281466 71908
rect 583526 71906 583586 72798
rect 281460 71846 583586 71906
rect 281460 71844 281466 71846
rect -960 71634 480 71724
rect 3509 71634 3575 71637
rect -960 71632 3575 71634
rect -960 71576 3514 71632
rect 3570 71576 3575 71632
rect -960 71574 3575 71576
rect -960 71484 480 71574
rect 3509 71571 3575 71574
rect 162710 71028 162716 71092
rect 162780 71090 162786 71092
rect 580257 71090 580323 71093
rect 162780 71088 580323 71090
rect 162780 71032 580262 71088
rect 580318 71032 580323 71088
rect 162780 71030 580323 71032
rect 162780 71028 162786 71030
rect 580257 71027 580323 71030
rect 187366 69532 187372 69596
rect 187436 69594 187442 69596
rect 318057 69594 318123 69597
rect 187436 69592 318123 69594
rect 187436 69536 318062 69592
rect 318118 69536 318123 69592
rect 187436 69534 318123 69536
rect 187436 69532 187442 69534
rect 318057 69531 318123 69534
rect 189942 64092 189948 64156
rect 190012 64154 190018 64156
rect 354673 64154 354739 64157
rect 190012 64152 354739 64154
rect 190012 64096 354678 64152
rect 354734 64096 354739 64152
rect 190012 64094 354739 64096
rect 190012 64092 190018 64094
rect 354673 64091 354739 64094
rect 191230 62732 191236 62796
rect 191300 62794 191306 62796
rect 361573 62794 361639 62797
rect 191300 62792 361639 62794
rect 191300 62736 361578 62792
rect 361634 62736 361639 62792
rect 191300 62734 361639 62736
rect 191300 62732 191306 62734
rect 361573 62731 361639 62734
rect 191414 61372 191420 61436
rect 191484 61434 191490 61436
rect 368473 61434 368539 61437
rect 191484 61432 368539 61434
rect 191484 61376 368478 61432
rect 368534 61376 368539 61432
rect 191484 61374 368539 61376
rect 191484 61372 191490 61374
rect 368473 61371 368539 61374
rect 583520 59666 584960 59756
rect 567150 59606 584960 59666
rect 333094 59332 333100 59396
rect 333164 59394 333170 59396
rect 567150 59394 567210 59606
rect 583520 59516 584960 59606
rect 333164 59334 567210 59394
rect 333164 59332 333170 59334
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 190862 58516 190868 58580
rect 190932 58578 190938 58580
rect 372613 58578 372679 58581
rect 190932 58576 372679 58578
rect 190932 58520 372618 58576
rect 372674 58520 372679 58576
rect 190932 58518 372679 58520
rect 190932 58516 190938 58518
rect 372613 58515 372679 58518
rect 193990 54436 193996 54500
rect 194060 54498 194066 54500
rect 407205 54498 407271 54501
rect 194060 54496 407271 54498
rect 194060 54440 407210 54496
rect 407266 54440 407271 54496
rect 194060 54438 407271 54440
rect 194060 54436 194066 54438
rect 407205 54435 407271 54438
rect 194174 53076 194180 53140
rect 194244 53138 194250 53140
rect 411253 53138 411319 53141
rect 194244 53136 411319 53138
rect 194244 53080 411258 53136
rect 411314 53080 411319 53136
rect 194244 53078 411319 53080
rect 194244 53076 194250 53078
rect 411253 53075 411319 53078
rect 580257 46338 580323 46341
rect 583520 46338 584960 46428
rect 580257 46336 584960 46338
rect 580257 46280 580262 46336
rect 580318 46280 584960 46336
rect 580257 46278 584960 46280
rect 580257 46275 580323 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3509 45522 3575 45525
rect -960 45520 3575 45522
rect -960 45464 3514 45520
rect 3570 45464 3575 45520
rect -960 45462 3575 45464
rect -960 45372 480 45462
rect 3509 45459 3575 45462
rect 201350 39204 201356 39268
rect 201420 39266 201426 39268
rect 487153 39266 487219 39269
rect 201420 39264 487219 39266
rect 201420 39208 487158 39264
rect 487214 39208 487219 39264
rect 201420 39206 487219 39208
rect 201420 39204 201426 39206
rect 487153 39203 487219 39206
rect 583520 33146 584960 33236
rect 583342 33086 584960 33146
rect 583342 33010 583402 33086
rect 583520 33010 584960 33086
rect 583342 32996 584960 33010
rect 583342 32950 583586 32996
rect -960 32466 480 32556
rect 2865 32466 2931 32469
rect -960 32464 2931 32466
rect -960 32408 2870 32464
rect 2926 32408 2931 32464
rect -960 32406 2931 32408
rect -960 32316 480 32406
rect 2865 32403 2931 32406
rect 183318 32404 183324 32468
rect 183388 32466 183394 32468
rect 269113 32466 269179 32469
rect 183388 32464 269179 32466
rect 183388 32408 269118 32464
rect 269174 32408 269179 32464
rect 183388 32406 269179 32408
rect 183388 32404 183394 32406
rect 269113 32403 269179 32406
rect 331806 31724 331812 31788
rect 331876 31786 331882 31788
rect 583526 31786 583586 32950
rect 331876 31726 583586 31786
rect 331876 31724 331882 31726
rect 177614 28188 177620 28252
rect 177684 28250 177690 28252
rect 193857 28250 193923 28253
rect 177684 28248 193923 28250
rect 177684 28192 193862 28248
rect 193918 28192 193923 28248
rect 177684 28190 193923 28192
rect 177684 28188 177690 28190
rect 193857 28187 193923 28190
rect 183870 26828 183876 26892
rect 183940 26890 183946 26892
rect 287053 26890 287119 26893
rect 183940 26888 287119 26890
rect 183940 26832 287058 26888
rect 287114 26832 287119 26888
rect 183940 26830 287119 26832
rect 183940 26828 183946 26830
rect 287053 26827 287119 26830
rect 194358 21252 194364 21316
rect 194428 21314 194434 21316
rect 397453 21314 397519 21317
rect 194428 21312 397519 21314
rect 194428 21256 397458 21312
rect 397514 21256 397519 21312
rect 194428 21254 397519 21256
rect 194428 21252 194434 21254
rect 397453 21251 397519 21254
rect 580073 19818 580139 19821
rect 583520 19818 584960 19908
rect 580073 19816 584960 19818
rect 580073 19760 580078 19816
rect 580134 19760 584960 19816
rect 580073 19758 584960 19760
rect 580073 19755 580139 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 177798 17172 177804 17236
rect 177868 17234 177874 17236
rect 196617 17234 196683 17237
rect 177868 17232 196683 17234
rect 177868 17176 196622 17232
rect 196678 17176 196683 17232
rect 177868 17174 196683 17176
rect 177868 17172 177874 17174
rect 196617 17171 196683 17174
rect 195646 14452 195652 14516
rect 195716 14514 195722 14516
rect 429193 14514 429259 14517
rect 195716 14512 429259 14514
rect 195716 14456 429198 14512
rect 429254 14456 429259 14512
rect 195716 14454 429259 14456
rect 195716 14452 195722 14454
rect 429193 14451 429259 14454
rect 187550 12956 187556 13020
rect 187620 13018 187626 13020
rect 322933 13018 322999 13021
rect 187620 13016 322999 13018
rect 187620 12960 322938 13016
rect 322994 12960 322999 13016
rect 187620 12958 322999 12960
rect 187620 12956 187626 12958
rect 322933 12955 322999 12958
rect 190126 9420 190132 9484
rect 190196 9482 190202 9484
rect 358721 9482 358787 9485
rect 190196 9480 358787 9482
rect 190196 9424 358726 9480
rect 358782 9424 358787 9480
rect 190196 9422 358787 9424
rect 190196 9420 190202 9422
rect 358721 9419 358787 9422
rect 195462 9284 195468 9348
rect 195532 9346 195538 9348
rect 415485 9346 415551 9349
rect 195532 9344 415551 9346
rect 195532 9288 415490 9344
rect 415546 9288 415551 9344
rect 195532 9286 415551 9288
rect 195532 9284 195538 9286
rect 415485 9283 415551 9286
rect 195094 9148 195100 9212
rect 195164 9210 195170 9212
rect 418981 9210 419047 9213
rect 195164 9208 419047 9210
rect 195164 9152 418986 9208
rect 419042 9152 419047 9208
rect 195164 9150 419047 9152
rect 195164 9148 195170 9150
rect 418981 9147 419047 9150
rect 196566 9012 196572 9076
rect 196636 9074 196642 9076
rect 436829 9074 436895 9077
rect 196636 9072 436895 9074
rect 196636 9016 436834 9072
rect 436890 9016 436895 9072
rect 196636 9014 436895 9016
rect 196636 9012 196642 9014
rect 436829 9011 436895 9014
rect 196934 8876 196940 8940
rect 197004 8938 197010 8940
rect 440325 8938 440391 8941
rect 197004 8936 440391 8938
rect 197004 8880 440330 8936
rect 440386 8880 440391 8936
rect 197004 8878 440391 8880
rect 197004 8876 197010 8878
rect 440325 8875 440391 8878
rect 188470 6836 188476 6900
rect 188540 6898 188546 6900
rect 330385 6898 330451 6901
rect 188540 6896 330451 6898
rect 188540 6840 330390 6896
rect 330446 6840 330451 6896
rect 188540 6838 330451 6840
rect 188540 6836 188546 6838
rect 330385 6835 330451 6838
rect 188838 6700 188844 6764
rect 188908 6762 188914 6764
rect 333881 6762 333947 6765
rect 188908 6760 333947 6762
rect 188908 6704 333886 6760
rect 333942 6704 333947 6760
rect 188908 6702 333947 6704
rect 188908 6700 188914 6702
rect 333881 6699 333947 6702
rect -960 6490 480 6580
rect 188654 6564 188660 6628
rect 188724 6626 188730 6628
rect 337469 6626 337535 6629
rect 188724 6624 337535 6626
rect 188724 6568 337474 6624
rect 337530 6568 337535 6624
rect 188724 6566 337535 6568
rect 188724 6564 188730 6566
rect 337469 6563 337535 6566
rect 580349 6626 580415 6629
rect 583520 6626 584960 6716
rect 580349 6624 584960 6626
rect 580349 6568 580354 6624
rect 580410 6568 584960 6624
rect 580349 6566 584960 6568
rect 580349 6563 580415 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 192702 6428 192708 6492
rect 192772 6490 192778 6492
rect 379973 6490 380039 6493
rect 192772 6488 380039 6490
rect 192772 6432 379978 6488
rect 380034 6432 380039 6488
rect 583520 6476 584960 6566
rect 192772 6430 380039 6432
rect 192772 6428 192778 6430
rect 379973 6427 380039 6430
rect 192518 6292 192524 6356
rect 192588 6354 192594 6356
rect 390645 6354 390711 6357
rect 192588 6352 390711 6354
rect 192588 6296 390650 6352
rect 390706 6296 390711 6352
rect 192588 6294 390711 6296
rect 192588 6292 192594 6294
rect 390645 6291 390711 6294
rect 192886 6156 192892 6220
rect 192956 6218 192962 6220
rect 394233 6218 394299 6221
rect 192956 6216 394299 6218
rect 192956 6160 394238 6216
rect 394294 6160 394299 6216
rect 192956 6158 394299 6160
rect 192956 6156 192962 6158
rect 394233 6155 394299 6158
rect 185158 6020 185164 6084
rect 185228 6082 185234 6084
rect 301957 6082 302023 6085
rect 185228 6080 302023 6082
rect 185228 6024 301962 6080
rect 302018 6024 302023 6080
rect 185228 6022 302023 6024
rect 185228 6020 185234 6022
rect 301957 6019 302023 6022
rect 190310 3708 190316 3772
rect 190380 3770 190386 3772
rect 351637 3770 351703 3773
rect 190380 3768 351703 3770
rect 190380 3712 351642 3768
rect 351698 3712 351703 3768
rect 190380 3710 351703 3712
rect 190380 3708 190386 3710
rect 351637 3707 351703 3710
rect 353334 3708 353340 3772
rect 353404 3770 353410 3772
rect 354029 3770 354095 3773
rect 353404 3768 354095 3770
rect 353404 3712 354034 3768
rect 354090 3712 354095 3768
rect 353404 3710 354095 3712
rect 353404 3708 353410 3710
rect 354029 3707 354095 3710
rect 198590 3572 198596 3636
rect 198660 3634 198666 3636
rect 458081 3634 458147 3637
rect 198660 3632 458147 3634
rect 198660 3576 458086 3632
rect 458142 3576 458147 3632
rect 198660 3574 458147 3576
rect 198660 3572 198666 3574
rect 458081 3571 458147 3574
rect 198406 3436 198412 3500
rect 198476 3498 198482 3500
rect 465165 3498 465231 3501
rect 198476 3496 465231 3498
rect 198476 3440 465170 3496
rect 465226 3440 465231 3496
rect 198476 3438 465231 3440
rect 198476 3436 198482 3438
rect 465165 3435 465231 3438
rect 199878 3300 199884 3364
rect 199948 3362 199954 3364
rect 482829 3362 482895 3365
rect 199948 3360 482895 3362
rect 199948 3304 482834 3360
rect 482890 3304 482895 3360
rect 199948 3302 482895 3304
rect 199948 3300 199954 3302
rect 482829 3299 482895 3302
<< via3 >>
rect 279924 452644 279988 452708
rect 372660 452568 372724 452572
rect 372660 452512 372674 452568
rect 372674 452512 372724 452568
rect 372660 452508 372724 452512
rect 374132 452568 374196 452572
rect 374132 452512 374146 452568
rect 374146 452512 374196 452568
rect 374132 452508 374196 452512
rect 343588 452100 343652 452164
rect 278636 451828 278700 451892
rect 357388 451556 357452 451620
rect 346348 451420 346412 451484
rect 368980 451420 369044 451484
rect 347636 451284 347700 451348
rect 355180 451284 355244 451348
rect 375972 451284 376036 451348
rect 343956 449380 344020 449444
rect 345244 449440 345308 449444
rect 345244 449384 345258 449440
rect 345258 449384 345308 449440
rect 345244 449380 345308 449384
rect 349660 449380 349724 449444
rect 353340 449440 353404 449444
rect 353340 449384 353390 449440
rect 353390 449384 353404 449440
rect 353340 449380 353404 449384
rect 344876 449244 344940 449308
rect 357572 449380 357636 449444
rect 370452 449380 370516 449444
rect 371556 449380 371620 449444
rect 372660 449380 372724 449444
rect 374132 449380 374196 449444
rect 382228 449380 382292 449444
rect 383884 449440 383948 449444
rect 383884 449384 383898 449440
rect 383898 449384 383948 449440
rect 383884 449380 383948 449384
rect 384252 449440 384316 449444
rect 384252 449384 384302 449440
rect 384302 449384 384316 449440
rect 384252 449380 384316 449384
rect 385356 449380 385420 449444
rect 373948 449244 374012 449308
rect 382964 449244 383028 449308
rect 346348 447748 346412 447812
rect 343588 446388 343652 446452
rect 343956 444892 344020 444956
rect 345244 401916 345308 401980
rect 352788 401780 352852 401844
rect 368980 401236 369044 401300
rect 375972 401100 376036 401164
rect 357572 400964 357636 401028
rect 347636 400828 347700 400892
rect 353524 400692 353588 400756
rect 343220 400556 343284 400620
rect 348556 400556 348620 400620
rect 354260 400556 354324 400620
rect 385724 400420 385788 400484
rect 381308 400284 381372 400348
rect 355180 400148 355244 400212
rect 344876 400012 344940 400076
rect 348556 400012 348620 400076
rect 351316 400012 351380 400076
rect 357388 400012 357452 400076
rect 346532 399876 346596 399940
rect 346900 399876 346964 399940
rect 347084 399936 347148 399940
rect 347084 399880 347088 399936
rect 347088 399880 347144 399936
rect 347144 399880 347148 399936
rect 347084 399876 347148 399880
rect 347820 399936 347884 399940
rect 347820 399880 347824 399936
rect 347824 399880 347880 399936
rect 347880 399880 347884 399936
rect 347820 399876 347884 399880
rect 348188 399876 348252 399940
rect 348740 399876 348804 399940
rect 349844 399876 349908 399940
rect 350212 399876 350276 399940
rect 351132 399876 351196 399940
rect 352420 399876 352484 399940
rect 353524 399876 353588 399940
rect 354306 399936 354370 399940
rect 354306 399880 354356 399936
rect 354356 399880 354370 399936
rect 354306 399876 354370 399880
rect 354812 399936 354876 399940
rect 354812 399880 354816 399936
rect 354816 399880 354872 399936
rect 354872 399880 354876 399936
rect 354812 399876 354876 399880
rect 354996 399876 355060 399940
rect 356468 399876 356532 399940
rect 356836 399876 356900 399940
rect 357572 399876 357636 399940
rect 358124 399876 358188 399940
rect 358676 399876 358740 399940
rect 359044 399876 359108 399940
rect 346348 399740 346412 399804
rect 346716 399800 346780 399804
rect 346716 399744 346766 399800
rect 346766 399744 346780 399800
rect 346716 399740 346780 399744
rect 347268 399740 347332 399804
rect 359780 399876 359844 399940
rect 360332 399876 360396 399940
rect 361068 399876 361132 399940
rect 363276 399936 363340 399940
rect 363276 399880 363280 399936
rect 363280 399880 363336 399936
rect 363336 399880 363340 399936
rect 363276 399876 363340 399880
rect 363828 399876 363892 399940
rect 359412 399740 359476 399804
rect 360516 399740 360580 399804
rect 361252 399740 361316 399804
rect 362908 399740 362972 399804
rect 364380 399876 364444 399940
rect 364932 399876 364996 399940
rect 368428 400012 368492 400076
rect 368060 399876 368124 399940
rect 369164 399936 369228 399940
rect 369164 399880 369168 399936
rect 369168 399880 369224 399936
rect 369224 399880 369228 399936
rect 369164 399876 369228 399880
rect 369532 399936 369596 399940
rect 369532 399880 369536 399936
rect 369536 399880 369592 399936
rect 369592 399880 369596 399936
rect 369532 399876 369596 399880
rect 370084 399876 370148 399940
rect 370636 399936 370700 399940
rect 370636 399880 370640 399936
rect 370640 399880 370696 399936
rect 370696 399880 370700 399936
rect 370636 399876 370700 399880
rect 364932 399740 364996 399804
rect 365300 399740 365364 399804
rect 366404 399740 366468 399804
rect 368244 399740 368308 399804
rect 368612 399740 368676 399804
rect 374132 400012 374196 400076
rect 346348 399468 346412 399532
rect 352788 399468 352852 399532
rect 353340 399468 353404 399532
rect 359044 399468 359108 399532
rect 360700 399468 360764 399532
rect 366588 399468 366652 399532
rect 370452 399528 370516 399532
rect 370452 399472 370502 399528
rect 370502 399472 370516 399528
rect 370452 399468 370516 399472
rect 348924 399332 348988 399396
rect 343220 399196 343284 399260
rect 354812 399196 354876 399260
rect 358860 399196 358924 399260
rect 287652 398924 287716 398988
rect 375052 399936 375116 399940
rect 375052 399880 375056 399936
rect 375056 399880 375112 399936
rect 375112 399880 375116 399936
rect 372844 399332 372908 399396
rect 375052 399876 375116 399880
rect 375788 399936 375852 399940
rect 375788 399880 375792 399936
rect 375792 399880 375848 399936
rect 375848 399880 375852 399936
rect 375788 399876 375852 399880
rect 376524 400012 376588 400076
rect 377260 400012 377324 400076
rect 376708 399936 376772 399940
rect 376708 399880 376712 399936
rect 376712 399880 376768 399936
rect 376768 399880 376772 399936
rect 376708 399876 376772 399880
rect 378732 399936 378796 399940
rect 378732 399880 378736 399936
rect 378736 399880 378792 399936
rect 378792 399880 378796 399936
rect 378732 399876 378796 399880
rect 380204 399876 380268 399940
rect 353892 398924 353956 398988
rect 372660 399060 372724 399124
rect 376892 399332 376956 399396
rect 378916 399740 378980 399804
rect 381078 399936 381142 399940
rect 381078 399880 381092 399936
rect 381092 399880 381142 399936
rect 381078 399876 381142 399880
rect 378180 399196 378244 399260
rect 379652 399196 379716 399260
rect 384988 400012 385052 400076
rect 381492 399876 381556 399940
rect 382228 399740 382292 399804
rect 381308 399664 381372 399668
rect 381308 399608 381322 399664
rect 381322 399608 381372 399664
rect 381308 399604 381372 399608
rect 381676 399604 381740 399668
rect 359044 398924 359108 398988
rect 360332 398924 360396 398988
rect 384436 399196 384500 399260
rect 385724 399604 385788 399668
rect 293172 398788 293236 398852
rect 346348 398788 346412 398852
rect 348924 398788 348988 398852
rect 360332 398788 360396 398852
rect 374500 398848 374564 398852
rect 374500 398792 374514 398848
rect 374514 398792 374564 398848
rect 374500 398788 374564 398792
rect 366588 398712 366652 398716
rect 366588 398656 366602 398712
rect 366602 398656 366652 398712
rect 366588 398652 366652 398656
rect 370084 398712 370148 398716
rect 370084 398656 370098 398712
rect 370098 398656 370148 398712
rect 370084 398652 370148 398656
rect 380756 398652 380820 398716
rect 381492 398652 381556 398716
rect 346532 398516 346596 398580
rect 351316 398516 351380 398580
rect 364748 398516 364812 398580
rect 370084 398516 370148 398580
rect 349292 398380 349356 398444
rect 352052 398380 352116 398444
rect 370636 398440 370700 398444
rect 370636 398384 370650 398440
rect 370650 398384 370700 398440
rect 356836 398244 356900 398308
rect 356836 398108 356900 398172
rect 345244 397972 345308 398036
rect 350764 397972 350828 398036
rect 355364 397972 355428 398036
rect 350580 397836 350644 397900
rect 362724 397972 362788 398036
rect 363460 398108 363524 398172
rect 370636 398380 370700 398384
rect 376708 398380 376772 398444
rect 383700 398380 383764 398444
rect 372660 398244 372724 398308
rect 367324 398108 367388 398172
rect 367692 398108 367756 398172
rect 368244 398032 368308 398036
rect 368244 397976 368294 398032
rect 368294 397976 368308 398032
rect 368244 397972 368308 397976
rect 368980 397972 369044 398036
rect 365300 397836 365364 397900
rect 369532 397836 369596 397900
rect 369900 397836 369964 397900
rect 372844 397836 372908 397900
rect 382780 397836 382844 397900
rect 348004 397564 348068 397628
rect 370268 397700 370332 397764
rect 369164 397564 369228 397628
rect 382228 397564 382292 397628
rect 351868 397428 351932 397492
rect 353340 397488 353404 397492
rect 353340 397432 353354 397488
rect 353354 397432 353404 397488
rect 353340 397428 353404 397432
rect 357388 397428 357452 397492
rect 371372 397428 371436 397492
rect 373212 397428 373276 397492
rect 378364 397428 378428 397492
rect 380940 397428 381004 397492
rect 363644 397292 363708 397356
rect 366588 397352 366652 397356
rect 366588 397296 366638 397352
rect 366638 397296 366652 397352
rect 366588 397292 366652 397296
rect 367140 397352 367204 397356
rect 367140 397296 367190 397352
rect 367190 397296 367204 397352
rect 367140 397292 367204 397296
rect 356652 397156 356716 397220
rect 364748 397156 364812 397220
rect 318564 397020 318628 397084
rect 315804 396884 315868 396948
rect 375788 396884 375852 396948
rect 380204 396884 380268 396948
rect 350212 396748 350276 396812
rect 350948 396748 351012 396812
rect 357940 396748 358004 396812
rect 361068 396748 361132 396812
rect 354996 396672 355060 396676
rect 354996 396616 355010 396672
rect 355010 396616 355060 396672
rect 354996 396612 355060 396616
rect 373948 396612 374012 396676
rect 359412 396476 359476 396540
rect 345060 396128 345124 396132
rect 345060 396072 345074 396128
rect 345074 396072 345124 396128
rect 345060 396068 345124 396072
rect 357020 396068 357084 396132
rect 368060 396068 368124 396132
rect 385172 396068 385236 396132
rect 283420 395932 283484 395996
rect 313044 395932 313108 395996
rect 343588 395796 343652 395860
rect 363276 395660 363340 395724
rect 355180 395524 355244 395588
rect 347084 395388 347148 395452
rect 347820 395388 347884 395452
rect 349844 395388 349908 395452
rect 359412 395388 359476 395452
rect 364380 395388 364444 395452
rect 358124 395252 358188 395316
rect 364380 395252 364444 395316
rect 375052 395252 375116 395316
rect 378732 395252 378796 395316
rect 378916 395252 378980 395316
rect 283604 395116 283668 395180
rect 346716 394980 346780 395044
rect 349108 394980 349172 395044
rect 359780 394980 359844 395044
rect 364932 394980 364996 395044
rect 348740 394844 348804 394908
rect 295564 394436 295628 394500
rect 363828 394436 363892 394500
rect 286916 394300 286980 394364
rect 296116 394164 296180 394228
rect 352052 394028 352116 394092
rect 358676 393892 358740 393956
rect 371372 393892 371436 393956
rect 297956 393756 298020 393820
rect 296484 393620 296548 393684
rect 351132 393484 351196 393548
rect 381124 393484 381188 393548
rect 302188 393076 302252 393140
rect 302004 392940 302068 393004
rect 361252 392940 361316 393004
rect 297036 392804 297100 392868
rect 357572 392804 357636 392868
rect 368612 392668 368676 392732
rect 360516 392532 360580 392596
rect 298508 392396 298572 392460
rect 292988 392260 293052 392324
rect 374500 392124 374564 392188
rect 285076 391852 285140 391916
rect 310284 391852 310348 391916
rect 295196 391716 295260 391780
rect 295012 391580 295076 391644
rect 292804 391444 292868 391508
rect 349292 391308 349356 391372
rect 375420 391308 375484 391372
rect 288940 391036 289004 391100
rect 307708 390628 307772 390692
rect 317276 390492 317340 390556
rect 320036 390356 320100 390420
rect 294644 390220 294708 390284
rect 357020 390220 357084 390284
rect 317092 390084 317156 390148
rect 346716 389812 346780 389876
rect 294828 389676 294892 389740
rect 348188 389132 348252 389196
rect 344140 388996 344204 389060
rect 383884 388996 383948 389060
rect 286364 388860 286428 388924
rect 288204 388724 288268 388788
rect 289492 388588 289556 388652
rect 345244 388452 345308 388516
rect 385356 388452 385420 388516
rect 348004 388316 348068 388380
rect 363644 388180 363708 388244
rect 371556 387636 371620 387700
rect 356468 387500 356532 387564
rect 283788 387364 283852 387428
rect 297588 387228 297652 387292
rect 359044 387092 359108 387156
rect 285444 386956 285508 387020
rect 343036 386820 343100 386884
rect 349660 386820 349724 386884
rect 342852 386684 342916 386748
rect 368980 386004 369044 386068
rect 330524 385868 330588 385932
rect 286548 385732 286612 385796
rect 382964 385732 383028 385796
rect 353340 385596 353404 385660
rect 295932 384372 295996 384436
rect 370268 384236 370332 384300
rect 355364 383420 355428 383484
rect 364564 383284 364628 383348
rect 304948 383148 305012 383212
rect 351868 383012 351932 383076
rect 356836 382876 356900 382940
rect 285260 381788 285324 381852
rect 290964 381652 291028 381716
rect 299980 381516 300044 381580
rect 297404 380156 297468 380220
rect 290780 379340 290844 379404
rect 291884 379204 291948 379268
rect 292252 379068 292316 379132
rect 306972 378932 307036 378996
rect 366588 378932 366652 378996
rect 289308 378796 289372 378860
rect 289124 378660 289188 378724
rect 314332 377708 314396 377772
rect 283972 377572 284036 377636
rect 343588 377572 343652 377636
rect 372660 377572 372724 377636
rect 308996 377436 309060 377500
rect 292068 377300 292132 377364
rect 277900 375396 277964 375460
rect 306236 373492 306300 373556
rect 291700 373356 291764 373420
rect 307524 373220 307588 373284
rect 367324 373220 367388 373284
rect 278452 372948 278516 373012
rect 221228 372676 221292 372740
rect 324268 372268 324332 372332
rect 282316 371920 282380 371924
rect 282316 371864 282330 371920
rect 282330 371864 282380 371920
rect 282316 371860 282380 371864
rect 344140 371860 344204 371924
rect 281028 371724 281092 371788
rect 279372 371588 279436 371652
rect 280844 371588 280908 371652
rect 276612 371452 276676 371516
rect 323164 371452 323228 371516
rect 343036 370636 343100 370700
rect 315620 370500 315684 370564
rect 280660 370228 280724 370292
rect 333100 370092 333164 370156
rect 331812 369956 331876 370020
rect 282132 369820 282196 369884
rect 285628 369548 285692 369612
rect 287284 369608 287348 369612
rect 287284 369552 287288 369608
rect 287288 369552 287344 369608
rect 287344 369552 287348 369608
rect 287284 369548 287348 369552
rect 279924 369276 279988 369340
rect 287284 369336 287348 369340
rect 287284 369280 287288 369336
rect 287288 369280 287344 369336
rect 287344 369280 287348 369336
rect 278636 369140 278700 369204
rect 281396 369140 281460 369204
rect 287284 369276 287348 369280
rect 315436 369684 315500 369748
rect 311020 369548 311084 369612
rect 313780 369548 313844 369612
rect 319300 369548 319364 369612
rect 320956 369548 321020 369612
rect 301452 369412 301516 369476
rect 302740 369412 302804 369476
rect 311204 369412 311268 369476
rect 312492 369412 312556 369476
rect 313596 369412 313660 369476
rect 318012 369412 318076 369476
rect 319668 369412 319732 369476
rect 321140 369412 321204 369476
rect 310100 369336 310164 369340
rect 310100 369280 310104 369336
rect 310104 369280 310160 369336
rect 310160 369280 310164 369336
rect 310100 369276 310164 369280
rect 285628 368732 285692 368796
rect 287284 368596 287348 368660
rect 310100 368324 310164 368388
rect 324268 366284 324332 366348
rect 323164 364924 323228 364988
rect 281028 363564 281092 363628
rect 280844 362204 280908 362268
rect 278452 358804 278516 358868
rect 282316 357988 282380 358052
rect 350948 357988 351012 358052
rect 323716 356628 323780 356692
rect 323900 342892 323964 342956
rect 325372 341396 325436 341460
rect 324636 340036 324700 340100
rect 376524 338132 376588 338196
rect 380756 335412 380820 335476
rect 380756 334596 380820 334660
rect 329236 330516 329300 330580
rect 325372 327116 325436 327180
rect 338620 326300 338684 326364
rect 370084 325212 370148 325276
rect 378364 325076 378428 325140
rect 323532 324396 323596 324460
rect 382228 324940 382292 325004
rect 276612 323580 276676 323644
rect 324084 323580 324148 323644
rect 327764 322900 327828 322964
rect 326660 322220 326724 322284
rect 330340 322220 330404 322284
rect 385172 322220 385236 322284
rect 324452 322084 324516 322148
rect 320772 321948 320836 322012
rect 308812 321812 308876 321876
rect 283972 321540 284036 321604
rect 327396 321600 327460 321604
rect 327396 321544 327446 321600
rect 327446 321544 327460 321600
rect 327396 321540 327460 321544
rect 320588 321404 320652 321468
rect 294460 321268 294524 321332
rect 320956 321268 321020 321332
rect 321508 321268 321572 321332
rect 322980 321268 323044 321332
rect 279372 321132 279436 321196
rect 294276 321132 294340 321196
rect 295196 321132 295260 321196
rect 301452 321132 301516 321196
rect 306972 321132 307036 321196
rect 318932 321132 318996 321196
rect 303292 320996 303356 321060
rect 321324 320996 321388 321060
rect 378180 320996 378244 321060
rect 283788 320724 283852 320788
rect 283972 320724 284036 320788
rect 287100 320860 287164 320924
rect 288204 320784 288268 320788
rect 288204 320728 288208 320784
rect 288208 320728 288264 320784
rect 288264 320728 288268 320784
rect 288204 320724 288268 320728
rect 290964 320724 291028 320788
rect 291700 320724 291764 320788
rect 292068 320724 292132 320788
rect 292436 320724 292500 320788
rect 295932 320724 295996 320788
rect 283604 320648 283668 320652
rect 283604 320592 283608 320648
rect 283608 320592 283664 320648
rect 283664 320592 283668 320648
rect 283604 320588 283668 320592
rect 283972 320588 284036 320652
rect 286364 320588 286428 320652
rect 283420 320452 283484 320516
rect 283972 320316 284036 320380
rect 284340 320376 284404 320380
rect 285260 320452 285324 320516
rect 285812 320452 285876 320516
rect 286916 320452 286980 320516
rect 288388 320452 288452 320516
rect 292068 320452 292132 320516
rect 292804 320452 292868 320516
rect 293356 320452 293420 320516
rect 294276 320452 294340 320516
rect 294644 320452 294708 320516
rect 295564 320588 295628 320652
rect 296300 320724 296364 320788
rect 296668 320724 296732 320788
rect 297956 320724 298020 320788
rect 298508 320724 298572 320788
rect 299060 320784 299124 320788
rect 299060 320728 299064 320784
rect 299064 320728 299120 320784
rect 299120 320728 299124 320784
rect 299060 320724 299124 320728
rect 302556 320724 302620 320788
rect 306972 320724 307036 320788
rect 308812 320784 308876 320788
rect 308812 320728 308816 320784
rect 308816 320728 308872 320784
rect 308872 320728 308876 320784
rect 308812 320724 308876 320728
rect 323532 320784 323596 320788
rect 323532 320728 323536 320784
rect 323536 320728 323592 320784
rect 323592 320728 323596 320784
rect 312676 320588 312740 320652
rect 314884 320588 314948 320652
rect 315804 320648 315868 320652
rect 315804 320592 315808 320648
rect 315808 320592 315864 320648
rect 315864 320592 315868 320648
rect 315804 320588 315868 320592
rect 316908 320588 316972 320652
rect 317460 320588 317524 320652
rect 318012 320648 318076 320652
rect 318012 320592 318016 320648
rect 318016 320592 318072 320648
rect 318072 320592 318076 320648
rect 318012 320588 318076 320592
rect 318196 320648 318260 320652
rect 318196 320592 318200 320648
rect 318200 320592 318256 320648
rect 318256 320592 318260 320648
rect 318196 320588 318260 320592
rect 318932 320648 318996 320652
rect 318932 320592 318936 320648
rect 318936 320592 318992 320648
rect 318992 320592 318996 320648
rect 318932 320588 318996 320592
rect 321324 320588 321388 320652
rect 296852 320452 296916 320516
rect 298324 320452 298388 320516
rect 298876 320452 298940 320516
rect 302188 320452 302252 320516
rect 305316 320452 305380 320516
rect 306052 320452 306116 320516
rect 307708 320452 307772 320516
rect 310836 320452 310900 320516
rect 322980 320588 323044 320652
rect 323532 320724 323596 320728
rect 324084 320784 324148 320788
rect 324084 320728 324088 320784
rect 324088 320728 324144 320784
rect 324144 320728 324148 320784
rect 324084 320724 324148 320728
rect 324820 320724 324884 320788
rect 325372 320724 325436 320788
rect 326660 320724 326724 320788
rect 322060 320512 322124 320516
rect 322060 320456 322064 320512
rect 322064 320456 322120 320512
rect 322120 320456 322124 320512
rect 284340 320320 284344 320376
rect 284344 320320 284400 320376
rect 284400 320320 284404 320376
rect 284340 320316 284404 320320
rect 285076 320316 285140 320380
rect 286548 320316 286612 320380
rect 287468 320316 287532 320380
rect 288388 320316 288452 320380
rect 289492 320376 289556 320380
rect 289492 320320 289496 320376
rect 289496 320320 289552 320376
rect 289552 320320 289556 320376
rect 289492 320316 289556 320320
rect 290780 320316 290844 320380
rect 292252 320316 292316 320380
rect 292620 320316 292684 320380
rect 294460 320316 294524 320380
rect 309548 320376 309612 320380
rect 309548 320320 309552 320376
rect 309552 320320 309608 320376
rect 309608 320320 309612 320376
rect 309548 320316 309612 320320
rect 309916 320316 309980 320380
rect 310284 320376 310348 320380
rect 310284 320320 310288 320376
rect 310288 320320 310344 320376
rect 310344 320320 310348 320376
rect 310284 320316 310348 320320
rect 310652 320376 310716 320380
rect 310652 320320 310656 320376
rect 310656 320320 310712 320376
rect 310712 320320 310716 320376
rect 310652 320316 310716 320320
rect 311020 320316 311084 320380
rect 311388 320376 311452 320380
rect 311388 320320 311392 320376
rect 311392 320320 311448 320376
rect 311448 320320 311452 320376
rect 311388 320316 311452 320320
rect 292804 320240 292868 320244
rect 292804 320184 292808 320240
rect 292808 320184 292864 320240
rect 292864 320184 292868 320240
rect 283972 320044 284036 320108
rect 284892 320044 284956 320108
rect 285444 320044 285508 320108
rect 285628 320044 285692 320108
rect 287100 320104 287164 320108
rect 287100 320048 287104 320104
rect 287104 320048 287160 320104
rect 287160 320048 287164 320104
rect 287100 320044 287164 320048
rect 286364 319636 286428 319700
rect 288756 320044 288820 320108
rect 289124 320044 289188 320108
rect 290596 320044 290660 320108
rect 291884 320044 291948 320108
rect 292804 320180 292868 320184
rect 292988 320180 293052 320244
rect 294828 320180 294892 320244
rect 295748 320180 295812 320244
rect 296484 320180 296548 320244
rect 297036 320240 297100 320244
rect 297036 320184 297040 320240
rect 297040 320184 297096 320240
rect 297096 320184 297100 320240
rect 297036 320180 297100 320184
rect 293172 320044 293236 320108
rect 291148 319696 291212 319700
rect 291148 319640 291162 319696
rect 291162 319640 291212 319696
rect 291148 319636 291212 319640
rect 294460 320104 294524 320108
rect 294460 320048 294464 320104
rect 294464 320048 294520 320104
rect 294520 320048 294524 320104
rect 294460 320044 294524 320048
rect 295196 320044 295260 320108
rect 295012 319908 295076 319972
rect 297588 320104 297652 320108
rect 297588 320048 297592 320104
rect 297592 320048 297648 320104
rect 297648 320048 297652 320104
rect 297588 320044 297652 320048
rect 296116 319832 296180 319836
rect 296116 319776 296166 319832
rect 296166 319776 296180 319832
rect 296116 319772 296180 319776
rect 292804 319500 292868 319564
rect 297588 319772 297652 319836
rect 299428 320180 299492 320244
rect 300900 320180 300964 320244
rect 302004 320240 302068 320244
rect 302004 320184 302008 320240
rect 302008 320184 302064 320240
rect 302064 320184 302068 320240
rect 302004 320180 302068 320184
rect 302188 320180 302252 320244
rect 307708 320180 307772 320244
rect 322060 320452 322124 320456
rect 322612 320452 322676 320516
rect 323348 320512 323412 320516
rect 323348 320456 323352 320512
rect 323352 320456 323408 320512
rect 323408 320456 323412 320512
rect 323348 320452 323412 320456
rect 323532 320452 323596 320516
rect 325004 320452 325068 320516
rect 299244 320104 299308 320108
rect 299244 320048 299248 320104
rect 299248 320048 299304 320104
rect 299304 320048 299308 320104
rect 299244 320044 299308 320048
rect 299796 320044 299860 320108
rect 301268 320044 301332 320108
rect 302372 320044 302436 320108
rect 297956 319908 298020 319972
rect 298508 319636 298572 319700
rect 299060 319636 299124 319700
rect 301636 319908 301700 319972
rect 303292 319696 303356 319700
rect 305500 320044 305564 320108
rect 305684 319908 305748 319972
rect 307524 320104 307588 320108
rect 307524 320048 307528 320104
rect 307528 320048 307584 320104
rect 307584 320048 307588 320104
rect 307524 320044 307588 320048
rect 307708 320044 307772 320108
rect 308996 320044 309060 320108
rect 303292 319640 303342 319696
rect 303342 319640 303356 319696
rect 303292 319636 303356 319640
rect 283604 319364 283668 319428
rect 302372 319364 302436 319428
rect 311204 320044 311268 320108
rect 311940 320104 312004 320108
rect 311940 320048 311944 320104
rect 311944 320048 312000 320104
rect 312000 320048 312004 320104
rect 311940 320044 312004 320048
rect 312492 320044 312556 320108
rect 313044 320044 313108 320108
rect 313964 320180 314028 320244
rect 314332 320180 314396 320244
rect 313596 320044 313660 320108
rect 314148 320044 314212 320108
rect 309548 319636 309612 319700
rect 315068 320044 315132 320108
rect 315620 320044 315684 320108
rect 318564 320180 318628 320244
rect 319300 320316 319364 320380
rect 320588 320316 320652 320380
rect 321324 320316 321388 320380
rect 322428 320316 322492 320380
rect 323900 320316 323964 320380
rect 324268 320376 324332 320380
rect 324268 320320 324272 320376
rect 324272 320320 324328 320376
rect 324328 320320 324332 320376
rect 324268 320316 324332 320320
rect 324452 320316 324516 320380
rect 326660 320316 326724 320380
rect 327396 320376 327460 320380
rect 327396 320320 327400 320376
rect 327400 320320 327456 320376
rect 327456 320320 327460 320376
rect 327396 320316 327460 320320
rect 327764 320316 327828 320380
rect 316724 320044 316788 320108
rect 317276 320044 317340 320108
rect 317644 320044 317708 320108
rect 319116 320104 319180 320108
rect 319116 320048 319120 320104
rect 319120 320048 319176 320104
rect 319176 320048 319180 320104
rect 313964 319636 314028 319700
rect 315436 319636 315500 319700
rect 319116 320044 319180 320048
rect 319484 320044 319548 320108
rect 320036 320044 320100 320108
rect 320404 320044 320468 320108
rect 321508 320044 321572 320108
rect 324636 320044 324700 320108
rect 326844 320104 326908 320108
rect 326844 320048 326848 320104
rect 326848 320048 326904 320104
rect 326904 320048 326908 320104
rect 326844 320044 326908 320048
rect 309916 319500 309980 319564
rect 310652 319560 310716 319564
rect 310652 319504 310702 319560
rect 310702 319504 310716 319560
rect 310652 319500 310716 319504
rect 317460 319500 317524 319564
rect 352420 319772 352484 319836
rect 322428 319636 322492 319700
rect 323900 319636 323964 319700
rect 324084 319696 324148 319700
rect 324084 319640 324098 319696
rect 324098 319640 324148 319696
rect 324084 319636 324148 319640
rect 324820 319636 324884 319700
rect 330524 319636 330588 319700
rect 362724 319636 362788 319700
rect 322060 319500 322124 319564
rect 326844 319560 326908 319564
rect 326844 319504 326858 319560
rect 326858 319504 326908 319560
rect 326844 319500 326908 319504
rect 367140 319500 367204 319564
rect 318196 319424 318260 319428
rect 318196 319368 318246 319424
rect 318246 319368 318260 319424
rect 318196 319364 318260 319368
rect 319300 319364 319364 319428
rect 320404 319424 320468 319428
rect 320404 319368 320454 319424
rect 320454 319368 320468 319424
rect 320404 319364 320468 319368
rect 321324 319364 321388 319428
rect 287468 319228 287532 319292
rect 288572 319288 288636 319292
rect 288572 319232 288622 319288
rect 288622 319232 288636 319288
rect 288572 319228 288636 319232
rect 292436 319228 292500 319292
rect 298324 319288 298388 319292
rect 298324 319232 298374 319288
rect 298374 319232 298388 319288
rect 298324 319228 298388 319232
rect 298692 319228 298756 319292
rect 310836 319228 310900 319292
rect 288756 319152 288820 319156
rect 288756 319096 288770 319152
rect 288770 319096 288820 319152
rect 288756 319092 288820 319096
rect 291700 319092 291764 319156
rect 318012 318956 318076 319020
rect 321140 318956 321204 319020
rect 322612 318956 322676 319020
rect 323348 318956 323412 319020
rect 324268 319016 324332 319020
rect 324268 318960 324282 319016
rect 324282 318960 324332 319016
rect 324268 318956 324332 318960
rect 325004 319016 325068 319020
rect 325004 318960 325054 319016
rect 325054 318960 325068 319016
rect 325004 318956 325068 318960
rect 326660 319016 326724 319020
rect 326660 318960 326710 319016
rect 326710 318960 326724 319016
rect 326660 318956 326724 318960
rect 327396 319016 327460 319020
rect 327396 318960 327446 319016
rect 327446 318960 327460 319016
rect 327396 318956 327460 318960
rect 283972 318820 284036 318884
rect 290596 318820 290660 318884
rect 291148 318820 291212 318884
rect 304212 318820 304276 318884
rect 305500 318820 305564 318884
rect 283788 318684 283852 318748
rect 287652 318684 287716 318748
rect 302372 318684 302436 318748
rect 316356 318684 316420 318748
rect 317092 318744 317156 318748
rect 317092 318688 317142 318744
rect 317142 318688 317156 318744
rect 317092 318684 317156 318688
rect 319668 318684 319732 318748
rect 283420 318548 283484 318612
rect 288940 318548 289004 318612
rect 302556 318548 302620 318612
rect 309364 318548 309428 318612
rect 310100 318548 310164 318612
rect 328500 318548 328564 318612
rect 284340 318412 284404 318476
rect 294460 318412 294524 318476
rect 316908 318472 316972 318476
rect 316908 318416 316922 318472
rect 316922 318416 316972 318472
rect 316908 318412 316972 318416
rect 323348 318412 323412 318476
rect 247540 318276 247604 318340
rect 285444 318276 285508 318340
rect 289308 318276 289372 318340
rect 306420 318276 306484 318340
rect 292068 318200 292132 318204
rect 292068 318144 292082 318200
rect 292082 318144 292132 318200
rect 292068 318140 292132 318144
rect 237972 318004 238036 318068
rect 291332 318004 291396 318068
rect 299428 318004 299492 318068
rect 303476 318004 303540 318068
rect 318748 318004 318812 318068
rect 369900 318004 369964 318068
rect 283236 317732 283300 317796
rect 291148 317732 291212 317796
rect 298140 317928 298204 317932
rect 298140 317872 298190 317928
rect 298190 317872 298204 317928
rect 298140 317868 298204 317872
rect 299612 317868 299676 317932
rect 302740 317868 302804 317932
rect 304580 317868 304644 317932
rect 306972 317868 307036 317932
rect 311756 317868 311820 317932
rect 313780 317928 313844 317932
rect 313780 317872 313830 317928
rect 313830 317872 313844 317928
rect 313780 317868 313844 317872
rect 320772 317868 320836 317932
rect 320220 317732 320284 317796
rect 323164 317928 323228 317932
rect 323164 317872 323214 317928
rect 323214 317872 323228 317928
rect 323164 317868 323228 317872
rect 329052 317868 329116 317932
rect 326660 317732 326724 317796
rect 328316 317732 328380 317796
rect 317276 317596 317340 317660
rect 327028 317596 327092 317660
rect 283052 317460 283116 317524
rect 295932 317460 295996 317524
rect 299428 317460 299492 317524
rect 301084 317460 301148 317524
rect 302924 317460 302988 317524
rect 304396 317520 304460 317524
rect 304396 317464 304446 317520
rect 304446 317464 304460 317520
rect 304396 317460 304460 317464
rect 307524 317460 307588 317524
rect 312676 317460 312740 317524
rect 315620 317460 315684 317524
rect 316540 317460 316604 317524
rect 318380 317520 318444 317524
rect 318380 317464 318430 317520
rect 318430 317464 318444 317520
rect 318380 317460 318444 317464
rect 321324 317460 321388 317524
rect 321692 317460 321756 317524
rect 223436 316916 223500 316980
rect 306972 316916 307036 316980
rect 366404 316916 366468 316980
rect 231716 316780 231780 316844
rect 297956 316644 298020 316708
rect 319116 316644 319180 316708
rect 326660 316372 326724 316436
rect 338620 316508 338684 316572
rect 328868 316236 328932 316300
rect 328684 316100 328748 316164
rect 295196 315964 295260 316028
rect 237236 315828 237300 315892
rect 296484 315828 296548 315892
rect 360148 315828 360212 315892
rect 235212 315692 235276 315756
rect 291332 315692 291396 315756
rect 296852 315692 296916 315756
rect 301636 315692 301700 315756
rect 224724 315556 224788 315620
rect 237052 315556 237116 315620
rect 297036 315556 297100 315620
rect 314148 315556 314212 315620
rect 382780 315556 382844 315620
rect 296116 315420 296180 315484
rect 295932 315284 295996 315348
rect 316724 315284 316788 315348
rect 299244 315012 299308 315076
rect 295748 314876 295812 314940
rect 307524 314664 307588 314668
rect 307524 314608 307574 314664
rect 307574 314608 307588 314664
rect 307524 314604 307588 314608
rect 232268 314468 232332 314532
rect 318748 314468 318812 314532
rect 241100 314332 241164 314396
rect 223988 314196 224052 314260
rect 298876 314196 298940 314260
rect 223252 314060 223316 314124
rect 244596 314060 244660 314124
rect 305316 314060 305380 314124
rect 232820 313924 232884 313988
rect 292988 313924 293052 313988
rect 239444 313788 239508 313852
rect 299428 313788 299492 313852
rect 241284 313652 241348 313716
rect 299612 313516 299676 313580
rect 301452 313516 301516 313580
rect 247908 313108 247972 313172
rect 249564 312972 249628 313036
rect 309364 312972 309428 313036
rect 252324 312836 252388 312900
rect 226196 312700 226260 312764
rect 251772 312700 251836 312764
rect 234292 312564 234356 312628
rect 292620 312564 292684 312628
rect 299796 312624 299860 312628
rect 299796 312568 299846 312624
rect 299846 312568 299860 312624
rect 299796 312564 299860 312568
rect 311940 312564 312004 312628
rect 327028 312564 327092 312628
rect 311388 312428 311452 312492
rect 234476 312292 234540 312356
rect 293356 312292 293420 312356
rect 310284 312156 310348 312220
rect 282868 311884 282932 311948
rect 283236 311884 283300 311948
rect 232636 311612 232700 311676
rect 291148 311612 291212 311676
rect 318380 311612 318444 311676
rect 318748 311612 318812 311676
rect 230060 311476 230124 311540
rect 231348 311340 231412 311404
rect 291884 311340 291948 311404
rect 231164 311204 231228 311268
rect 292252 311204 292316 311268
rect 380940 311340 381004 311404
rect 229324 311068 229388 311132
rect 290780 311068 290844 311132
rect 287652 310932 287716 310996
rect 318748 310796 318812 310860
rect 228956 310252 229020 310316
rect 298692 310388 298756 310452
rect 227484 310116 227548 310180
rect 228220 309980 228284 310044
rect 288204 309980 288268 310044
rect 244780 309844 244844 309908
rect 308260 309844 308324 309908
rect 315620 309844 315684 309908
rect 375972 309844 376036 309908
rect 225460 309708 225524 309772
rect 286364 309708 286428 309772
rect 312676 308756 312740 308820
rect 303476 308620 303540 308684
rect 355180 308620 355244 308684
rect 238524 308484 238588 308548
rect 342852 308484 342916 308548
rect 234108 308348 234172 308412
rect 294828 308348 294892 308412
rect 299980 308348 300044 308412
rect 236868 307668 236932 307732
rect 296484 307668 296548 307732
rect 283052 307532 283116 307596
rect 384988 307532 385052 307596
rect 289124 307396 289188 307460
rect 297588 307260 297652 307324
rect 357940 307396 358004 307460
rect 356652 307260 356716 307324
rect 301268 306988 301332 307052
rect 222700 306852 222764 306916
rect 329052 306852 329116 306916
rect 238708 306444 238772 306508
rect 238708 306232 238772 306236
rect 238708 306176 238722 306232
rect 238722 306176 238772 306232
rect 238708 306172 238772 306176
rect 377260 305900 377324 305964
rect 316540 305764 316604 305828
rect 327580 304948 327644 305012
rect 282868 304812 282932 304876
rect 320772 304812 320836 304876
rect 379468 304812 379532 304876
rect 304580 304676 304644 304740
rect 362908 304676 362972 304740
rect 367692 304540 367756 304604
rect 235580 304404 235644 304468
rect 363460 304404 363524 304468
rect 357572 304268 357636 304332
rect 350764 304132 350828 304196
rect 301084 303512 301148 303516
rect 301084 303456 301134 303512
rect 301134 303456 301148 303512
rect 301084 303452 301148 303456
rect 302924 303452 302988 303516
rect 373212 303316 373276 303380
rect 360700 303180 360764 303244
rect 239260 302228 239324 302292
rect 302556 302228 302620 302292
rect 302924 302228 302988 302292
rect 358860 302092 358924 302156
rect 304948 301956 305012 302020
rect 305500 301956 305564 302020
rect 383700 301956 383764 302020
rect 350580 301820 350644 301884
rect 240916 301684 240980 301748
rect 223804 301548 223868 301612
rect 246436 301548 246500 301612
rect 304948 301548 305012 301612
rect 235396 301412 235460 301476
rect 321508 301412 321572 301476
rect 274588 301276 274652 301340
rect 381492 300596 381556 300660
rect 302188 300248 302252 300252
rect 302188 300192 302238 300248
rect 302238 300192 302252 300248
rect 302188 300188 302252 300192
rect 238340 300052 238404 300116
rect 298140 300052 298204 300116
rect 368428 299372 368492 299436
rect 310468 299236 310532 299300
rect 311756 299236 311820 299300
rect 317276 299236 317340 299300
rect 376892 299236 376956 299300
rect 375420 299100 375484 299164
rect 228588 298964 228652 299028
rect 235028 298828 235092 298892
rect 233924 298692 233988 298756
rect 295012 298692 295076 298756
rect 304396 298012 304460 298076
rect 364380 298012 364444 298076
rect 359412 297876 359476 297940
rect 302740 297604 302804 297668
rect 238892 296788 238956 296852
rect 238708 296516 238772 296580
rect 226012 296380 226076 296444
rect 284340 296380 284404 296444
rect 226380 296244 226444 296308
rect 223068 296108 223132 296172
rect 226564 295972 226628 296036
rect 223620 295292 223684 295356
rect 349108 295156 349172 295220
rect 345060 295020 345124 295084
rect 229508 294884 229572 294948
rect 227300 294748 227364 294812
rect 285812 294748 285876 294812
rect 225276 294612 225340 294676
rect 285628 294612 285692 294676
rect 228404 294476 228468 294540
rect 232452 294340 232516 294404
rect 229876 294204 229940 294268
rect 288388 294204 288452 294268
rect 251956 293660 252020 293724
rect 310652 293660 310716 293724
rect 242940 293524 243004 293588
rect 302740 293524 302804 293588
rect 238156 293388 238220 293452
rect 239076 293252 239140 293316
rect 235948 293116 236012 293180
rect 215892 292572 215956 292636
rect 282132 292436 282196 292500
rect 221044 292164 221108 292228
rect 280660 292300 280724 292364
rect 218652 292028 218716 292092
rect 277900 291892 277964 291956
rect 248092 291756 248156 291820
rect 353892 291756 353956 291820
rect 220124 291484 220188 291548
rect 220308 291348 220372 291412
rect 221228 291212 221292 291276
rect 253060 290940 253124 291004
rect 312124 290940 312188 291004
rect 245148 290804 245212 290868
rect 253244 290668 253308 290732
rect 313780 290668 313844 290732
rect 262076 290532 262140 290596
rect 246252 290396 246316 290460
rect 238892 290124 238956 290188
rect 244228 290184 244292 290188
rect 244228 290128 244278 290184
rect 244278 290128 244292 290184
rect 244228 290124 244292 290128
rect 231532 289912 231596 289916
rect 231532 289856 231582 289912
rect 231582 289856 231596 289912
rect 231532 289852 231596 289856
rect 244228 289716 244292 289780
rect 244964 289716 245028 289780
rect 245332 289444 245396 289508
rect 249380 289172 249444 289236
rect 245332 289036 245396 289100
rect 231532 288356 231596 288420
rect 231532 287676 231596 287740
rect 269620 287676 269684 287740
rect 221044 286316 221108 286380
rect 220308 278020 220372 278084
rect 220124 276660 220188 276724
rect 221228 275164 221292 275228
rect 271092 273804 271156 273868
rect 260604 272444 260668 272508
rect 318932 272444 318996 272508
rect 266676 271084 266740 271148
rect 259316 268364 259380 268428
rect 317644 268364 317708 268428
rect 255636 267004 255700 267068
rect 257108 264420 257172 264484
rect 316356 264420 316420 264484
rect 264836 264284 264900 264348
rect 256372 264148 256436 264212
rect 259132 262788 259196 262852
rect 261892 261428 261956 261492
rect 320404 261428 320468 261492
rect 263548 258844 263612 258908
rect 323348 258844 323412 258908
rect 255452 258708 255516 258772
rect 260420 257212 260484 257276
rect 266124 255852 266188 255916
rect 324452 255852 324516 255916
rect 267412 253268 267476 253332
rect 261708 253132 261772 253196
rect 256004 251772 256068 251836
rect 263548 250548 263612 250612
rect 324636 250548 324700 250612
rect 266124 249052 266188 249116
rect 258948 247964 259012 248028
rect 263364 247692 263428 247756
rect 265388 246604 265452 246668
rect 317828 246468 317892 246532
rect 266124 246196 266188 246260
rect 323164 245108 323228 245172
rect 264284 244972 264348 245036
rect 256924 244836 256988 244900
rect 218652 243476 218716 243540
rect 267412 242252 267476 242316
rect 259500 242116 259564 242180
rect 245700 241980 245764 242044
rect 241836 241844 241900 241908
rect 222700 241708 222764 241772
rect 252692 241708 252756 241772
rect 225460 241572 225524 241636
rect 257292 241572 257356 241636
rect 269620 241572 269684 241636
rect 225644 241436 225708 241500
rect 247540 241436 247604 241500
rect 258580 241436 258644 241500
rect 224172 241300 224236 241364
rect 230796 241164 230860 241228
rect 232084 241028 232148 241092
rect 233372 241028 233436 241092
rect 292620 241028 292684 241092
rect 227668 240892 227732 240956
rect 229140 240756 229204 240820
rect 234844 240756 234908 240820
rect 294460 240756 294524 240820
rect 233188 240620 233252 240684
rect 233740 240620 233804 240684
rect 234476 240620 234540 240684
rect 237972 240620 238036 240684
rect 258396 240620 258460 240684
rect 259868 240620 259932 240684
rect 224172 240484 224236 240548
rect 230428 240484 230492 240548
rect 237788 240484 237852 240548
rect 222516 240348 222580 240412
rect 233004 240348 233068 240412
rect 239812 240212 239876 240276
rect 265204 240348 265268 240412
rect 274588 240620 274652 240684
rect 222516 239940 222580 240004
rect 223068 239940 223132 240004
rect 223804 239940 223868 240004
rect 223988 239940 224052 240004
rect 223252 239804 223316 239868
rect 226380 239940 226444 240004
rect 230980 240076 231044 240140
rect 241836 240076 241900 240140
rect 242020 240076 242084 240140
rect 246252 240076 246316 240140
rect 224172 239864 224236 239868
rect 224172 239808 224186 239864
rect 224186 239808 224236 239864
rect 224172 239804 224236 239808
rect 224724 239804 224788 239868
rect 225092 239864 225156 239868
rect 225092 239808 225096 239864
rect 225096 239808 225152 239864
rect 225152 239808 225156 239864
rect 225092 239804 225156 239808
rect 226196 239804 226260 239868
rect 227300 239804 227364 239868
rect 229508 239804 229572 239868
rect 230060 239804 230124 239868
rect 230980 239804 231044 239868
rect 231716 239804 231780 239868
rect 232636 239804 232700 239868
rect 232820 239804 232884 239868
rect 233372 239864 233436 239868
rect 233372 239808 233422 239864
rect 233422 239808 233436 239864
rect 233372 239804 233436 239808
rect 233924 239804 233988 239868
rect 223436 239668 223500 239732
rect 223620 239668 223684 239732
rect 225276 239532 225340 239596
rect 222700 239396 222764 239460
rect 226012 239396 226076 239460
rect 225644 239260 225708 239324
rect 226748 239668 226812 239732
rect 227668 239668 227732 239732
rect 228588 239668 228652 239732
rect 229140 239668 229204 239732
rect 229876 239668 229940 239732
rect 230796 239668 230860 239732
rect 231348 239668 231412 239732
rect 231532 239728 231596 239732
rect 231532 239672 231546 239728
rect 231546 239672 231596 239728
rect 231532 239668 231596 239672
rect 232084 239668 232148 239732
rect 233188 239668 233252 239732
rect 233740 239728 233804 239732
rect 233740 239672 233754 239728
rect 233754 239672 233804 239728
rect 233740 239668 233804 239672
rect 234108 239668 234172 239732
rect 226380 239532 226444 239596
rect 226564 239396 226628 239460
rect 227484 239456 227548 239460
rect 227484 239400 227498 239456
rect 227498 239400 227548 239456
rect 227484 239396 227548 239400
rect 227852 239396 227916 239460
rect 228956 239532 229020 239596
rect 229508 239592 229572 239596
rect 229508 239536 229558 239592
rect 229558 239536 229572 239592
rect 229508 239532 229572 239536
rect 231164 239532 231228 239596
rect 232268 239532 232332 239596
rect 233004 239532 233068 239596
rect 236684 239940 236748 240004
rect 234844 239864 234908 239868
rect 234844 239808 234848 239864
rect 234848 239808 234904 239864
rect 234904 239808 234908 239864
rect 234844 239804 234908 239808
rect 236868 239804 236932 239868
rect 237972 239804 238036 239868
rect 239628 239940 239692 240004
rect 239076 239804 239140 239868
rect 240180 239804 240244 239868
rect 240548 239804 240612 239868
rect 241100 239804 241164 239868
rect 235028 239728 235092 239732
rect 235028 239672 235078 239728
rect 235078 239672 235092 239728
rect 235028 239668 235092 239672
rect 235396 239668 235460 239732
rect 236132 239728 236196 239732
rect 236132 239672 236146 239728
rect 236146 239672 236196 239728
rect 236132 239668 236196 239672
rect 237236 239668 237300 239732
rect 238340 239668 238404 239732
rect 238708 239668 238772 239732
rect 242940 239668 243004 239732
rect 244964 239804 245028 239868
rect 245148 239804 245212 239868
rect 245884 239804 245948 239868
rect 249196 239940 249260 240004
rect 246436 239804 246500 239868
rect 248276 239804 248340 239868
rect 248644 239864 248708 239868
rect 248644 239808 248648 239864
rect 248648 239808 248704 239864
rect 248704 239808 248708 239864
rect 248644 239804 248708 239808
rect 249380 239804 249444 239868
rect 244596 239668 244660 239732
rect 245332 239668 245396 239732
rect 246804 239668 246868 239732
rect 247908 239668 247972 239732
rect 248460 239668 248524 239732
rect 250852 239804 250916 239868
rect 251956 239804 252020 239868
rect 252692 239804 252756 239868
rect 254900 239804 254964 239868
rect 250116 239668 250180 239732
rect 251772 239668 251836 239732
rect 253428 239668 253492 239732
rect 258396 240212 258460 240276
rect 256004 239804 256068 239868
rect 255452 239668 255516 239732
rect 257108 239728 257172 239732
rect 258396 239940 258460 240004
rect 261708 239804 261772 239868
rect 262444 239804 262508 239868
rect 262996 239804 263060 239868
rect 263548 239804 263612 239868
rect 263916 239804 263980 239868
rect 264836 239804 264900 239868
rect 265388 239864 265452 239868
rect 265388 239808 265392 239864
rect 265392 239808 265448 239864
rect 265448 239808 265452 239864
rect 265388 239804 265452 239808
rect 266308 239804 266372 239868
rect 257108 239672 257158 239728
rect 257158 239672 257172 239728
rect 257108 239668 257172 239672
rect 259500 239728 259564 239732
rect 259500 239672 259514 239728
rect 259514 239672 259564 239728
rect 259500 239668 259564 239672
rect 259684 239668 259748 239732
rect 260420 239668 260484 239732
rect 261524 239668 261588 239732
rect 262076 239668 262140 239732
rect 262260 239668 262324 239732
rect 263364 239668 263428 239732
rect 264100 239668 264164 239732
rect 265204 239668 265268 239732
rect 265756 239668 265820 239732
rect 266124 239668 266188 239732
rect 266676 239668 266740 239732
rect 228220 239396 228284 239460
rect 229324 239396 229388 239460
rect 230428 239396 230492 239460
rect 234292 239396 234356 239460
rect 235212 239396 235276 239460
rect 236316 239396 236380 239460
rect 237052 239456 237116 239460
rect 237052 239400 237066 239456
rect 237066 239400 237116 239456
rect 237052 239396 237116 239400
rect 238156 239396 238220 239460
rect 238524 239396 238588 239460
rect 238892 239456 238956 239460
rect 238892 239400 238942 239456
rect 238942 239400 238956 239456
rect 238892 239396 238956 239400
rect 239260 239456 239324 239460
rect 239260 239400 239310 239456
rect 239310 239400 239324 239456
rect 239260 239396 239324 239400
rect 239812 239396 239876 239460
rect 243124 239396 243188 239460
rect 244780 239396 244844 239460
rect 247540 239396 247604 239460
rect 248092 239396 248156 239460
rect 249564 239456 249628 239460
rect 249564 239400 249578 239456
rect 249578 239400 249628 239456
rect 249564 239396 249628 239400
rect 252324 239396 252388 239460
rect 253060 239456 253124 239460
rect 253060 239400 253074 239456
rect 253074 239400 253124 239456
rect 253060 239396 253124 239400
rect 253244 239396 253308 239460
rect 256372 239396 256436 239460
rect 257292 239396 257356 239460
rect 258580 239396 258644 239460
rect 259132 239396 259196 239460
rect 259316 239396 259380 239460
rect 261156 239396 261220 239460
rect 263364 239396 263428 239460
rect 263732 239396 263796 239460
rect 223804 238988 223868 239052
rect 225460 238988 225524 239052
rect 228404 238716 228468 238780
rect 231164 238776 231228 238780
rect 231164 238720 231178 238776
rect 231178 238720 231228 238776
rect 231164 238716 231228 238720
rect 232452 238716 232516 238780
rect 233740 238716 233804 238780
rect 235580 238716 235644 238780
rect 239444 238716 239508 238780
rect 240916 238716 240980 238780
rect 233924 238580 233988 238644
rect 241100 238640 241164 238644
rect 245700 238716 245764 238780
rect 249932 238716 249996 238780
rect 241100 238584 241150 238640
rect 241150 238584 241164 238640
rect 241100 238580 241164 238584
rect 245332 238640 245396 238644
rect 245332 238584 245382 238640
rect 245382 238584 245396 238640
rect 245332 238580 245396 238584
rect 250300 238580 250364 238644
rect 255636 238580 255700 238644
rect 256924 238716 256988 238780
rect 259500 238716 259564 238780
rect 260420 238776 260484 238780
rect 260420 238720 260434 238776
rect 260434 238720 260484 238776
rect 260420 238716 260484 238720
rect 260604 238716 260668 238780
rect 264100 238776 264164 238780
rect 264100 238720 264150 238776
rect 264150 238720 264164 238776
rect 264100 238716 264164 238720
rect 265388 238716 265452 238780
rect 271828 238716 271892 238780
rect 234292 238444 234356 238508
rect 259316 238444 259380 238508
rect 186820 238308 186884 238372
rect 175964 238172 176028 238236
rect 223988 238172 224052 238236
rect 227300 238172 227364 238236
rect 231716 238172 231780 238236
rect 233556 238172 233620 238236
rect 236132 238172 236196 238236
rect 236684 238172 236748 238236
rect 239260 238172 239324 238236
rect 241284 238172 241348 238236
rect 242388 238172 242452 238236
rect 258396 238308 258460 238372
rect 258948 238172 259012 238236
rect 259868 238308 259932 238372
rect 260604 238308 260668 238372
rect 263548 238232 263612 238236
rect 263548 238176 263598 238232
rect 263598 238176 263612 238232
rect 263548 238172 263612 238176
rect 185164 238036 185228 238100
rect 227116 238036 227180 238100
rect 234292 238036 234356 238100
rect 175780 237900 175844 237964
rect 230612 237900 230676 237964
rect 255452 237960 255516 237964
rect 255452 237904 255466 237960
rect 255466 237904 255516 237960
rect 255452 237900 255516 237904
rect 258764 238036 258828 238100
rect 262812 237900 262876 237964
rect 268332 237900 268396 237964
rect 229692 237764 229756 237828
rect 251036 237764 251100 237828
rect 230060 237492 230124 237556
rect 236868 237492 236932 237556
rect 239628 237492 239692 237556
rect 263180 237628 263244 237692
rect 271092 237628 271156 237692
rect 287652 237356 287716 237420
rect 265756 237144 265820 237148
rect 265756 237088 265770 237144
rect 265770 237088 265820 237144
rect 265756 237084 265820 237088
rect 268332 237084 268396 237148
rect 236500 236812 236564 236876
rect 239076 236676 239140 236740
rect 240732 236676 240796 236740
rect 241836 236736 241900 236740
rect 241836 236680 241886 236736
rect 241886 236680 241900 236736
rect 241836 236676 241900 236680
rect 249932 236736 249996 236740
rect 249932 236680 249946 236736
rect 249946 236680 249996 236736
rect 249932 236676 249996 236680
rect 252508 236676 252572 236740
rect 256372 236676 256436 236740
rect 258580 236676 258644 236740
rect 266124 236676 266188 236740
rect 232452 236540 232516 236604
rect 229692 236404 229756 236468
rect 248644 236404 248708 236468
rect 252876 236404 252940 236468
rect 224724 236268 224788 236332
rect 235212 236268 235276 236332
rect 237052 236132 237116 236196
rect 261340 236192 261404 236196
rect 261340 236136 261390 236192
rect 261390 236136 261404 236192
rect 261340 236132 261404 236136
rect 229876 235996 229940 236060
rect 233740 235996 233804 236060
rect 234476 235996 234540 236060
rect 226748 235860 226812 235924
rect 274588 235860 274652 235924
rect 328684 235860 328748 235924
rect 230612 235724 230676 235788
rect 232636 235724 232700 235788
rect 238524 235724 238588 235788
rect 253244 235724 253308 235788
rect 183140 235588 183204 235652
rect 261708 235588 261772 235652
rect 169524 235452 169588 235516
rect 176516 235180 176580 235244
rect 235028 235452 235092 235516
rect 239628 235452 239692 235516
rect 328868 235452 328932 235516
rect 244780 235316 244844 235380
rect 257108 235044 257172 235108
rect 261524 235044 261588 235108
rect 183324 234636 183388 234700
rect 243124 234636 243188 234700
rect 182956 234500 183020 234564
rect 261156 234500 261220 234564
rect 181484 234364 181548 234428
rect 254900 234364 254964 234428
rect 181300 234228 181364 234292
rect 250116 234228 250180 234292
rect 182772 234092 182836 234156
rect 173756 233956 173820 234020
rect 233372 233956 233436 234020
rect 180564 233820 180628 233884
rect 184428 233684 184492 233748
rect 235396 233684 235460 233748
rect 258580 233276 258644 233340
rect 165476 233140 165540 233204
rect 240548 233140 240612 233204
rect 246436 233140 246500 233204
rect 190868 233004 190932 233068
rect 175044 232868 175108 232932
rect 162900 232732 162964 232796
rect 193628 232732 193692 232796
rect 299980 232732 300044 232796
rect 163820 232596 163884 232660
rect 265756 232596 265820 232660
rect 330340 232596 330404 232660
rect 168236 232460 168300 232524
rect 191420 232324 191484 232388
rect 259500 232324 259564 232388
rect 192708 232188 192772 232252
rect 252140 232188 252204 232252
rect 262444 232188 262508 232252
rect 168052 231780 168116 231844
rect 227852 231644 227916 231708
rect 234476 231644 234540 231708
rect 172284 231508 172348 231572
rect 295932 231508 295996 231572
rect 174860 231372 174924 231436
rect 166764 231236 166828 231300
rect 170628 231100 170692 231164
rect 262996 230828 263060 230892
rect 166580 230012 166644 230076
rect 173572 229876 173636 229940
rect 225092 229740 225156 229804
rect 241836 230284 241900 230348
rect 262812 230208 262876 230212
rect 262812 230152 262862 230208
rect 262862 230152 262876 230208
rect 262812 230148 262876 230152
rect 310468 230148 310532 230212
rect 252508 230072 252572 230076
rect 252508 230016 252522 230072
rect 252522 230016 252572 230072
rect 252508 230012 252572 230016
rect 262444 229740 262508 229804
rect 327580 228652 327644 228716
rect 307708 228516 307772 228580
rect 252876 228380 252940 228444
rect 242388 228244 242452 228308
rect 249748 228244 249812 228308
rect 250852 228244 250916 228308
rect 258580 227564 258644 227628
rect 249748 227292 249812 227356
rect 328500 227292 328564 227356
rect 249196 227156 249260 227220
rect 190316 226884 190380 226948
rect 249196 226884 249260 226948
rect 181116 226340 181180 226404
rect 163452 225660 163516 225724
rect 246988 226204 247052 226268
rect 248276 226204 248340 226268
rect 260420 226204 260484 226268
rect 323532 226204 323596 226268
rect 243124 226068 243188 226132
rect 302556 226068 302620 226132
rect 227668 225932 227732 225996
rect 248276 225932 248340 225996
rect 306420 225932 306484 225996
rect 233740 225796 233804 225860
rect 234476 225524 234540 225588
rect 243124 224980 243188 225044
rect 180380 224300 180444 224364
rect 240180 224844 240244 224908
rect 261340 224708 261404 224772
rect 320220 224708 320284 224772
rect 246436 224436 246500 224500
rect 304212 224572 304276 224636
rect 251588 224300 251652 224364
rect 165292 224164 165356 224228
rect 246988 224164 247052 224228
rect 225092 223484 225156 223548
rect 263180 223484 263244 223548
rect 320772 223348 320836 223412
rect 300900 223212 300964 223276
rect 314332 223076 314396 223140
rect 178908 222804 178972 222868
rect 239628 222940 239692 223004
rect 240732 222804 240796 222868
rect 251036 222124 251100 222188
rect 256372 221988 256436 222052
rect 308260 221988 308324 222052
rect 233188 221852 233252 221916
rect 233556 221852 233620 221916
rect 263364 221716 263428 221780
rect 180932 221580 180996 221644
rect 233188 221444 233252 221508
rect 260972 221444 261036 221508
rect 264100 221308 264164 221372
rect 170076 220356 170140 220420
rect 230428 220628 230492 220692
rect 231164 220628 231228 220692
rect 230980 220492 231044 220556
rect 231532 220492 231596 220556
rect 290596 220356 290660 220420
rect 174676 220220 174740 220284
rect 314884 220220 314948 220284
rect 230428 220084 230492 220148
rect 250300 219268 250364 219332
rect 315068 219132 315132 219196
rect 165108 218860 165172 218924
rect 247540 218860 247604 218924
rect 306972 218996 307036 219060
rect 253428 218860 253492 218924
rect 312308 218860 312372 218924
rect 163636 218724 163700 218788
rect 250300 218724 250364 218788
rect 179092 218588 179156 218652
rect 238892 218588 238956 218652
rect 246804 218588 246868 218652
rect 253428 218044 253492 218108
rect 166396 217908 166460 217972
rect 167868 217772 167932 217836
rect 170444 217636 170508 217700
rect 167684 217500 167748 217564
rect 169340 217364 169404 217428
rect 170260 217228 170324 217292
rect 172100 217092 172164 217156
rect 171916 215868 171980 215932
rect 176148 215052 176212 215116
rect 195836 214916 195900 214980
rect 191236 214780 191300 214844
rect 195652 214644 195716 214708
rect 192892 214508 192956 214572
rect 180196 213828 180260 213892
rect 177620 213692 177684 213756
rect 173388 213556 173452 213620
rect 184612 213420 184676 213484
rect 173204 213284 173268 213348
rect 174492 213148 174556 213212
rect 177804 213012 177868 213076
rect 215892 212060 215956 212124
rect 169156 211924 169220 211988
rect 180012 211788 180076 211852
rect 239444 211788 239508 211852
rect 161980 211108 162044 211172
rect 162716 211108 162780 211172
rect 203380 211108 203444 211172
rect 164740 209612 164804 209676
rect 166212 209612 166276 209676
rect 184060 209612 184124 209676
rect 171180 209476 171244 209540
rect 183876 209476 183940 209540
rect 188292 209476 188356 209540
rect 191052 209476 191116 209540
rect 192340 209476 192404 209540
rect 193996 209476 194060 209540
rect 195468 209476 195532 209540
rect 196756 209612 196820 209676
rect 197860 209612 197924 209676
rect 199332 209612 199396 209676
rect 199700 209612 199764 209676
rect 196388 209476 196452 209540
rect 196572 209340 196636 209404
rect 199516 209476 199580 209540
rect 198596 207572 198660 207636
rect 256740 207572 256804 207636
rect 203380 201316 203444 201380
rect 205956 190980 206020 191044
rect 207612 182820 207676 182884
rect 204116 179964 204180 180028
rect 207980 178604 208044 178668
rect 205404 177244 205468 177308
rect 209084 173300 209148 173364
rect 207796 173164 207860 173228
rect 206876 171668 206940 171732
rect 209268 169084 209332 169148
rect 205220 168948 205284 169012
rect 263916 168948 263980 169012
rect 204668 165956 204732 166020
rect 203932 165004 203996 165068
rect 206508 164868 206572 164932
rect 203564 163508 203628 163572
rect 204852 163372 204916 163436
rect 206692 162148 206756 162212
rect 203196 162012 203260 162076
rect 170996 161876 171060 161940
rect 201356 161876 201420 161940
rect 169156 161740 169220 161804
rect 197860 161196 197924 161260
rect 164372 160788 164436 160852
rect 165108 160788 165172 160852
rect 167132 160652 167196 160716
rect 175964 160652 176028 160716
rect 167316 160516 167380 160580
rect 166028 160380 166092 160444
rect 163820 159836 163884 159900
rect 163268 159700 163332 159764
rect 163636 159564 163700 159628
rect 167132 160108 167196 160172
rect 164372 159836 164436 159900
rect 166764 159972 166828 160036
rect 186820 160788 186884 160852
rect 181484 160244 181548 160308
rect 169340 159972 169404 160036
rect 164924 159836 164988 159900
rect 166396 159836 166460 159900
rect 166580 159836 166644 159900
rect 167316 159836 167380 159900
rect 167868 159836 167932 159900
rect 168972 159836 169036 159900
rect 165292 159700 165356 159764
rect 165476 159760 165540 159764
rect 165476 159704 165526 159760
rect 165526 159704 165540 159760
rect 165476 159700 165540 159704
rect 166212 159760 166276 159764
rect 166212 159704 166226 159760
rect 166226 159704 166276 159760
rect 166212 159700 166276 159704
rect 167684 159700 167748 159764
rect 168604 159700 168668 159764
rect 169156 159700 169220 159764
rect 169524 159700 169588 159764
rect 166028 159564 166092 159628
rect 168236 159564 168300 159628
rect 170076 159836 170140 159900
rect 170628 159836 170692 159900
rect 172284 159972 172348 160036
rect 171916 159836 171980 159900
rect 173204 159972 173268 160036
rect 172836 159896 172900 159900
rect 172836 159840 172886 159896
rect 172886 159840 172900 159896
rect 170628 159760 170692 159764
rect 170628 159704 170642 159760
rect 170642 159704 170692 159760
rect 170628 159700 170692 159704
rect 170996 159760 171060 159764
rect 170996 159704 171010 159760
rect 171010 159704 171060 159760
rect 170996 159700 171060 159704
rect 172100 159700 172164 159764
rect 172836 159836 172900 159840
rect 173388 159836 173452 159900
rect 173572 159836 173636 159900
rect 175044 159972 175108 160036
rect 180748 159972 180812 160036
rect 203380 160788 203444 160852
rect 202828 160516 202892 160580
rect 245700 160516 245764 160580
rect 174860 159836 174924 159900
rect 176516 159836 176580 159900
rect 177620 159836 177684 159900
rect 178908 159896 178972 159900
rect 178908 159840 178958 159896
rect 178958 159840 178972 159896
rect 178908 159836 178972 159840
rect 180012 159896 180076 159900
rect 180012 159840 180062 159896
rect 180062 159840 180076 159896
rect 180012 159836 180076 159840
rect 180380 159896 180444 159900
rect 180380 159840 180394 159896
rect 180394 159840 180444 159896
rect 180380 159836 180444 159840
rect 180564 159896 180628 159900
rect 180564 159840 180614 159896
rect 180614 159840 180628 159896
rect 180564 159836 180628 159840
rect 180932 159836 180996 159900
rect 181300 159836 181364 159900
rect 173020 159700 173084 159764
rect 173388 159760 173452 159764
rect 173388 159704 173438 159760
rect 173438 159704 173452 159760
rect 173388 159700 173452 159704
rect 173756 159700 173820 159764
rect 170444 159564 170508 159628
rect 174676 159700 174740 159764
rect 176884 159700 176948 159764
rect 177804 159700 177868 159764
rect 179092 159700 179156 159764
rect 180196 159700 180260 159764
rect 181484 159700 181548 159764
rect 182588 159972 182652 160036
rect 183140 159972 183204 160036
rect 182772 159896 182836 159900
rect 182772 159840 182822 159896
rect 182822 159840 182836 159896
rect 182772 159836 182836 159840
rect 183324 159896 183388 159900
rect 183324 159840 183338 159896
rect 183338 159840 183388 159896
rect 183324 159836 183388 159840
rect 184612 159972 184676 160036
rect 184428 159836 184492 159900
rect 188292 159896 188356 159900
rect 188292 159840 188342 159896
rect 188342 159840 188356 159896
rect 188292 159836 188356 159840
rect 190868 159972 190932 160036
rect 190316 159836 190380 159900
rect 191052 159836 191116 159900
rect 196388 159972 196452 160036
rect 192340 159836 192404 159900
rect 192892 159836 192956 159900
rect 193812 159836 193876 159900
rect 194180 159836 194244 159900
rect 195100 159836 195164 159900
rect 195468 159836 195532 159900
rect 195652 159836 195716 159900
rect 196572 159836 196636 159900
rect 197860 160108 197924 160172
rect 198412 159836 198476 159900
rect 199700 160108 199764 160172
rect 199516 159972 199580 160036
rect 199332 159896 199396 159900
rect 199332 159840 199382 159896
rect 199382 159840 199396 159896
rect 199332 159836 199396 159840
rect 201356 159896 201420 159900
rect 201356 159840 201370 159896
rect 201370 159840 201420 159896
rect 201356 159836 201420 159840
rect 203564 159896 203628 159900
rect 203564 159840 203578 159896
rect 203578 159840 203628 159896
rect 203564 159836 203628 159840
rect 204116 159836 204180 159900
rect 205036 159836 205100 159900
rect 205404 159836 205468 159900
rect 182956 159700 183020 159764
rect 183324 159760 183388 159764
rect 183324 159704 183374 159760
rect 183374 159704 183388 159760
rect 183324 159700 183388 159704
rect 184060 159700 184124 159764
rect 191420 159700 191484 159764
rect 192708 159700 192772 159764
rect 195836 159700 195900 159764
rect 196940 159700 197004 159764
rect 198596 159700 198660 159764
rect 203196 159700 203260 159764
rect 203380 159760 203444 159764
rect 203380 159704 203430 159760
rect 203430 159704 203444 159760
rect 203380 159700 203444 159704
rect 203932 159700 203996 159764
rect 204852 159700 204916 159764
rect 205956 159836 206020 159900
rect 206508 159896 206572 159900
rect 206508 159840 206558 159896
rect 206558 159840 206572 159896
rect 206508 159836 206572 159840
rect 206876 159896 206940 159900
rect 206876 159840 206890 159896
rect 206890 159840 206940 159896
rect 206876 159836 206940 159840
rect 207796 159836 207860 159900
rect 207612 159700 207676 159764
rect 172652 159564 172716 159628
rect 174492 159564 174556 159628
rect 175780 159428 175844 159492
rect 168604 159292 168668 159356
rect 183876 159428 183940 159492
rect 191236 159428 191300 159492
rect 176884 159292 176948 159356
rect 185164 159292 185228 159356
rect 165844 159080 165908 159084
rect 165844 159024 165894 159080
rect 165894 159024 165908 159080
rect 165844 159020 165908 159024
rect 201356 159080 201420 159084
rect 201356 159024 201406 159080
rect 201406 159024 201420 159080
rect 201356 159020 201420 159024
rect 204668 159020 204732 159084
rect 168604 158944 168668 158948
rect 168604 158888 168618 158944
rect 168618 158888 168668 158944
rect 168604 158884 168668 158888
rect 173020 158884 173084 158948
rect 176516 158748 176580 158812
rect 186452 158748 186516 158812
rect 163084 158672 163148 158676
rect 163084 158616 163098 158672
rect 163098 158616 163148 158672
rect 163084 158612 163148 158616
rect 164924 158612 164988 158676
rect 166764 158672 166828 158676
rect 166764 158616 166814 158672
rect 166814 158616 166828 158672
rect 166764 158612 166828 158616
rect 168052 158612 168116 158676
rect 168420 158612 168484 158676
rect 169524 158612 169588 158676
rect 170076 158612 170140 158676
rect 171548 158612 171612 158676
rect 171916 158612 171980 158676
rect 173572 158612 173636 158676
rect 174676 158672 174740 158676
rect 174676 158616 174690 158672
rect 174690 158616 174740 158672
rect 174676 158612 174740 158616
rect 176148 158612 176212 158676
rect 163452 158476 163516 158540
rect 165292 158476 165356 158540
rect 165660 158476 165724 158540
rect 177620 158672 177684 158676
rect 177620 158616 177634 158672
rect 177634 158616 177684 158672
rect 177620 158612 177684 158616
rect 178724 158612 178788 158676
rect 179828 158612 179892 158676
rect 180564 158612 180628 158676
rect 181116 158612 181180 158676
rect 182956 158612 183020 158676
rect 183140 158672 183204 158676
rect 183140 158616 183154 158672
rect 183154 158616 183204 158672
rect 183140 158612 183204 158616
rect 184980 158672 185044 158676
rect 184980 158616 185030 158672
rect 185030 158616 185044 158672
rect 184980 158612 185044 158616
rect 185164 158612 185228 158676
rect 187004 158612 187068 158676
rect 187372 158612 187436 158676
rect 187556 158672 187620 158676
rect 187556 158616 187570 158672
rect 187570 158616 187620 158672
rect 187556 158612 187620 158616
rect 188476 158612 188540 158676
rect 188660 158672 188724 158676
rect 188660 158616 188674 158672
rect 188674 158616 188724 158672
rect 188660 158612 188724 158616
rect 189764 158612 189828 158676
rect 189948 158672 190012 158676
rect 189948 158616 189998 158672
rect 189998 158616 190012 158672
rect 189948 158612 190012 158616
rect 190132 158612 190196 158676
rect 191236 158612 191300 158676
rect 192708 158612 192772 158676
rect 192892 158612 192956 158676
rect 193996 158612 194060 158676
rect 195284 158612 195348 158676
rect 195836 158672 195900 158676
rect 195836 158616 195886 158672
rect 195886 158616 195900 158672
rect 195836 158612 195900 158616
rect 196204 158612 196268 158676
rect 196756 158612 196820 158676
rect 198228 158672 198292 158676
rect 198228 158616 198278 158672
rect 198278 158616 198292 158672
rect 198228 158612 198292 158616
rect 199332 158612 199396 158676
rect 199884 158672 199948 158676
rect 199884 158616 199898 158672
rect 199898 158616 199948 158672
rect 199884 158612 199948 158616
rect 200620 158612 200684 158676
rect 200988 158672 201052 158676
rect 200988 158616 201002 158672
rect 201002 158616 201052 158672
rect 200988 158612 201052 158616
rect 202644 158612 202708 158676
rect 203748 158612 203812 158676
rect 203932 158672 203996 158676
rect 203932 158616 203982 158672
rect 203982 158616 203996 158672
rect 203932 158612 203996 158616
rect 205036 158612 205100 158676
rect 209084 158612 209148 158676
rect 162900 158340 162964 158404
rect 168236 158340 168300 158404
rect 166948 158204 167012 158268
rect 168972 158204 169036 158268
rect 170996 158340 171060 158404
rect 171180 158340 171244 158404
rect 175044 158340 175108 158404
rect 175964 158340 176028 158404
rect 198044 158340 198108 158404
rect 199516 158340 199580 158404
rect 201172 158340 201236 158404
rect 201356 158400 201420 158404
rect 201356 158344 201406 158400
rect 201406 158344 201420 158400
rect 201356 158340 201420 158344
rect 202460 158340 202524 158404
rect 204668 158340 204732 158404
rect 169892 158204 169956 158268
rect 170628 158204 170692 158268
rect 173388 158204 173452 158268
rect 174492 158204 174556 158268
rect 165844 158068 165908 158132
rect 168604 158068 168668 158132
rect 170260 158068 170324 158132
rect 170812 158068 170876 158132
rect 176332 158068 176396 158132
rect 206692 158204 206756 158268
rect 177436 158068 177500 158132
rect 181484 158068 181548 158132
rect 187188 158068 187252 158132
rect 194364 158068 194428 158132
rect 195468 158068 195532 158132
rect 196388 158068 196452 158132
rect 207980 158068 208044 158132
rect 177252 157932 177316 157996
rect 201356 157932 201420 157996
rect 202092 157932 202156 157996
rect 244780 157932 244844 157996
rect 164372 157856 164436 157860
rect 164372 157800 164386 157856
rect 164386 157800 164436 157856
rect 164372 157796 164436 157800
rect 177988 157796 178052 157860
rect 186452 157796 186516 157860
rect 166764 157660 166828 157724
rect 168236 157660 168300 157724
rect 202828 157660 202892 157724
rect 209268 157660 209332 157724
rect 169708 157524 169772 157588
rect 192340 157584 192404 157588
rect 192340 157528 192390 157584
rect 192390 157528 192404 157584
rect 192340 157524 192404 157528
rect 200804 157388 200868 157452
rect 164372 157252 164436 157316
rect 170444 157252 170508 157316
rect 173756 157252 173820 157316
rect 188292 157252 188356 157316
rect 192340 157312 192404 157316
rect 192340 157256 192390 157312
rect 192390 157256 192404 157312
rect 162900 157116 162964 157180
rect 192340 157252 192404 157256
rect 199884 157116 199948 157180
rect 168420 156844 168484 156908
rect 163268 156436 163332 156500
rect 202276 156028 202340 156092
rect 195284 155348 195348 155412
rect 199700 154532 199764 154596
rect 200988 154124 201052 154188
rect 177988 153988 178052 154052
rect 203932 153852 203996 153916
rect 174676 153716 174740 153780
rect 171732 153036 171796 153100
rect 176148 153096 176212 153100
rect 176148 153040 176198 153096
rect 176198 153040 176212 153096
rect 176148 153036 176212 153040
rect 175964 152900 176028 152964
rect 199332 152900 199396 152964
rect 258580 152900 258644 152964
rect 236500 152628 236564 152692
rect 199332 152492 199396 152556
rect 199700 152492 199764 152556
rect 198044 152356 198108 152420
rect 196756 152220 196820 152284
rect 226932 151132 226996 151196
rect 178908 150996 178972 151060
rect 172836 149908 172900 149972
rect 170076 149772 170140 149836
rect 177436 149772 177500 149836
rect 173572 149500 173636 149564
rect 175964 149092 176028 149156
rect 178724 148548 178788 148612
rect 173572 148412 173636 148476
rect 171180 147596 171244 147660
rect 265572 147596 265636 147660
rect 169892 147460 169956 147524
rect 174492 147460 174556 147524
rect 233740 147460 233804 147524
rect 173756 147324 173820 147388
rect 177620 147188 177684 147252
rect 232452 147052 232516 147116
rect 202644 146236 202708 146300
rect 262812 146236 262876 146300
rect 201356 146100 201420 146164
rect 203748 145964 203812 146028
rect 262260 145964 262324 146028
rect 202460 145828 202524 145892
rect 261156 145828 261220 145892
rect 205036 145692 205100 145756
rect 163084 145556 163148 145620
rect 235212 144740 235276 144804
rect 187004 144604 187068 144668
rect 171548 144468 171612 144532
rect 230980 144468 231044 144532
rect 196204 144332 196268 144396
rect 200620 144332 200684 144396
rect 202092 144332 202156 144396
rect 259684 144332 259748 144396
rect 199516 143924 199580 143988
rect 199884 143924 199948 143988
rect 202276 144060 202340 144124
rect 201172 143788 201236 143852
rect 261340 143788 261404 143852
rect 189764 143380 189828 143444
rect 248460 143380 248524 143444
rect 189948 143244 190012 143308
rect 187188 143108 187252 143172
rect 242020 143108 242084 143172
rect 187372 142972 187436 143036
rect 188660 142836 188724 142900
rect 255820 142836 255884 142900
rect 185164 142700 185228 142764
rect 187556 142564 187620 142628
rect 181484 142020 181548 142084
rect 181116 141884 181180 141948
rect 240732 141884 240796 141948
rect 183140 141748 183204 141812
rect 238708 141748 238772 141812
rect 268332 141748 268396 141812
rect 188476 141612 188540 141676
rect 177804 141476 177868 141540
rect 192892 141476 192956 141540
rect 174492 141340 174556 141404
rect 177804 141340 177868 141404
rect 177252 140796 177316 140860
rect 177804 140796 177868 140860
rect 184980 140796 185044 140860
rect 198228 140660 198292 140724
rect 168236 140524 168300 140588
rect 173020 139980 173084 140044
rect 179092 139980 179156 140044
rect 194364 139164 194428 139228
rect 257108 139164 257172 139228
rect 195468 139028 195532 139092
rect 254900 139028 254964 139092
rect 191236 138892 191300 138956
rect 190132 138756 190196 138820
rect 193996 138620 194060 138684
rect 192708 138484 192772 138548
rect 271828 137940 271892 138004
rect 168236 137260 168300 137324
rect 171732 136036 171796 136100
rect 168972 135900 169036 135964
rect 165660 131684 165724 131748
rect 168604 130460 168668 130524
rect 164372 130324 164436 130388
rect 182956 130324 183020 130388
rect 182588 127604 182652 127668
rect 172468 126380 172532 126444
rect 168420 126244 168484 126308
rect 180380 124748 180444 124812
rect 169708 122164 169772 122228
rect 181116 122164 181180 122228
rect 162900 122028 162964 122092
rect 203748 122028 203812 122092
rect 180012 120940 180076 121004
rect 195284 120804 195348 120868
rect 205036 120668 205100 120732
rect 196756 117948 196820 118012
rect 177436 116452 177500 116516
rect 198044 116452 198108 116516
rect 199700 115092 199764 115156
rect 165844 113732 165908 113796
rect 189764 113732 189828 113796
rect 180748 112372 180812 112436
rect 200988 111012 201052 111076
rect 184612 109652 184676 109716
rect 184428 108292 184492 108356
rect 187004 106932 187068 106996
rect 201172 106796 201236 106860
rect 202276 105436 202340 105500
rect 202460 104076 202524 104140
rect 191052 102852 191116 102916
rect 202644 102716 202708 102780
rect 187188 100132 187252 100196
rect 161980 99996 162044 100060
rect 179828 98772 179892 98836
rect 176516 98636 176580 98700
rect 203196 98636 203260 98700
rect 183140 97276 183204 97340
rect 204116 97140 204180 97204
rect 181484 95916 181548 95980
rect 205220 95780 205284 95844
rect 184060 94420 184124 94484
rect 205404 93060 205468 93124
rect 193812 82044 193876 82108
rect 198228 76468 198292 76532
rect 188292 72388 188356 72452
rect 281396 71844 281460 71908
rect 162716 71028 162780 71092
rect 187372 69532 187436 69596
rect 189948 64092 190012 64156
rect 191236 62732 191300 62796
rect 191420 61372 191484 61436
rect 333100 59332 333164 59396
rect 190868 58516 190932 58580
rect 193996 54436 194060 54500
rect 194180 53076 194244 53140
rect 201356 39204 201420 39268
rect 183324 32404 183388 32468
rect 331812 31724 331876 31788
rect 177620 28188 177684 28252
rect 183876 26828 183940 26892
rect 194364 21252 194428 21316
rect 177804 17172 177868 17236
rect 195652 14452 195716 14516
rect 187556 12956 187620 13020
rect 190132 9420 190196 9484
rect 195468 9284 195532 9348
rect 195100 9148 195164 9212
rect 196572 9012 196636 9076
rect 196940 8876 197004 8940
rect 188476 6836 188540 6900
rect 188844 6700 188908 6764
rect 188660 6564 188724 6628
rect 192708 6428 192772 6492
rect 192524 6292 192588 6356
rect 192892 6156 192956 6220
rect 185164 6020 185228 6084
rect 190316 3708 190380 3772
rect 353340 3708 353404 3772
rect 198596 3572 198660 3636
rect 198412 3436 198476 3500
rect 199884 3300 199948 3364
<< metal4 >>
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691174 -2346 705242
rect -2966 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 -2346 691174
rect -2966 690854 -2346 690938
rect -2966 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 -2346 690854
rect -2966 655174 -2346 690618
rect -2966 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 -2346 655174
rect -2966 654854 -2346 654938
rect -2966 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 -2346 654854
rect -2966 619174 -2346 654618
rect -2966 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 -2346 619174
rect -2966 618854 -2346 618938
rect -2966 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 -2346 618854
rect -2966 583174 -2346 618618
rect -2966 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 -2346 583174
rect -2966 582854 -2346 582938
rect -2966 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 -2346 582854
rect -2966 547174 -2346 582618
rect -2966 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 -2346 547174
rect -2966 546854 -2346 546938
rect -2966 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 -2346 546854
rect -2966 511174 -2346 546618
rect -2966 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 -2346 511174
rect -2966 510854 -2346 510938
rect -2966 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 -2346 510854
rect -2966 475174 -2346 510618
rect -2966 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 -2346 475174
rect -2966 474854 -2346 474938
rect -2966 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 -2346 474854
rect -2966 439174 -2346 474618
rect -2966 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 -2346 439174
rect -2966 438854 -2346 438938
rect -2966 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 -2346 438854
rect -2966 403174 -2346 438618
rect -2966 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 -2346 403174
rect -2966 402854 -2346 402938
rect -2966 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 -2346 402854
rect -2966 367174 -2346 402618
rect -2966 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 -2346 367174
rect -2966 366854 -2346 366938
rect -2966 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 -2346 366854
rect -2966 331174 -2346 366618
rect -2966 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 -2346 331174
rect -2966 330854 -2346 330938
rect -2966 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 -2346 330854
rect -2966 295174 -2346 330618
rect -2966 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 -2346 295174
rect -2966 294854 -2346 294938
rect -2966 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 -2346 294854
rect -2966 259174 -2346 294618
rect -2966 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 -2346 259174
rect -2966 258854 -2346 258938
rect -2966 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 -2346 258854
rect -2966 223174 -2346 258618
rect -2966 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 -2346 223174
rect -2966 222854 -2346 222938
rect -2966 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 -2346 222854
rect -2966 187174 -2346 222618
rect -2966 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 -2346 187174
rect -2966 186854 -2346 186938
rect -2966 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 -2346 186854
rect -2966 151174 -2346 186618
rect -2966 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 -2346 151174
rect -2966 150854 -2346 150938
rect -2966 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 -2346 150854
rect -2966 115174 -2346 150618
rect -2966 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 -2346 115174
rect -2966 114854 -2346 114938
rect -2966 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 -2346 114854
rect -2966 79174 -2346 114618
rect -2966 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 -2346 79174
rect -2966 78854 -2346 78938
rect -2966 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 -2346 78854
rect -2966 43174 -2346 78618
rect -2966 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 -2346 43174
rect -2966 42854 -2346 42938
rect -2966 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 -2346 42854
rect -2966 7174 -2346 42618
rect -2966 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 -2346 7174
rect -2966 6854 -2346 6938
rect -2966 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 -2346 6854
rect -2966 -1306 -2346 6618
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 705798 6134 705830
rect 5514 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 6134 705798
rect 5514 705478 6134 705562
rect 5514 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 6134 705478
rect 5514 691174 6134 705242
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect 5514 -1306 6134 6618
rect 5514 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 6134 -1306
rect 5514 -1626 6134 -1542
rect 5514 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 6134 -1626
rect 5514 -1894 6134 -1862
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 705798 42134 705830
rect 41514 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 42134 705798
rect 41514 705478 42134 705562
rect 41514 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 42134 705478
rect 41514 691174 42134 705242
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -1306 42134 6618
rect 41514 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 42134 -1306
rect 41514 -1626 42134 -1542
rect 41514 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 42134 -1626
rect 41514 -1894 42134 -1862
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 705798 78134 705830
rect 77514 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 78134 705798
rect 77514 705478 78134 705562
rect 77514 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 78134 705478
rect 77514 691174 78134 705242
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583174 78134 618618
rect 77514 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 78134 583174
rect 77514 582854 78134 582938
rect 77514 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 78134 582854
rect 77514 547174 78134 582618
rect 77514 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 78134 547174
rect 77514 546854 78134 546938
rect 77514 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 78134 546854
rect 77514 511174 78134 546618
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 439174 78134 474618
rect 77514 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 78134 439174
rect 77514 438854 78134 438938
rect 77514 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 78134 438854
rect 77514 403174 78134 438618
rect 77514 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 78134 403174
rect 77514 402854 78134 402938
rect 77514 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 78134 402854
rect 77514 367174 78134 402618
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 331174 78134 366618
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77514 295174 78134 330618
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 259174 78134 294618
rect 77514 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 78134 259174
rect 77514 258854 78134 258938
rect 77514 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 78134 258854
rect 77514 223174 78134 258618
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 151174 78134 186618
rect 77514 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 78134 151174
rect 77514 150854 78134 150938
rect 77514 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 78134 150854
rect 77514 115174 78134 150618
rect 77514 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 78134 115174
rect 77514 114854 78134 114938
rect 77514 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 78134 114854
rect 77514 79174 78134 114618
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -1306 78134 6618
rect 77514 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 78134 -1306
rect 77514 -1626 78134 -1542
rect 77514 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 78134 -1626
rect 77514 -1894 78134 -1862
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 705798 114134 705830
rect 113514 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 114134 705798
rect 113514 705478 114134 705562
rect 113514 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 114134 705478
rect 113514 691174 114134 705242
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 439174 114134 474618
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 113514 403174 114134 438618
rect 113514 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 114134 403174
rect 113514 402854 114134 402938
rect 113514 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 114134 402854
rect 113514 367174 114134 402618
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 331174 114134 366618
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 113514 295174 114134 330618
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 113514 259174 114134 294618
rect 113514 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 114134 259174
rect 113514 258854 114134 258938
rect 113514 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 114134 258854
rect 113514 223174 114134 258618
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 187174 114134 222618
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 113514 151174 114134 186618
rect 113514 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 114134 151174
rect 113514 150854 114134 150938
rect 113514 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 114134 150854
rect 113514 115174 114134 150618
rect 113514 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 114134 115174
rect 113514 114854 114134 114938
rect 113514 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 114134 114854
rect 113514 79174 114134 114618
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -1306 114134 6618
rect 113514 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 114134 -1306
rect 113514 -1626 114134 -1542
rect 113514 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 114134 -1626
rect 113514 -1894 114134 -1862
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 705798 150134 705830
rect 149514 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 150134 705798
rect 149514 705478 150134 705562
rect 149514 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 150134 705478
rect 149514 691174 150134 705242
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 149514 295174 150134 330618
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 149514 259174 150134 294618
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 223174 150134 258618
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 175963 238236 176029 238237
rect 175963 238172 175964 238236
rect 176028 238172 176029 238236
rect 175963 238171 176029 238172
rect 175779 237964 175845 237965
rect 175779 237900 175780 237964
rect 175844 237900 175845 237964
rect 175779 237899 175845 237900
rect 169523 235516 169589 235517
rect 169523 235452 169524 235516
rect 169588 235452 169589 235516
rect 169523 235451 169589 235452
rect 165475 233204 165541 233205
rect 165475 233140 165476 233204
rect 165540 233140 165541 233204
rect 165475 233139 165541 233140
rect 162899 232796 162965 232797
rect 162899 232732 162900 232796
rect 162964 232732 162965 232796
rect 162899 232731 162965 232732
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 187174 150134 222618
rect 161979 211172 162045 211173
rect 161979 211108 161980 211172
rect 162044 211108 162045 211172
rect 161979 211107 162045 211108
rect 162715 211172 162781 211173
rect 162715 211108 162716 211172
rect 162780 211108 162781 211172
rect 162715 211107 162781 211108
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 149514 151174 150134 186618
rect 149514 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 150134 151174
rect 149514 150854 150134 150938
rect 149514 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 150134 150854
rect 149514 115174 150134 150618
rect 149514 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 150134 115174
rect 149514 114854 150134 114938
rect 149514 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 150134 114854
rect 149514 79174 150134 114618
rect 161982 100061 162042 211107
rect 161979 100060 162045 100061
rect 161979 99996 161980 100060
rect 162044 99996 162045 100060
rect 161979 99995 162045 99996
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 162718 71093 162778 211107
rect 162902 158405 162962 232731
rect 163819 232660 163885 232661
rect 163819 232596 163820 232660
rect 163884 232596 163885 232660
rect 163819 232595 163885 232596
rect 163451 225724 163517 225725
rect 163451 225660 163452 225724
rect 163516 225660 163517 225724
rect 163451 225659 163517 225660
rect 163267 159764 163333 159765
rect 163267 159700 163268 159764
rect 163332 159700 163333 159764
rect 163267 159699 163333 159700
rect 163083 158676 163149 158677
rect 163083 158612 163084 158676
rect 163148 158612 163149 158676
rect 163083 158611 163149 158612
rect 162899 158404 162965 158405
rect 162899 158340 162900 158404
rect 162964 158340 162965 158404
rect 162899 158339 162965 158340
rect 162899 157180 162965 157181
rect 162899 157116 162900 157180
rect 162964 157116 162965 157180
rect 162899 157115 162965 157116
rect 162902 122093 162962 157115
rect 163086 145621 163146 158611
rect 163270 156501 163330 159699
rect 163454 158541 163514 225659
rect 163635 218788 163701 218789
rect 163635 218724 163636 218788
rect 163700 218724 163701 218788
rect 163635 218723 163701 218724
rect 163638 159629 163698 218723
rect 163822 159901 163882 232595
rect 165291 224228 165357 224229
rect 165291 224164 165292 224228
rect 165356 224164 165357 224228
rect 165291 224163 165357 224164
rect 165107 218924 165173 218925
rect 165107 218860 165108 218924
rect 165172 218860 165173 218924
rect 165107 218859 165173 218860
rect 164739 209676 164805 209677
rect 164739 209612 164740 209676
rect 164804 209612 164805 209676
rect 164739 209611 164805 209612
rect 164208 183454 164528 183486
rect 164208 183218 164250 183454
rect 164486 183218 164528 183454
rect 164208 183134 164528 183218
rect 164208 182898 164250 183134
rect 164486 182898 164528 183134
rect 164208 182866 164528 182898
rect 164742 167010 164802 209611
rect 164742 166950 164986 167010
rect 164371 160852 164437 160853
rect 164371 160788 164372 160852
rect 164436 160788 164437 160852
rect 164371 160787 164437 160788
rect 164374 159901 164434 160787
rect 164926 159901 164986 166950
rect 165110 160853 165170 218859
rect 165107 160852 165173 160853
rect 165107 160788 165108 160852
rect 165172 160788 165173 160852
rect 165107 160787 165173 160788
rect 163819 159900 163885 159901
rect 163819 159836 163820 159900
rect 163884 159836 163885 159900
rect 163819 159835 163885 159836
rect 164371 159900 164437 159901
rect 164371 159836 164372 159900
rect 164436 159836 164437 159900
rect 164371 159835 164437 159836
rect 164923 159900 164989 159901
rect 164923 159836 164924 159900
rect 164988 159836 164989 159900
rect 164923 159835 164989 159836
rect 163635 159628 163701 159629
rect 163635 159564 163636 159628
rect 163700 159564 163701 159628
rect 163635 159563 163701 159564
rect 163451 158540 163517 158541
rect 163451 158476 163452 158540
rect 163516 158476 163517 158540
rect 163451 158475 163517 158476
rect 164374 157861 164434 159835
rect 164926 158677 164986 159835
rect 165294 159765 165354 224163
rect 165478 159765 165538 233139
rect 168235 232524 168301 232525
rect 168235 232460 168236 232524
rect 168300 232460 168301 232524
rect 168235 232459 168301 232460
rect 168051 231844 168117 231845
rect 168051 231780 168052 231844
rect 168116 231780 168117 231844
rect 168051 231779 168117 231780
rect 166763 231300 166829 231301
rect 166763 231236 166764 231300
rect 166828 231236 166829 231300
rect 166763 231235 166829 231236
rect 166579 230076 166645 230077
rect 166579 230012 166580 230076
rect 166644 230012 166645 230076
rect 166579 230011 166645 230012
rect 166395 217972 166461 217973
rect 166395 217908 166396 217972
rect 166460 217908 166461 217972
rect 166395 217907 166461 217908
rect 166211 209676 166277 209677
rect 166211 209612 166212 209676
rect 166276 209612 166277 209676
rect 166211 209611 166277 209612
rect 166027 160444 166093 160445
rect 166027 160380 166028 160444
rect 166092 160380 166093 160444
rect 166027 160379 166093 160380
rect 165291 159764 165357 159765
rect 165291 159700 165292 159764
rect 165356 159700 165357 159764
rect 165291 159699 165357 159700
rect 165475 159764 165541 159765
rect 165475 159700 165476 159764
rect 165540 159700 165541 159764
rect 165475 159699 165541 159700
rect 164923 158676 164989 158677
rect 164923 158612 164924 158676
rect 164988 158612 164989 158676
rect 164923 158611 164989 158612
rect 165294 158541 165354 159699
rect 166030 159629 166090 160379
rect 166214 159765 166274 209611
rect 166398 159901 166458 217907
rect 166582 159901 166642 230011
rect 166766 160037 166826 231235
rect 167867 217836 167933 217837
rect 167867 217772 167868 217836
rect 167932 217772 167933 217836
rect 167867 217771 167933 217772
rect 167683 217564 167749 217565
rect 167683 217500 167684 217564
rect 167748 217500 167749 217564
rect 167683 217499 167749 217500
rect 167131 160716 167197 160717
rect 167131 160652 167132 160716
rect 167196 160652 167197 160716
rect 167131 160651 167197 160652
rect 167134 160173 167194 160651
rect 167315 160580 167381 160581
rect 167315 160516 167316 160580
rect 167380 160516 167381 160580
rect 167315 160515 167381 160516
rect 167131 160172 167197 160173
rect 167131 160108 167132 160172
rect 167196 160108 167197 160172
rect 167131 160107 167197 160108
rect 166763 160036 166829 160037
rect 166763 159972 166764 160036
rect 166828 159972 166829 160036
rect 166763 159971 166829 159972
rect 166395 159900 166461 159901
rect 166395 159836 166396 159900
rect 166460 159836 166461 159900
rect 166395 159835 166461 159836
rect 166579 159900 166645 159901
rect 166579 159836 166580 159900
rect 166644 159836 166645 159900
rect 166579 159835 166645 159836
rect 166211 159764 166277 159765
rect 166211 159700 166212 159764
rect 166276 159700 166277 159764
rect 166211 159699 166277 159700
rect 166027 159628 166093 159629
rect 166027 159564 166028 159628
rect 166092 159564 166093 159628
rect 166027 159563 166093 159564
rect 165843 159084 165909 159085
rect 165843 159020 165844 159084
rect 165908 159020 165909 159084
rect 165843 159019 165909 159020
rect 165291 158540 165357 158541
rect 165291 158476 165292 158540
rect 165356 158476 165357 158540
rect 165291 158475 165357 158476
rect 165659 158540 165725 158541
rect 165659 158476 165660 158540
rect 165724 158476 165725 158540
rect 165659 158475 165725 158476
rect 164371 157860 164437 157861
rect 164371 157796 164372 157860
rect 164436 157796 164437 157860
rect 164371 157795 164437 157796
rect 164371 157316 164437 157317
rect 164371 157252 164372 157316
rect 164436 157252 164437 157316
rect 164371 157251 164437 157252
rect 163267 156500 163333 156501
rect 163267 156436 163268 156500
rect 163332 156436 163333 156500
rect 163267 156435 163333 156436
rect 163083 145620 163149 145621
rect 163083 145556 163084 145620
rect 163148 145556 163149 145620
rect 163083 145555 163149 145556
rect 164374 130389 164434 157251
rect 165662 131749 165722 158475
rect 165846 158133 165906 159019
rect 166766 158677 166826 159971
rect 167318 159901 167378 160515
rect 167315 159900 167381 159901
rect 167315 159836 167316 159900
rect 167380 159836 167381 159900
rect 167315 159835 167381 159836
rect 167686 159765 167746 217499
rect 167870 159901 167930 217771
rect 167867 159900 167933 159901
rect 167867 159836 167868 159900
rect 167932 159836 167933 159900
rect 167867 159835 167933 159836
rect 167683 159764 167749 159765
rect 167683 159700 167684 159764
rect 167748 159700 167749 159764
rect 167683 159699 167749 159700
rect 168054 158677 168114 231779
rect 168238 159629 168298 232459
rect 169339 217428 169405 217429
rect 169339 217364 169340 217428
rect 169404 217364 169405 217428
rect 169339 217363 169405 217364
rect 169155 211988 169221 211989
rect 169155 211924 169156 211988
rect 169220 211924 169221 211988
rect 169155 211923 169221 211924
rect 169158 167010 169218 211923
rect 168974 166950 169218 167010
rect 168974 159901 169034 166950
rect 169155 161804 169221 161805
rect 169155 161740 169156 161804
rect 169220 161740 169221 161804
rect 169155 161739 169221 161740
rect 168971 159900 169037 159901
rect 168971 159836 168972 159900
rect 169036 159836 169037 159900
rect 168971 159835 169037 159836
rect 169158 159765 169218 161739
rect 169342 160037 169402 217363
rect 169339 160036 169405 160037
rect 169339 159972 169340 160036
rect 169404 159972 169405 160036
rect 169339 159971 169405 159972
rect 169526 159765 169586 235451
rect 173755 234020 173821 234021
rect 173755 233956 173756 234020
rect 173820 233956 173821 234020
rect 173755 233955 173821 233956
rect 172283 231572 172349 231573
rect 172283 231508 172284 231572
rect 172348 231508 172349 231572
rect 172283 231507 172349 231508
rect 170627 231164 170693 231165
rect 170627 231100 170628 231164
rect 170692 231100 170693 231164
rect 170627 231099 170693 231100
rect 170075 220420 170141 220421
rect 170075 220356 170076 220420
rect 170140 220356 170141 220420
rect 170075 220355 170141 220356
rect 170078 159901 170138 220355
rect 170443 217700 170509 217701
rect 170443 217636 170444 217700
rect 170508 217636 170509 217700
rect 170443 217635 170509 217636
rect 170259 217292 170325 217293
rect 170259 217228 170260 217292
rect 170324 217228 170325 217292
rect 170259 217227 170325 217228
rect 170075 159900 170141 159901
rect 170075 159836 170076 159900
rect 170140 159836 170141 159900
rect 170075 159835 170141 159836
rect 168603 159764 168669 159765
rect 168603 159700 168604 159764
rect 168668 159700 168669 159764
rect 168603 159699 168669 159700
rect 169155 159764 169221 159765
rect 169155 159700 169156 159764
rect 169220 159700 169221 159764
rect 169155 159699 169221 159700
rect 169523 159764 169589 159765
rect 169523 159700 169524 159764
rect 169588 159700 169589 159764
rect 169523 159699 169589 159700
rect 168235 159628 168301 159629
rect 168235 159564 168236 159628
rect 168300 159564 168301 159628
rect 168235 159563 168301 159564
rect 166763 158676 166829 158677
rect 166763 158612 166764 158676
rect 166828 158612 166829 158676
rect 166763 158611 166829 158612
rect 168051 158676 168117 158677
rect 168051 158612 168052 158676
rect 168116 158612 168117 158676
rect 168051 158611 168117 158612
rect 168238 158405 168298 159563
rect 168606 159357 168666 159699
rect 168603 159356 168669 159357
rect 168603 159292 168604 159356
rect 168668 159292 168669 159356
rect 168603 159291 168669 159292
rect 168606 158949 168666 159291
rect 168603 158948 168669 158949
rect 168603 158884 168604 158948
rect 168668 158884 168669 158948
rect 168603 158883 168669 158884
rect 169526 158677 169586 159699
rect 168419 158676 168485 158677
rect 168419 158612 168420 158676
rect 168484 158612 168485 158676
rect 168419 158611 168485 158612
rect 169523 158676 169589 158677
rect 169523 158612 169524 158676
rect 169588 158612 169589 158676
rect 169523 158611 169589 158612
rect 170075 158676 170141 158677
rect 170075 158612 170076 158676
rect 170140 158612 170141 158676
rect 170075 158611 170141 158612
rect 168235 158404 168301 158405
rect 168235 158340 168236 158404
rect 168300 158340 168301 158404
rect 168235 158339 168301 158340
rect 166947 158268 167013 158269
rect 166947 158204 166948 158268
rect 167012 158204 167013 158268
rect 166947 158203 167013 158204
rect 165843 158132 165909 158133
rect 165843 158068 165844 158132
rect 165908 158068 165909 158132
rect 166950 158130 167010 158203
rect 165843 158067 165909 158068
rect 166766 158070 167010 158130
rect 165659 131748 165725 131749
rect 165659 131684 165660 131748
rect 165724 131684 165725 131748
rect 165659 131683 165725 131684
rect 164371 130388 164437 130389
rect 164371 130324 164372 130388
rect 164436 130324 164437 130388
rect 164371 130323 164437 130324
rect 162899 122092 162965 122093
rect 162899 122028 162900 122092
rect 162964 122028 162965 122092
rect 162899 122027 162965 122028
rect 165846 113797 165906 158067
rect 166766 157725 166826 158070
rect 166763 157724 166829 157725
rect 166763 157660 166764 157724
rect 166828 157660 166829 157724
rect 166763 157659 166829 157660
rect 168235 157724 168301 157725
rect 168235 157660 168236 157724
rect 168300 157660 168301 157724
rect 168235 157659 168301 157660
rect 168238 140589 168298 157659
rect 168422 156909 168482 158611
rect 168971 158268 169037 158269
rect 168971 158204 168972 158268
rect 169036 158204 169037 158268
rect 168971 158203 169037 158204
rect 169891 158268 169957 158269
rect 169891 158204 169892 158268
rect 169956 158204 169957 158268
rect 169891 158203 169957 158204
rect 168603 158132 168669 158133
rect 168603 158068 168604 158132
rect 168668 158068 168669 158132
rect 168603 158067 168669 158068
rect 168419 156908 168485 156909
rect 168419 156844 168420 156908
rect 168484 156844 168485 156908
rect 168419 156843 168485 156844
rect 168235 140588 168301 140589
rect 168235 140524 168236 140588
rect 168300 140524 168301 140588
rect 168235 140523 168301 140524
rect 168238 137325 168298 140523
rect 168235 137324 168301 137325
rect 168235 137260 168236 137324
rect 168300 137260 168301 137324
rect 168235 137259 168301 137260
rect 168422 126309 168482 156843
rect 168606 130525 168666 158067
rect 168974 135965 169034 158203
rect 169707 157588 169773 157589
rect 169707 157524 169708 157588
rect 169772 157524 169773 157588
rect 169707 157523 169773 157524
rect 168971 135964 169037 135965
rect 168971 135900 168972 135964
rect 169036 135900 169037 135964
rect 168971 135899 169037 135900
rect 168603 130524 168669 130525
rect 168603 130460 168604 130524
rect 168668 130460 168669 130524
rect 168603 130459 168669 130460
rect 168419 126308 168485 126309
rect 168419 126244 168420 126308
rect 168484 126244 168485 126308
rect 168419 126243 168485 126244
rect 169710 122229 169770 157523
rect 169894 147525 169954 158203
rect 170078 149837 170138 158611
rect 170262 158133 170322 217227
rect 170446 159762 170506 217635
rect 170630 159901 170690 231099
rect 172099 217156 172165 217157
rect 172099 217092 172100 217156
rect 172164 217092 172165 217156
rect 172099 217091 172165 217092
rect 171915 215932 171981 215933
rect 171915 215868 171916 215932
rect 171980 215868 171981 215932
rect 171915 215867 171981 215868
rect 171179 209540 171245 209541
rect 171179 209476 171180 209540
rect 171244 209476 171245 209540
rect 171179 209475 171245 209476
rect 170995 161940 171061 161941
rect 170995 161876 170996 161940
rect 171060 161876 171061 161940
rect 170995 161875 171061 161876
rect 170627 159900 170693 159901
rect 170627 159836 170628 159900
rect 170692 159898 170693 159900
rect 170692 159838 170874 159898
rect 170692 159836 170693 159838
rect 170627 159835 170693 159836
rect 170627 159764 170693 159765
rect 170627 159762 170628 159764
rect 170446 159702 170628 159762
rect 170627 159700 170628 159702
rect 170692 159700 170693 159764
rect 170627 159699 170693 159700
rect 170443 159628 170509 159629
rect 170443 159564 170444 159628
rect 170508 159564 170509 159628
rect 170443 159563 170509 159564
rect 170259 158132 170325 158133
rect 170259 158068 170260 158132
rect 170324 158068 170325 158132
rect 170259 158067 170325 158068
rect 170446 157317 170506 159563
rect 170630 158269 170690 159699
rect 170627 158268 170693 158269
rect 170627 158204 170628 158268
rect 170692 158204 170693 158268
rect 170627 158203 170693 158204
rect 170814 158133 170874 159838
rect 170998 159765 171058 161875
rect 170995 159764 171061 159765
rect 170995 159700 170996 159764
rect 171060 159700 171061 159764
rect 170995 159699 171061 159700
rect 171182 158810 171242 209475
rect 171918 159901 171978 215867
rect 171915 159900 171981 159901
rect 171915 159836 171916 159900
rect 171980 159836 171981 159900
rect 171915 159835 171981 159836
rect 170998 158750 171242 158810
rect 170998 158405 171058 158750
rect 171918 158677 171978 159835
rect 172102 159765 172162 217091
rect 172286 160037 172346 231507
rect 173571 229940 173637 229941
rect 173571 229876 173572 229940
rect 173636 229876 173637 229940
rect 173571 229875 173637 229876
rect 173387 213620 173453 213621
rect 173387 213556 173388 213620
rect 173452 213556 173453 213620
rect 173387 213555 173453 213556
rect 173203 213348 173269 213349
rect 173203 213284 173204 213348
rect 173268 213284 173269 213348
rect 173203 213283 173269 213284
rect 173206 160037 173266 213283
rect 172283 160036 172349 160037
rect 172283 159972 172284 160036
rect 172348 159972 172349 160036
rect 172283 159971 172349 159972
rect 173203 160036 173269 160037
rect 173203 159972 173204 160036
rect 173268 159972 173269 160036
rect 173203 159971 173269 159972
rect 173390 159901 173450 213555
rect 173574 159901 173634 229875
rect 172835 159900 172901 159901
rect 172835 159836 172836 159900
rect 172900 159836 172901 159900
rect 172835 159835 172901 159836
rect 173387 159900 173453 159901
rect 173387 159836 173388 159900
rect 173452 159836 173453 159900
rect 173387 159835 173453 159836
rect 173571 159900 173637 159901
rect 173571 159836 173572 159900
rect 173636 159836 173637 159900
rect 173571 159835 173637 159836
rect 172099 159764 172165 159765
rect 172099 159700 172100 159764
rect 172164 159700 172165 159764
rect 172099 159699 172165 159700
rect 172651 159628 172717 159629
rect 172651 159564 172652 159628
rect 172716 159564 172717 159628
rect 172651 159563 172717 159564
rect 171547 158676 171613 158677
rect 171547 158612 171548 158676
rect 171612 158612 171613 158676
rect 171547 158611 171613 158612
rect 171915 158676 171981 158677
rect 171915 158612 171916 158676
rect 171980 158612 171981 158676
rect 171915 158611 171981 158612
rect 170995 158404 171061 158405
rect 170995 158340 170996 158404
rect 171060 158340 171061 158404
rect 170995 158339 171061 158340
rect 171179 158404 171245 158405
rect 171179 158340 171180 158404
rect 171244 158340 171245 158404
rect 171179 158339 171245 158340
rect 170811 158132 170877 158133
rect 170811 158068 170812 158132
rect 170876 158068 170877 158132
rect 170811 158067 170877 158068
rect 170443 157316 170509 157317
rect 170443 157252 170444 157316
rect 170508 157252 170509 157316
rect 170443 157251 170509 157252
rect 170075 149836 170141 149837
rect 170075 149772 170076 149836
rect 170140 149772 170141 149836
rect 170075 149771 170141 149772
rect 171182 147661 171242 158339
rect 171179 147660 171245 147661
rect 171179 147596 171180 147660
rect 171244 147596 171245 147660
rect 171179 147595 171245 147596
rect 169891 147524 169957 147525
rect 169891 147460 169892 147524
rect 169956 147460 169957 147524
rect 169891 147459 169957 147460
rect 171550 144533 171610 158611
rect 172654 153210 172714 159563
rect 172470 153150 172714 153210
rect 171731 153100 171797 153101
rect 171731 153036 171732 153100
rect 171796 153036 171797 153100
rect 171731 153035 171797 153036
rect 171547 144532 171613 144533
rect 171547 144468 171548 144532
rect 171612 144468 171613 144532
rect 171547 144467 171613 144468
rect 171734 136101 171794 153035
rect 171731 136100 171797 136101
rect 171731 136036 171732 136100
rect 171796 136036 171797 136100
rect 171731 136035 171797 136036
rect 172470 126445 172530 153150
rect 172838 149973 172898 159835
rect 173758 159765 173818 233955
rect 175043 232932 175109 232933
rect 175043 232868 175044 232932
rect 175108 232868 175109 232932
rect 175043 232867 175109 232868
rect 174859 231436 174925 231437
rect 174859 231372 174860 231436
rect 174924 231372 174925 231436
rect 174859 231371 174925 231372
rect 174675 220284 174741 220285
rect 174675 220220 174676 220284
rect 174740 220220 174741 220284
rect 174675 220219 174741 220220
rect 174491 213212 174557 213213
rect 174491 213148 174492 213212
rect 174556 213148 174557 213212
rect 174491 213147 174557 213148
rect 173019 159764 173085 159765
rect 173019 159700 173020 159764
rect 173084 159700 173085 159764
rect 173019 159699 173085 159700
rect 173387 159764 173453 159765
rect 173387 159700 173388 159764
rect 173452 159700 173453 159764
rect 173387 159699 173453 159700
rect 173755 159764 173821 159765
rect 173755 159700 173756 159764
rect 173820 159700 173821 159764
rect 173755 159699 173821 159700
rect 173022 158949 173082 159699
rect 173019 158948 173085 158949
rect 173019 158884 173020 158948
rect 173084 158884 173085 158948
rect 173019 158883 173085 158884
rect 173390 158269 173450 159699
rect 174494 159629 174554 213147
rect 174678 159765 174738 220219
rect 174862 159901 174922 231371
rect 175046 160037 175106 232867
rect 175043 160036 175109 160037
rect 175043 159972 175044 160036
rect 175108 159972 175109 160036
rect 175043 159971 175109 159972
rect 174859 159900 174925 159901
rect 174859 159836 174860 159900
rect 174924 159836 174925 159900
rect 174859 159835 174925 159836
rect 174675 159764 174741 159765
rect 174675 159700 174676 159764
rect 174740 159700 174741 159764
rect 174675 159699 174741 159700
rect 174491 159628 174557 159629
rect 174491 159564 174492 159628
rect 174556 159564 174557 159628
rect 174491 159563 174557 159564
rect 173571 158676 173637 158677
rect 173571 158612 173572 158676
rect 173636 158612 173637 158676
rect 173571 158611 173637 158612
rect 173387 158268 173453 158269
rect 173387 158204 173388 158268
rect 173452 158204 173453 158268
rect 173387 158203 173453 158204
rect 172835 149972 172901 149973
rect 172835 149908 172836 149972
rect 172900 149908 172901 149972
rect 172835 149907 172901 149908
rect 173574 149565 173634 158611
rect 174494 158269 174554 159563
rect 175782 159493 175842 237899
rect 175966 160717 176026 238171
rect 176515 235244 176581 235245
rect 176515 235180 176516 235244
rect 176580 235180 176581 235244
rect 176515 235179 176581 235180
rect 176147 215116 176213 215117
rect 176147 215052 176148 215116
rect 176212 215052 176213 215116
rect 176147 215051 176213 215052
rect 176150 167010 176210 215051
rect 176150 166950 176394 167010
rect 175963 160716 176029 160717
rect 175963 160652 175964 160716
rect 176028 160652 176029 160716
rect 175963 160651 176029 160652
rect 175779 159492 175845 159493
rect 175779 159428 175780 159492
rect 175844 159428 175845 159492
rect 175779 159427 175845 159428
rect 174675 158676 174741 158677
rect 174675 158612 174676 158676
rect 174740 158612 174741 158676
rect 174675 158611 174741 158612
rect 176147 158676 176213 158677
rect 176147 158612 176148 158676
rect 176212 158612 176213 158676
rect 176147 158611 176213 158612
rect 174491 158268 174557 158269
rect 174491 158204 174492 158268
rect 174556 158204 174557 158268
rect 174491 158203 174557 158204
rect 173755 157316 173821 157317
rect 173755 157252 173756 157316
rect 173820 157252 173821 157316
rect 173755 157251 173821 157252
rect 173571 149564 173637 149565
rect 173571 149500 173572 149564
rect 173636 149500 173637 149564
rect 173571 149499 173637 149500
rect 173574 148477 173634 149499
rect 173571 148476 173637 148477
rect 173571 148412 173572 148476
rect 173636 148412 173637 148476
rect 173571 148411 173637 148412
rect 173758 147389 173818 157251
rect 174678 153781 174738 158611
rect 175043 158404 175109 158405
rect 175043 158340 175044 158404
rect 175108 158340 175109 158404
rect 175043 158339 175109 158340
rect 175963 158404 176029 158405
rect 175963 158340 175964 158404
rect 176028 158340 176029 158404
rect 175963 158339 176029 158340
rect 174675 153780 174741 153781
rect 174675 153716 174676 153780
rect 174740 153716 174741 153780
rect 174675 153715 174741 153716
rect 175046 151830 175106 158339
rect 175966 152965 176026 158339
rect 176150 153101 176210 158611
rect 176334 158133 176394 166950
rect 176518 159901 176578 235179
rect 181483 234428 181549 234429
rect 181483 234364 181484 234428
rect 181548 234364 181549 234428
rect 181483 234363 181549 234364
rect 181299 234292 181365 234293
rect 181299 234228 181300 234292
rect 181364 234228 181365 234292
rect 181299 234227 181365 234228
rect 180563 233884 180629 233885
rect 180563 233820 180564 233884
rect 180628 233820 180629 233884
rect 180563 233819 180629 233820
rect 180379 224364 180445 224365
rect 180379 224300 180380 224364
rect 180444 224300 180445 224364
rect 180379 224299 180445 224300
rect 178907 222868 178973 222869
rect 178907 222804 178908 222868
rect 178972 222804 178973 222868
rect 178907 222803 178973 222804
rect 177619 213756 177685 213757
rect 177619 213692 177620 213756
rect 177684 213692 177685 213756
rect 177619 213691 177685 213692
rect 177622 159901 177682 213691
rect 177803 213076 177869 213077
rect 177803 213012 177804 213076
rect 177868 213012 177869 213076
rect 177803 213011 177869 213012
rect 176515 159900 176581 159901
rect 176515 159836 176516 159900
rect 176580 159836 176581 159900
rect 176515 159835 176581 159836
rect 177619 159900 177685 159901
rect 177619 159836 177620 159900
rect 177684 159836 177685 159900
rect 177619 159835 177685 159836
rect 177806 159765 177866 213011
rect 178910 159901 178970 222803
rect 179091 218652 179157 218653
rect 179091 218588 179092 218652
rect 179156 218588 179157 218652
rect 179091 218587 179157 218588
rect 178907 159900 178973 159901
rect 178907 159836 178908 159900
rect 178972 159836 178973 159900
rect 178907 159835 178973 159836
rect 176883 159764 176949 159765
rect 176883 159700 176884 159764
rect 176948 159700 176949 159764
rect 176883 159699 176949 159700
rect 177803 159764 177869 159765
rect 177803 159700 177804 159764
rect 177868 159700 177869 159764
rect 177803 159699 177869 159700
rect 176886 159357 176946 159699
rect 176883 159356 176949 159357
rect 176883 159292 176884 159356
rect 176948 159292 176949 159356
rect 176883 159291 176949 159292
rect 176515 158812 176581 158813
rect 176515 158748 176516 158812
rect 176580 158748 176581 158812
rect 176515 158747 176581 158748
rect 176331 158132 176397 158133
rect 176331 158068 176332 158132
rect 176396 158068 176397 158132
rect 176331 158067 176397 158068
rect 176147 153100 176213 153101
rect 176147 153036 176148 153100
rect 176212 153036 176213 153100
rect 176147 153035 176213 153036
rect 175963 152964 176029 152965
rect 175963 152900 175964 152964
rect 176028 152900 176029 152964
rect 175963 152899 176029 152900
rect 174494 151770 175106 151830
rect 174494 147525 174554 151770
rect 175966 149157 176026 152899
rect 175963 149156 176029 149157
rect 175963 149092 175964 149156
rect 176028 149092 176029 149156
rect 175963 149091 176029 149092
rect 174491 147524 174557 147525
rect 174491 147460 174492 147524
rect 174556 147460 174557 147524
rect 174491 147459 174557 147460
rect 173755 147388 173821 147389
rect 173755 147324 173756 147388
rect 173820 147324 173821 147388
rect 173755 147323 173821 147324
rect 173758 142170 173818 147323
rect 173022 142110 173818 142170
rect 173022 140045 173082 142110
rect 174494 141405 174554 147459
rect 174491 141404 174557 141405
rect 174491 141340 174492 141404
rect 174556 141340 174557 141404
rect 174491 141339 174557 141340
rect 173019 140044 173085 140045
rect 173019 139980 173020 140044
rect 173084 139980 173085 140044
rect 173019 139979 173085 139980
rect 172467 126444 172533 126445
rect 172467 126380 172468 126444
rect 172532 126380 172533 126444
rect 172467 126379 172533 126380
rect 169707 122228 169773 122229
rect 169707 122164 169708 122228
rect 169772 122164 169773 122228
rect 169707 122163 169773 122164
rect 165843 113796 165909 113797
rect 165843 113732 165844 113796
rect 165908 113732 165909 113796
rect 165843 113731 165909 113732
rect 176518 98701 176578 158747
rect 177619 158676 177685 158677
rect 177619 158612 177620 158676
rect 177684 158612 177685 158676
rect 177619 158611 177685 158612
rect 178723 158676 178789 158677
rect 178723 158612 178724 158676
rect 178788 158612 178789 158676
rect 178723 158611 178789 158612
rect 177435 158132 177501 158133
rect 177435 158068 177436 158132
rect 177500 158068 177501 158132
rect 177435 158067 177501 158068
rect 177251 157996 177317 157997
rect 177251 157932 177252 157996
rect 177316 157932 177317 157996
rect 177251 157931 177317 157932
rect 177254 140861 177314 157931
rect 177438 149837 177498 158067
rect 177435 149836 177501 149837
rect 177435 149772 177436 149836
rect 177500 149772 177501 149836
rect 177435 149771 177501 149772
rect 177251 140860 177317 140861
rect 177251 140796 177252 140860
rect 177316 140796 177317 140860
rect 177251 140795 177317 140796
rect 177438 116517 177498 149771
rect 177622 147253 177682 158611
rect 177987 157860 178053 157861
rect 177987 157796 177988 157860
rect 178052 157796 178053 157860
rect 177987 157795 178053 157796
rect 177990 154053 178050 157795
rect 177987 154052 178053 154053
rect 177987 153988 177988 154052
rect 178052 153988 178053 154052
rect 177987 153987 178053 153988
rect 177619 147252 177685 147253
rect 177619 147188 177620 147252
rect 177684 147188 177685 147252
rect 177619 147187 177685 147188
rect 177435 116516 177501 116517
rect 177435 116452 177436 116516
rect 177500 116452 177501 116516
rect 177435 116451 177501 116452
rect 176515 98700 176581 98701
rect 176515 98636 176516 98700
rect 176580 98636 176581 98700
rect 176515 98635 176581 98636
rect 162715 71092 162781 71093
rect 162715 71028 162716 71092
rect 162780 71028 162781 71092
rect 162715 71027 162781 71028
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 177622 28253 177682 147187
rect 177990 142170 178050 153987
rect 178726 148613 178786 158611
rect 178910 151061 178970 159835
rect 179094 159765 179154 218587
rect 180195 213892 180261 213893
rect 180195 213828 180196 213892
rect 180260 213828 180261 213892
rect 180195 213827 180261 213828
rect 180011 211852 180077 211853
rect 180011 211788 180012 211852
rect 180076 211788 180077 211852
rect 180011 211787 180077 211788
rect 179568 187174 179888 187206
rect 179568 186938 179610 187174
rect 179846 186938 179888 187174
rect 179568 186854 179888 186938
rect 179568 186618 179610 186854
rect 179846 186618 179888 186854
rect 179568 186586 179888 186618
rect 180014 159901 180074 211787
rect 180011 159900 180077 159901
rect 180011 159836 180012 159900
rect 180076 159836 180077 159900
rect 180011 159835 180077 159836
rect 179091 159764 179157 159765
rect 179091 159700 179092 159764
rect 179156 159700 179157 159764
rect 179091 159699 179157 159700
rect 178907 151060 178973 151061
rect 178907 150996 178908 151060
rect 178972 150996 178973 151060
rect 178907 150995 178973 150996
rect 178723 148612 178789 148613
rect 178723 148548 178724 148612
rect 178788 148548 178789 148612
rect 178723 148547 178789 148548
rect 177806 142110 178050 142170
rect 177806 141541 177866 142110
rect 177803 141540 177869 141541
rect 177803 141476 177804 141540
rect 177868 141476 177869 141540
rect 177803 141475 177869 141476
rect 177803 141404 177869 141405
rect 177803 141340 177804 141404
rect 177868 141340 177869 141404
rect 177803 141339 177869 141340
rect 177806 140861 177866 141339
rect 177803 140860 177869 140861
rect 177803 140796 177804 140860
rect 177868 140796 177869 140860
rect 177803 140795 177869 140796
rect 177619 28252 177685 28253
rect 177619 28188 177620 28252
rect 177684 28188 177685 28252
rect 177619 28187 177685 28188
rect 177806 17237 177866 140795
rect 179094 140045 179154 159699
rect 179827 158676 179893 158677
rect 179827 158612 179828 158676
rect 179892 158612 179893 158676
rect 179827 158611 179893 158612
rect 179091 140044 179157 140045
rect 179091 139980 179092 140044
rect 179156 139980 179157 140044
rect 179091 139979 179157 139980
rect 179830 98837 179890 158611
rect 180014 121005 180074 159835
rect 180198 159765 180258 213827
rect 180382 159901 180442 224299
rect 180566 159901 180626 233819
rect 181115 226404 181181 226405
rect 181115 226340 181116 226404
rect 181180 226340 181181 226404
rect 181115 226339 181181 226340
rect 180931 221644 180997 221645
rect 180931 221580 180932 221644
rect 180996 221580 180997 221644
rect 180931 221579 180997 221580
rect 180747 160036 180813 160037
rect 180747 159972 180748 160036
rect 180812 159972 180813 160036
rect 180747 159971 180813 159972
rect 180379 159900 180445 159901
rect 180379 159836 180380 159900
rect 180444 159836 180445 159900
rect 180379 159835 180445 159836
rect 180563 159900 180629 159901
rect 180563 159836 180564 159900
rect 180628 159836 180629 159900
rect 180563 159835 180629 159836
rect 180195 159764 180261 159765
rect 180195 159700 180196 159764
rect 180260 159700 180261 159764
rect 180195 159699 180261 159700
rect 180382 124813 180442 159835
rect 180566 158677 180626 159835
rect 180563 158676 180629 158677
rect 180563 158612 180564 158676
rect 180628 158612 180629 158676
rect 180563 158611 180629 158612
rect 180750 147690 180810 159971
rect 180934 159901 180994 221579
rect 180931 159900 180997 159901
rect 180931 159836 180932 159900
rect 180996 159836 180997 159900
rect 181118 159898 181178 226339
rect 181302 160170 181362 234227
rect 181486 160309 181546 234363
rect 181794 219454 182414 254898
rect 185514 705798 186134 705830
rect 185514 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 186134 705798
rect 185514 705478 186134 705562
rect 185514 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 186134 705478
rect 185514 691174 186134 705242
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 439174 186134 474618
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 367174 186134 402618
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 295174 186134 330618
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185514 259174 186134 294618
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 221514 705798 222134 705830
rect 221514 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 222134 705798
rect 221514 705478 222134 705562
rect 221514 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 222134 705478
rect 221514 691174 222134 705242
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 439174 222134 474618
rect 221514 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 222134 439174
rect 221514 438854 222134 438938
rect 221514 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 222134 438854
rect 221514 403174 222134 438618
rect 221514 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 222134 403174
rect 221514 402854 222134 402938
rect 221514 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 222134 402854
rect 221227 372740 221293 372741
rect 221227 372676 221228 372740
rect 221292 372676 221293 372740
rect 221227 372675 221293 372676
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 215891 292636 215957 292637
rect 215891 292572 215892 292636
rect 215956 292572 215957 292636
rect 215891 292571 215957 292572
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185163 238100 185229 238101
rect 185163 238036 185164 238100
rect 185228 238036 185229 238100
rect 185163 238035 185229 238036
rect 183139 235652 183205 235653
rect 183139 235588 183140 235652
rect 183204 235588 183205 235652
rect 183139 235587 183205 235588
rect 182955 234564 183021 234565
rect 182955 234500 182956 234564
rect 183020 234500 183021 234564
rect 182955 234499 183021 234500
rect 182771 234156 182837 234157
rect 182771 234092 182772 234156
rect 182836 234092 182837 234156
rect 182771 234091 182837 234092
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181483 160308 181549 160309
rect 181483 160244 181484 160308
rect 181548 160244 181549 160308
rect 181483 160243 181549 160244
rect 181302 160110 181546 160170
rect 181299 159900 181365 159901
rect 181299 159898 181300 159900
rect 181118 159838 181300 159898
rect 180931 159835 180997 159836
rect 181299 159836 181300 159838
rect 181364 159836 181365 159900
rect 181299 159835 181365 159836
rect 181486 159765 181546 160110
rect 181483 159764 181549 159765
rect 181483 159700 181484 159764
rect 181548 159700 181549 159764
rect 181483 159699 181549 159700
rect 181115 158676 181181 158677
rect 181115 158612 181116 158676
rect 181180 158612 181181 158676
rect 181115 158611 181181 158612
rect 180566 147630 180810 147690
rect 180379 124812 180445 124813
rect 180379 124748 180380 124812
rect 180444 124748 180445 124812
rect 180379 124747 180445 124748
rect 180011 121004 180077 121005
rect 180011 120940 180012 121004
rect 180076 120940 180077 121004
rect 180011 120939 180077 120940
rect 180566 112570 180626 147630
rect 181118 141949 181178 158611
rect 181483 158132 181549 158133
rect 181483 158068 181484 158132
rect 181548 158068 181549 158132
rect 181483 158067 181549 158068
rect 181486 142085 181546 158067
rect 181794 147454 182414 182898
rect 182587 160036 182653 160037
rect 182587 159972 182588 160036
rect 182652 159972 182653 160036
rect 182587 159971 182653 159972
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181483 142084 181549 142085
rect 181483 142020 181484 142084
rect 181548 142020 181549 142084
rect 181483 142019 181549 142020
rect 181115 141948 181181 141949
rect 181115 141884 181116 141948
rect 181180 141884 181181 141948
rect 181115 141883 181181 141884
rect 181118 122229 181178 141883
rect 181115 122228 181181 122229
rect 181115 122164 181116 122228
rect 181180 122164 181181 122228
rect 181115 122163 181181 122164
rect 180566 112510 180810 112570
rect 180750 112437 180810 112510
rect 180747 112436 180813 112437
rect 180747 112372 180748 112436
rect 180812 112372 180813 112436
rect 180747 112371 180813 112372
rect 179827 98836 179893 98837
rect 179827 98772 179828 98836
rect 179892 98772 179893 98836
rect 179827 98771 179893 98772
rect 181486 95981 181546 142019
rect 181794 111454 182414 146898
rect 182590 127669 182650 159971
rect 182774 159901 182834 234091
rect 182771 159900 182837 159901
rect 182771 159836 182772 159900
rect 182836 159836 182837 159900
rect 182771 159835 182837 159836
rect 182958 159765 183018 234499
rect 183142 160037 183202 235587
rect 183323 234700 183389 234701
rect 183323 234636 183324 234700
rect 183388 234636 183389 234700
rect 183323 234635 183389 234636
rect 183139 160036 183205 160037
rect 183139 159972 183140 160036
rect 183204 159972 183205 160036
rect 183139 159971 183205 159972
rect 183326 159901 183386 234635
rect 184427 233748 184493 233749
rect 184427 233684 184428 233748
rect 184492 233684 184493 233748
rect 184427 233683 184493 233684
rect 184059 209676 184125 209677
rect 184059 209612 184060 209676
rect 184124 209612 184125 209676
rect 184059 209611 184125 209612
rect 183875 209540 183941 209541
rect 183875 209476 183876 209540
rect 183940 209476 183941 209540
rect 183875 209475 183941 209476
rect 183323 159900 183389 159901
rect 183323 159836 183324 159900
rect 183388 159836 183389 159900
rect 183323 159835 183389 159836
rect 182955 159764 183021 159765
rect 182955 159700 182956 159764
rect 183020 159700 183021 159764
rect 182955 159699 183021 159700
rect 183323 159764 183389 159765
rect 183323 159700 183324 159764
rect 183388 159700 183389 159764
rect 183323 159699 183389 159700
rect 182955 158676 183021 158677
rect 182955 158612 182956 158676
rect 183020 158612 183021 158676
rect 182955 158611 183021 158612
rect 183139 158676 183205 158677
rect 183139 158612 183140 158676
rect 183204 158612 183205 158676
rect 183139 158611 183205 158612
rect 182958 130389 183018 158611
rect 183142 141813 183202 158611
rect 183139 141812 183205 141813
rect 183139 141748 183140 141812
rect 183204 141748 183205 141812
rect 183139 141747 183205 141748
rect 182955 130388 183021 130389
rect 182955 130324 182956 130388
rect 183020 130324 183021 130388
rect 182955 130323 183021 130324
rect 182587 127668 182653 127669
rect 182587 127604 182588 127668
rect 182652 127604 182653 127668
rect 182587 127603 182653 127604
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181483 95980 181549 95981
rect 181483 95916 181484 95980
rect 181548 95916 181549 95980
rect 181483 95915 181549 95916
rect 181794 75454 182414 110898
rect 183142 97341 183202 141747
rect 183139 97340 183205 97341
rect 183139 97276 183140 97340
rect 183204 97276 183205 97340
rect 183139 97275 183205 97276
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 177803 17236 177869 17237
rect 177803 17172 177804 17236
rect 177868 17172 177869 17236
rect 177803 17171 177869 17172
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -1306 150134 6618
rect 149514 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 150134 -1306
rect 149514 -1626 150134 -1542
rect 149514 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 150134 -1626
rect 149514 -1894 150134 -1862
rect 181794 3454 182414 38898
rect 183326 32469 183386 159699
rect 183878 159493 183938 209475
rect 184062 159765 184122 209611
rect 184430 159901 184490 233683
rect 184611 213484 184677 213485
rect 184611 213420 184612 213484
rect 184676 213420 184677 213484
rect 184611 213419 184677 213420
rect 184614 160037 184674 213419
rect 184611 160036 184677 160037
rect 184611 159972 184612 160036
rect 184676 159972 184677 160036
rect 184611 159971 184677 159972
rect 184427 159900 184493 159901
rect 184427 159836 184428 159900
rect 184492 159836 184493 159900
rect 184427 159835 184493 159836
rect 184059 159764 184125 159765
rect 184059 159700 184060 159764
rect 184124 159700 184125 159764
rect 184059 159699 184125 159700
rect 183875 159492 183941 159493
rect 183875 159428 183876 159492
rect 183940 159428 183941 159492
rect 183875 159427 183941 159428
rect 183323 32468 183389 32469
rect 183323 32404 183324 32468
rect 183388 32404 183389 32468
rect 183323 32403 183389 32404
rect 183878 26893 183938 159427
rect 184062 94485 184122 159699
rect 184430 108357 184490 159835
rect 184614 109717 184674 159971
rect 185166 159357 185226 238035
rect 185514 223174 186134 258618
rect 186819 238372 186885 238373
rect 186819 238308 186820 238372
rect 186884 238308 186885 238372
rect 186819 238307 186885 238308
rect 185514 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 186134 223174
rect 185514 222854 186134 222938
rect 185514 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 186134 222854
rect 185514 187174 186134 222618
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 185163 159356 185229 159357
rect 185163 159292 185164 159356
rect 185228 159292 185229 159356
rect 185163 159291 185229 159292
rect 184979 158676 185045 158677
rect 184979 158612 184980 158676
rect 185044 158612 185045 158676
rect 184979 158611 185045 158612
rect 185163 158676 185229 158677
rect 185163 158612 185164 158676
rect 185228 158612 185229 158676
rect 185163 158611 185229 158612
rect 184982 140861 185042 158611
rect 185166 142765 185226 158611
rect 185514 151174 186134 186618
rect 186822 160853 186882 238307
rect 190867 233068 190933 233069
rect 190867 233004 190868 233068
rect 190932 233004 190933 233068
rect 190867 233003 190933 233004
rect 190315 226948 190381 226949
rect 190315 226884 190316 226948
rect 190380 226884 190381 226948
rect 190315 226883 190381 226884
rect 188291 209540 188357 209541
rect 188291 209476 188292 209540
rect 188356 209476 188357 209540
rect 188291 209475 188357 209476
rect 186819 160852 186885 160853
rect 186819 160788 186820 160852
rect 186884 160788 186885 160852
rect 186819 160787 186885 160788
rect 188294 159901 188354 209475
rect 190318 159901 190378 226883
rect 190870 160037 190930 233003
rect 193627 232796 193693 232797
rect 193627 232732 193628 232796
rect 193692 232732 193693 232796
rect 193627 232731 193693 232732
rect 191419 232388 191485 232389
rect 191419 232324 191420 232388
rect 191484 232324 191485 232388
rect 191419 232323 191485 232324
rect 191235 214844 191301 214845
rect 191235 214780 191236 214844
rect 191300 214780 191301 214844
rect 191235 214779 191301 214780
rect 191051 209540 191117 209541
rect 191051 209476 191052 209540
rect 191116 209476 191117 209540
rect 191051 209475 191117 209476
rect 190867 160036 190933 160037
rect 190867 159972 190868 160036
rect 190932 159972 190933 160036
rect 190867 159971 190933 159972
rect 188291 159900 188357 159901
rect 188291 159836 188292 159900
rect 188356 159836 188357 159900
rect 188291 159835 188357 159836
rect 190315 159900 190381 159901
rect 190315 159836 190316 159900
rect 190380 159836 190381 159900
rect 190315 159835 190381 159836
rect 188294 159490 188354 159835
rect 188294 159430 188906 159490
rect 186451 158812 186517 158813
rect 186451 158748 186452 158812
rect 186516 158748 186517 158812
rect 186451 158747 186517 158748
rect 186454 157861 186514 158747
rect 187003 158676 187069 158677
rect 187003 158612 187004 158676
rect 187068 158612 187069 158676
rect 187003 158611 187069 158612
rect 187371 158676 187437 158677
rect 187371 158612 187372 158676
rect 187436 158612 187437 158676
rect 187371 158611 187437 158612
rect 187555 158676 187621 158677
rect 187555 158612 187556 158676
rect 187620 158612 187621 158676
rect 187555 158611 187621 158612
rect 188475 158676 188541 158677
rect 188475 158612 188476 158676
rect 188540 158612 188541 158676
rect 188475 158611 188541 158612
rect 188659 158676 188725 158677
rect 188659 158612 188660 158676
rect 188724 158612 188725 158676
rect 188659 158611 188725 158612
rect 186451 157860 186517 157861
rect 186451 157796 186452 157860
rect 186516 157796 186517 157860
rect 186451 157795 186517 157796
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185163 142764 185229 142765
rect 185163 142700 185164 142764
rect 185228 142700 185229 142764
rect 185163 142699 185229 142700
rect 184979 140860 185045 140861
rect 184979 140796 184980 140860
rect 185044 140796 185045 140860
rect 184979 140795 185045 140796
rect 184611 109716 184677 109717
rect 184611 109652 184612 109716
rect 184676 109652 184677 109716
rect 184611 109651 184677 109652
rect 184427 108356 184493 108357
rect 184427 108292 184428 108356
rect 184492 108292 184493 108356
rect 184427 108291 184493 108292
rect 184059 94484 184125 94485
rect 184059 94420 184060 94484
rect 184124 94420 184125 94484
rect 184059 94419 184125 94420
rect 183875 26892 183941 26893
rect 183875 26828 183876 26892
rect 183940 26828 183941 26892
rect 183875 26827 183941 26828
rect 185166 6085 185226 142699
rect 185514 115174 186134 150618
rect 187006 144669 187066 158611
rect 187187 158132 187253 158133
rect 187187 158068 187188 158132
rect 187252 158068 187253 158132
rect 187187 158067 187253 158068
rect 187003 144668 187069 144669
rect 187003 144604 187004 144668
rect 187068 144604 187069 144668
rect 187003 144603 187069 144604
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 187006 106997 187066 144603
rect 187190 143173 187250 158067
rect 187187 143172 187253 143173
rect 187187 143108 187188 143172
rect 187252 143108 187253 143172
rect 187187 143107 187253 143108
rect 187003 106996 187069 106997
rect 187003 106932 187004 106996
rect 187068 106932 187069 106996
rect 187003 106931 187069 106932
rect 187190 100197 187250 143107
rect 187374 143037 187434 158611
rect 187371 143036 187437 143037
rect 187371 142972 187372 143036
rect 187436 142972 187437 143036
rect 187371 142971 187437 142972
rect 187187 100196 187253 100197
rect 187187 100132 187188 100196
rect 187252 100132 187253 100196
rect 187187 100131 187253 100132
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 187374 69597 187434 142971
rect 187558 142629 187618 158611
rect 188291 157316 188357 157317
rect 188291 157252 188292 157316
rect 188356 157252 188357 157316
rect 188291 157251 188357 157252
rect 187555 142628 187621 142629
rect 187555 142564 187556 142628
rect 187620 142564 187621 142628
rect 187555 142563 187621 142564
rect 187371 69596 187437 69597
rect 187371 69532 187372 69596
rect 187436 69532 187437 69596
rect 187371 69531 187437 69532
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 187558 13021 187618 142563
rect 188294 72453 188354 157251
rect 188478 141677 188538 158611
rect 188662 142901 188722 158611
rect 188659 142900 188725 142901
rect 188659 142836 188660 142900
rect 188724 142836 188725 142900
rect 188659 142835 188725 142836
rect 188475 141676 188541 141677
rect 188475 141612 188476 141676
rect 188540 141612 188541 141676
rect 188475 141611 188541 141612
rect 188291 72452 188357 72453
rect 188291 72388 188292 72452
rect 188356 72388 188357 72452
rect 188291 72387 188357 72388
rect 187555 13020 187621 13021
rect 187555 12956 187556 13020
rect 187620 12956 187621 13020
rect 187555 12955 187621 12956
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 188478 6901 188538 141611
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 188475 6900 188541 6901
rect 188475 6836 188476 6900
rect 188540 6836 188541 6900
rect 188475 6835 188541 6836
rect 188662 6629 188722 142835
rect 188846 6765 188906 159430
rect 189763 158676 189829 158677
rect 189763 158612 189764 158676
rect 189828 158612 189829 158676
rect 189763 158611 189829 158612
rect 189947 158676 190013 158677
rect 189947 158612 189948 158676
rect 190012 158612 190013 158676
rect 189947 158611 190013 158612
rect 190131 158676 190197 158677
rect 190131 158612 190132 158676
rect 190196 158612 190197 158676
rect 190131 158611 190197 158612
rect 189766 143445 189826 158611
rect 189763 143444 189829 143445
rect 189763 143380 189764 143444
rect 189828 143380 189829 143444
rect 189763 143379 189829 143380
rect 189766 113797 189826 143379
rect 189950 143309 190010 158611
rect 189947 143308 190013 143309
rect 189947 143244 189948 143308
rect 190012 143244 190013 143308
rect 189947 143243 190013 143244
rect 189763 113796 189829 113797
rect 189763 113732 189764 113796
rect 189828 113732 189829 113796
rect 189763 113731 189829 113732
rect 189950 64157 190010 143243
rect 190134 138821 190194 158611
rect 190131 138820 190197 138821
rect 190131 138756 190132 138820
rect 190196 138756 190197 138820
rect 190131 138755 190197 138756
rect 189947 64156 190013 64157
rect 189947 64092 189948 64156
rect 190012 64092 190013 64156
rect 189947 64091 190013 64092
rect 190134 9485 190194 138755
rect 190131 9484 190197 9485
rect 190131 9420 190132 9484
rect 190196 9420 190197 9484
rect 190131 9419 190197 9420
rect 188843 6764 188909 6765
rect 188843 6700 188844 6764
rect 188908 6700 188909 6764
rect 188843 6699 188909 6700
rect 185163 6084 185229 6085
rect 185163 6020 185164 6084
rect 185228 6020 185229 6084
rect 185163 6019 185229 6020
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 -1306 186134 6618
rect 188659 6628 188725 6629
rect 188659 6564 188660 6628
rect 188724 6564 188725 6628
rect 188659 6563 188725 6564
rect 190318 3773 190378 159835
rect 190870 58581 190930 159971
rect 191054 159901 191114 209475
rect 191051 159900 191117 159901
rect 191051 159836 191052 159900
rect 191116 159836 191117 159900
rect 191051 159835 191117 159836
rect 191054 102917 191114 159835
rect 191238 159493 191298 214779
rect 191422 159765 191482 232323
rect 192707 232252 192773 232253
rect 192707 232188 192708 232252
rect 192772 232188 192773 232252
rect 192707 232187 192773 232188
rect 192339 209540 192405 209541
rect 192339 209476 192340 209540
rect 192404 209476 192405 209540
rect 192339 209475 192405 209476
rect 192342 159901 192402 209475
rect 192339 159900 192405 159901
rect 192339 159836 192340 159900
rect 192404 159836 192405 159900
rect 192339 159835 192405 159836
rect 192710 159765 192770 232187
rect 192891 214572 192957 214573
rect 192891 214508 192892 214572
rect 192956 214508 192957 214572
rect 192891 214507 192957 214508
rect 192894 159901 192954 214507
rect 193630 171150 193690 232731
rect 195835 214980 195901 214981
rect 195835 214916 195836 214980
rect 195900 214916 195901 214980
rect 195835 214915 195901 214916
rect 195651 214708 195717 214709
rect 195651 214644 195652 214708
rect 195716 214644 195717 214708
rect 195651 214643 195717 214644
rect 193995 209540 194061 209541
rect 193995 209476 193996 209540
rect 194060 209476 194061 209540
rect 193995 209475 194061 209476
rect 195467 209540 195533 209541
rect 195467 209476 195468 209540
rect 195532 209476 195533 209540
rect 195467 209475 195533 209476
rect 193998 171150 194058 209475
rect 194928 183454 195248 183486
rect 194928 183218 194970 183454
rect 195206 183218 195248 183454
rect 194928 183134 195248 183218
rect 194928 182898 194970 183134
rect 195206 182898 195248 183134
rect 194928 182866 195248 182898
rect 193630 171090 193874 171150
rect 193998 171090 194242 171150
rect 193814 159901 193874 171090
rect 194182 159901 194242 171090
rect 195470 159901 195530 209475
rect 195654 159901 195714 214643
rect 192891 159900 192957 159901
rect 192891 159836 192892 159900
rect 192956 159836 192957 159900
rect 192891 159835 192957 159836
rect 193811 159900 193877 159901
rect 193811 159836 193812 159900
rect 193876 159836 193877 159900
rect 193811 159835 193877 159836
rect 194179 159900 194245 159901
rect 194179 159836 194180 159900
rect 194244 159836 194245 159900
rect 194179 159835 194245 159836
rect 195099 159900 195165 159901
rect 195099 159836 195100 159900
rect 195164 159836 195165 159900
rect 195099 159835 195165 159836
rect 195467 159900 195533 159901
rect 195467 159836 195468 159900
rect 195532 159836 195533 159900
rect 195467 159835 195533 159836
rect 195651 159900 195717 159901
rect 195651 159836 195652 159900
rect 195716 159836 195717 159900
rect 195651 159835 195717 159836
rect 191419 159764 191485 159765
rect 191419 159700 191420 159764
rect 191484 159700 191485 159764
rect 191419 159699 191485 159700
rect 192707 159764 192773 159765
rect 192707 159700 192708 159764
rect 192772 159700 192773 159764
rect 192707 159699 192773 159700
rect 191235 159492 191301 159493
rect 191235 159428 191236 159492
rect 191300 159428 191301 159492
rect 191235 159427 191301 159428
rect 191235 158676 191301 158677
rect 191235 158612 191236 158676
rect 191300 158612 191301 158676
rect 191235 158611 191301 158612
rect 191238 138957 191298 158611
rect 191235 138956 191301 138957
rect 191235 138892 191236 138956
rect 191300 138892 191301 138956
rect 191235 138891 191301 138892
rect 191051 102916 191117 102917
rect 191051 102852 191052 102916
rect 191116 102852 191117 102916
rect 191051 102851 191117 102852
rect 191238 62797 191298 138891
rect 191235 62796 191301 62797
rect 191235 62732 191236 62796
rect 191300 62732 191301 62796
rect 191235 62731 191301 62732
rect 191422 61437 191482 159699
rect 192894 159490 192954 159835
rect 192526 159430 192954 159490
rect 192339 157588 192405 157589
rect 192339 157524 192340 157588
rect 192404 157524 192405 157588
rect 192339 157523 192405 157524
rect 192342 157317 192402 157523
rect 192339 157316 192405 157317
rect 192339 157252 192340 157316
rect 192404 157252 192405 157316
rect 192339 157251 192405 157252
rect 191419 61436 191485 61437
rect 191419 61372 191420 61436
rect 191484 61372 191485 61436
rect 191419 61371 191485 61372
rect 190867 58580 190933 58581
rect 190867 58516 190868 58580
rect 190932 58516 190933 58580
rect 190867 58515 190933 58516
rect 192526 6357 192586 159430
rect 192707 158676 192773 158677
rect 192707 158612 192708 158676
rect 192772 158612 192773 158676
rect 192707 158611 192773 158612
rect 192891 158676 192957 158677
rect 192891 158612 192892 158676
rect 192956 158612 192957 158676
rect 192891 158611 192957 158612
rect 192710 138549 192770 158611
rect 192894 141541 192954 158611
rect 192891 141540 192957 141541
rect 192891 141476 192892 141540
rect 192956 141476 192957 141540
rect 192891 141475 192957 141476
rect 192707 138548 192773 138549
rect 192707 138484 192708 138548
rect 192772 138484 192773 138548
rect 192707 138483 192773 138484
rect 192710 6493 192770 138483
rect 192707 6492 192773 6493
rect 192707 6428 192708 6492
rect 192772 6428 192773 6492
rect 192707 6427 192773 6428
rect 192523 6356 192589 6357
rect 192523 6292 192524 6356
rect 192588 6292 192589 6356
rect 192523 6291 192589 6292
rect 192894 6221 192954 141475
rect 193814 82109 193874 159835
rect 193995 158676 194061 158677
rect 193995 158612 193996 158676
rect 194060 158612 194061 158676
rect 193995 158611 194061 158612
rect 193998 138685 194058 158611
rect 193995 138684 194061 138685
rect 193995 138620 193996 138684
rect 194060 138620 194061 138684
rect 193995 138619 194061 138620
rect 193811 82108 193877 82109
rect 193811 82044 193812 82108
rect 193876 82044 193877 82108
rect 193811 82043 193877 82044
rect 193998 54501 194058 138619
rect 193995 54500 194061 54501
rect 193995 54436 193996 54500
rect 194060 54436 194061 54500
rect 193995 54435 194061 54436
rect 194182 53141 194242 159835
rect 194363 158132 194429 158133
rect 194363 158068 194364 158132
rect 194428 158068 194429 158132
rect 194363 158067 194429 158068
rect 194366 139229 194426 158067
rect 194363 139228 194429 139229
rect 194363 139164 194364 139228
rect 194428 139164 194429 139228
rect 194363 139163 194429 139164
rect 194179 53140 194245 53141
rect 194179 53076 194180 53140
rect 194244 53076 194245 53140
rect 194179 53075 194245 53076
rect 194366 21317 194426 139163
rect 194363 21316 194429 21317
rect 194363 21252 194364 21316
rect 194428 21252 194429 21316
rect 194363 21251 194429 21252
rect 195102 9213 195162 159835
rect 195283 158676 195349 158677
rect 195283 158612 195284 158676
rect 195348 158612 195349 158676
rect 195283 158611 195349 158612
rect 195286 155413 195346 158611
rect 195467 158132 195533 158133
rect 195467 158068 195468 158132
rect 195532 158068 195533 158132
rect 195467 158067 195533 158068
rect 195283 155412 195349 155413
rect 195283 155348 195284 155412
rect 195348 155348 195349 155412
rect 195283 155347 195349 155348
rect 195286 120869 195346 155347
rect 195470 139093 195530 158067
rect 195467 139092 195533 139093
rect 195467 139028 195468 139092
rect 195532 139028 195533 139092
rect 195467 139027 195533 139028
rect 195283 120868 195349 120869
rect 195283 120804 195284 120868
rect 195348 120804 195349 120868
rect 195283 120803 195349 120804
rect 195470 9349 195530 139027
rect 195654 14517 195714 159835
rect 195838 159765 195898 214915
rect 215894 212125 215954 292571
rect 217794 291454 218414 326898
rect 221043 292228 221109 292229
rect 221043 292164 221044 292228
rect 221108 292164 221109 292228
rect 221043 292163 221109 292164
rect 218651 292092 218717 292093
rect 218651 292028 218652 292092
rect 218716 292028 218717 292092
rect 218651 292027 218717 292028
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 218654 243541 218714 292027
rect 220123 291548 220189 291549
rect 220123 291484 220124 291548
rect 220188 291484 220189 291548
rect 220123 291483 220189 291484
rect 220126 276725 220186 291483
rect 220307 291412 220373 291413
rect 220307 291348 220308 291412
rect 220372 291348 220373 291412
rect 220307 291347 220373 291348
rect 220310 278085 220370 291347
rect 221046 286381 221106 292163
rect 221230 291277 221290 372675
rect 221514 367174 222134 402618
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 331174 222134 366618
rect 221514 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 222134 331174
rect 221514 330854 222134 330938
rect 221514 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 222134 330854
rect 221514 295174 222134 330618
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 247539 318340 247605 318341
rect 247539 318276 247540 318340
rect 247604 318276 247605 318340
rect 247539 318275 247605 318276
rect 237971 318068 238037 318069
rect 237971 318004 237972 318068
rect 238036 318004 238037 318068
rect 237971 318003 238037 318004
rect 223435 316980 223501 316981
rect 223435 316916 223436 316980
rect 223500 316916 223501 316980
rect 223435 316915 223501 316916
rect 223251 314124 223317 314125
rect 223251 314060 223252 314124
rect 223316 314060 223317 314124
rect 223251 314059 223317 314060
rect 222699 306916 222765 306917
rect 222699 306852 222700 306916
rect 222764 306852 222765 306916
rect 222699 306851 222765 306852
rect 221514 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 222134 295174
rect 221514 294854 222134 294938
rect 221514 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 222134 294854
rect 221227 291276 221293 291277
rect 221227 291212 221228 291276
rect 221292 291212 221293 291276
rect 221227 291211 221293 291212
rect 221043 286380 221109 286381
rect 221043 286316 221044 286380
rect 221108 286316 221109 286380
rect 221043 286315 221109 286316
rect 220307 278084 220373 278085
rect 220307 278020 220308 278084
rect 220372 278020 220373 278084
rect 220307 278019 220373 278020
rect 220123 276724 220189 276725
rect 220123 276660 220124 276724
rect 220188 276660 220189 276724
rect 220123 276659 220189 276660
rect 221230 275229 221290 291211
rect 221227 275228 221293 275229
rect 221227 275164 221228 275228
rect 221292 275164 221293 275228
rect 221227 275163 221293 275164
rect 221514 259174 222134 294618
rect 221514 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 222134 259174
rect 221514 258854 222134 258938
rect 221514 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 222134 258854
rect 218651 243540 218717 243541
rect 218651 243476 218652 243540
rect 218716 243476 218717 243540
rect 218651 243475 218717 243476
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 215891 212124 215957 212125
rect 215891 212060 215892 212124
rect 215956 212060 215957 212124
rect 215891 212059 215957 212060
rect 203379 211172 203445 211173
rect 203379 211108 203380 211172
rect 203444 211108 203445 211172
rect 203379 211107 203445 211108
rect 196755 209676 196821 209677
rect 196755 209612 196756 209676
rect 196820 209612 196821 209676
rect 196755 209611 196821 209612
rect 197859 209676 197925 209677
rect 197859 209612 197860 209676
rect 197924 209612 197925 209676
rect 197859 209611 197925 209612
rect 199331 209676 199397 209677
rect 199331 209612 199332 209676
rect 199396 209612 199397 209676
rect 199331 209611 199397 209612
rect 199699 209676 199765 209677
rect 199699 209612 199700 209676
rect 199764 209612 199765 209676
rect 199699 209611 199765 209612
rect 196387 209540 196453 209541
rect 196387 209476 196388 209540
rect 196452 209476 196453 209540
rect 196387 209475 196453 209476
rect 196390 160037 196450 209475
rect 196571 209404 196637 209405
rect 196571 209340 196572 209404
rect 196636 209340 196637 209404
rect 196571 209339 196637 209340
rect 196387 160036 196453 160037
rect 196387 159972 196388 160036
rect 196452 159972 196453 160036
rect 196387 159971 196453 159972
rect 195835 159764 195901 159765
rect 195835 159700 195836 159764
rect 195900 159700 195901 159764
rect 195835 159699 195901 159700
rect 195838 158677 195898 159699
rect 195835 158676 195901 158677
rect 195835 158612 195836 158676
rect 195900 158612 195901 158676
rect 195835 158611 195901 158612
rect 196203 158676 196269 158677
rect 196203 158612 196204 158676
rect 196268 158612 196269 158676
rect 196203 158611 196269 158612
rect 196206 144397 196266 158611
rect 196390 158133 196450 159971
rect 196574 159901 196634 209339
rect 196758 171150 196818 209611
rect 197862 171150 197922 209611
rect 198595 207636 198661 207637
rect 198595 207572 198596 207636
rect 198660 207572 198661 207636
rect 198595 207571 198661 207572
rect 196758 171090 197002 171150
rect 197862 171090 198474 171150
rect 196571 159900 196637 159901
rect 196571 159836 196572 159900
rect 196636 159836 196637 159900
rect 196571 159835 196637 159836
rect 196387 158132 196453 158133
rect 196387 158068 196388 158132
rect 196452 158068 196453 158132
rect 196387 158067 196453 158068
rect 196203 144396 196269 144397
rect 196203 144332 196204 144396
rect 196268 144332 196269 144396
rect 196203 144331 196269 144332
rect 195651 14516 195717 14517
rect 195651 14452 195652 14516
rect 195716 14452 195717 14516
rect 195651 14451 195717 14452
rect 195467 9348 195533 9349
rect 195467 9284 195468 9348
rect 195532 9284 195533 9348
rect 195467 9283 195533 9284
rect 195099 9212 195165 9213
rect 195099 9148 195100 9212
rect 195164 9148 195165 9212
rect 195099 9147 195165 9148
rect 196574 9077 196634 159835
rect 196942 159765 197002 171090
rect 197859 161260 197925 161261
rect 197859 161196 197860 161260
rect 197924 161196 197925 161260
rect 197859 161195 197925 161196
rect 197862 160173 197922 161195
rect 197859 160172 197925 160173
rect 197859 160108 197860 160172
rect 197924 160108 197925 160172
rect 197859 160107 197925 160108
rect 198414 159901 198474 171090
rect 198411 159900 198477 159901
rect 198411 159836 198412 159900
rect 198476 159836 198477 159900
rect 198411 159835 198477 159836
rect 196939 159764 197005 159765
rect 196939 159700 196940 159764
rect 197004 159700 197005 159764
rect 196939 159699 197005 159700
rect 196755 158676 196821 158677
rect 196755 158612 196756 158676
rect 196820 158612 196821 158676
rect 196755 158611 196821 158612
rect 196758 152285 196818 158611
rect 196755 152284 196821 152285
rect 196755 152220 196756 152284
rect 196820 152220 196821 152284
rect 196755 152219 196821 152220
rect 196758 118013 196818 152219
rect 196755 118012 196821 118013
rect 196755 117948 196756 118012
rect 196820 117948 196821 118012
rect 196755 117947 196821 117948
rect 196571 9076 196637 9077
rect 196571 9012 196572 9076
rect 196636 9012 196637 9076
rect 196571 9011 196637 9012
rect 196942 8941 197002 159699
rect 198227 158676 198293 158677
rect 198227 158612 198228 158676
rect 198292 158612 198293 158676
rect 198227 158611 198293 158612
rect 198043 158404 198109 158405
rect 198043 158340 198044 158404
rect 198108 158340 198109 158404
rect 198043 158339 198109 158340
rect 198046 152421 198106 158339
rect 198043 152420 198109 152421
rect 198043 152356 198044 152420
rect 198108 152356 198109 152420
rect 198043 152355 198109 152356
rect 198046 116517 198106 152355
rect 198230 140725 198290 158611
rect 198227 140724 198293 140725
rect 198227 140660 198228 140724
rect 198292 140660 198293 140724
rect 198227 140659 198293 140660
rect 198043 116516 198109 116517
rect 198043 116452 198044 116516
rect 198108 116452 198109 116516
rect 198043 116451 198109 116452
rect 198230 76533 198290 140659
rect 198227 76532 198293 76533
rect 198227 76468 198228 76532
rect 198292 76468 198293 76532
rect 198227 76467 198293 76468
rect 196939 8940 197005 8941
rect 196939 8876 196940 8940
rect 197004 8876 197005 8940
rect 196939 8875 197005 8876
rect 192891 6220 192957 6221
rect 192891 6156 192892 6220
rect 192956 6156 192957 6220
rect 192891 6155 192957 6156
rect 190315 3772 190381 3773
rect 190315 3708 190316 3772
rect 190380 3708 190381 3772
rect 190315 3707 190381 3708
rect 198414 3501 198474 159835
rect 198598 159765 198658 207571
rect 199334 159901 199394 209611
rect 199515 209540 199581 209541
rect 199515 209476 199516 209540
rect 199580 209476 199581 209540
rect 199515 209475 199581 209476
rect 199518 160037 199578 209475
rect 199702 160173 199762 209611
rect 203382 201381 203442 211107
rect 203379 201380 203445 201381
rect 203379 201316 203380 201380
rect 203444 201316 203445 201380
rect 203379 201315 203445 201316
rect 205955 191044 206021 191045
rect 205955 190980 205956 191044
rect 206020 190980 206021 191044
rect 205955 190979 206021 190980
rect 204115 180028 204181 180029
rect 204115 179964 204116 180028
rect 204180 179964 204181 180028
rect 204115 179963 204181 179964
rect 203931 165068 203997 165069
rect 203931 165004 203932 165068
rect 203996 165004 203997 165068
rect 203931 165003 203997 165004
rect 203563 163572 203629 163573
rect 203563 163508 203564 163572
rect 203628 163508 203629 163572
rect 203563 163507 203629 163508
rect 203195 162076 203261 162077
rect 203195 162012 203196 162076
rect 203260 162012 203261 162076
rect 203195 162011 203261 162012
rect 201355 161940 201421 161941
rect 201355 161876 201356 161940
rect 201420 161876 201421 161940
rect 201355 161875 201421 161876
rect 199699 160172 199765 160173
rect 199699 160108 199700 160172
rect 199764 160108 199765 160172
rect 199699 160107 199765 160108
rect 199515 160036 199581 160037
rect 199515 159972 199516 160036
rect 199580 159972 199581 160036
rect 199515 159971 199581 159972
rect 201358 159901 201418 161875
rect 202827 160580 202893 160581
rect 202827 160516 202828 160580
rect 202892 160516 202893 160580
rect 202827 160515 202893 160516
rect 199331 159900 199397 159901
rect 199331 159836 199332 159900
rect 199396 159898 199397 159900
rect 201355 159900 201421 159901
rect 201355 159898 201356 159900
rect 199396 159838 199762 159898
rect 199396 159836 199397 159838
rect 199331 159835 199397 159836
rect 198595 159764 198661 159765
rect 198595 159700 198596 159764
rect 198660 159700 198661 159764
rect 198595 159699 198661 159700
rect 198598 3637 198658 159699
rect 199331 158676 199397 158677
rect 199331 158612 199332 158676
rect 199396 158612 199397 158676
rect 199331 158611 199397 158612
rect 199334 152965 199394 158611
rect 199515 158404 199581 158405
rect 199515 158340 199516 158404
rect 199580 158340 199581 158404
rect 199515 158339 199581 158340
rect 199331 152964 199397 152965
rect 199331 152900 199332 152964
rect 199396 152900 199397 152964
rect 199331 152899 199397 152900
rect 199334 152557 199394 152899
rect 199331 152556 199397 152557
rect 199331 152492 199332 152556
rect 199396 152492 199397 152556
rect 199331 152491 199397 152492
rect 199518 143989 199578 158339
rect 199702 154597 199762 159838
rect 200806 159838 201356 159898
rect 199883 158676 199949 158677
rect 199883 158612 199884 158676
rect 199948 158612 199949 158676
rect 199883 158611 199949 158612
rect 200619 158676 200685 158677
rect 200619 158612 200620 158676
rect 200684 158612 200685 158676
rect 200619 158611 200685 158612
rect 199886 157181 199946 158611
rect 199883 157180 199949 157181
rect 199883 157116 199884 157180
rect 199948 157116 199949 157180
rect 199883 157115 199949 157116
rect 199699 154596 199765 154597
rect 199699 154532 199700 154596
rect 199764 154532 199765 154596
rect 199699 154531 199765 154532
rect 199699 152556 199765 152557
rect 199699 152492 199700 152556
rect 199764 152492 199765 152556
rect 199699 152491 199765 152492
rect 199515 143988 199581 143989
rect 199515 143924 199516 143988
rect 199580 143924 199581 143988
rect 199515 143923 199581 143924
rect 199702 115157 199762 152491
rect 200622 144397 200682 158611
rect 200806 157453 200866 159838
rect 201355 159836 201356 159838
rect 201420 159836 201421 159900
rect 201355 159835 201421 159836
rect 201355 159084 201421 159085
rect 201355 159020 201356 159084
rect 201420 159020 201421 159084
rect 201355 159019 201421 159020
rect 200987 158676 201053 158677
rect 200987 158612 200988 158676
rect 201052 158612 201053 158676
rect 200987 158611 201053 158612
rect 200803 157452 200869 157453
rect 200803 157388 200804 157452
rect 200868 157388 200869 157452
rect 200803 157387 200869 157388
rect 200990 154189 201050 158611
rect 201358 158405 201418 159019
rect 202643 158676 202709 158677
rect 202643 158612 202644 158676
rect 202708 158612 202709 158676
rect 202643 158611 202709 158612
rect 201171 158404 201237 158405
rect 201171 158340 201172 158404
rect 201236 158340 201237 158404
rect 201171 158339 201237 158340
rect 201355 158404 201421 158405
rect 201355 158340 201356 158404
rect 201420 158340 201421 158404
rect 201355 158339 201421 158340
rect 202459 158404 202525 158405
rect 202459 158340 202460 158404
rect 202524 158340 202525 158404
rect 202459 158339 202525 158340
rect 200987 154188 201053 154189
rect 200987 154124 200988 154188
rect 201052 154124 201053 154188
rect 200987 154123 201053 154124
rect 200619 144396 200685 144397
rect 200619 144332 200620 144396
rect 200684 144332 200685 144396
rect 200619 144331 200685 144332
rect 199883 143988 199949 143989
rect 199883 143924 199884 143988
rect 199948 143924 199949 143988
rect 199883 143923 199949 143924
rect 199699 115156 199765 115157
rect 199699 115092 199700 115156
rect 199764 115092 199765 115156
rect 199699 115091 199765 115092
rect 198595 3636 198661 3637
rect 198595 3572 198596 3636
rect 198660 3572 198661 3636
rect 198595 3571 198661 3572
rect 198411 3500 198477 3501
rect 198411 3436 198412 3500
rect 198476 3436 198477 3500
rect 198411 3435 198477 3436
rect 199886 3365 199946 143923
rect 200622 142170 200682 144331
rect 201174 143853 201234 158339
rect 201355 157996 201421 157997
rect 201355 157932 201356 157996
rect 201420 157932 201421 157996
rect 201355 157931 201421 157932
rect 202091 157996 202157 157997
rect 202091 157932 202092 157996
rect 202156 157932 202157 157996
rect 202091 157931 202157 157932
rect 201358 146165 201418 157931
rect 201355 146164 201421 146165
rect 201355 146100 201356 146164
rect 201420 146100 201421 146164
rect 201355 146099 201421 146100
rect 201171 143852 201237 143853
rect 201171 143788 201172 143852
rect 201236 143788 201237 143852
rect 201171 143787 201237 143788
rect 200622 142110 201050 142170
rect 200990 111077 201050 142110
rect 200987 111076 201053 111077
rect 200987 111012 200988 111076
rect 201052 111012 201053 111076
rect 200987 111011 201053 111012
rect 201174 106861 201234 143787
rect 201171 106860 201237 106861
rect 201171 106796 201172 106860
rect 201236 106796 201237 106860
rect 201171 106795 201237 106796
rect 201358 39269 201418 146099
rect 202094 144397 202154 157931
rect 202275 156092 202341 156093
rect 202275 156028 202276 156092
rect 202340 156028 202341 156092
rect 202275 156027 202341 156028
rect 202091 144396 202157 144397
rect 202091 144332 202092 144396
rect 202156 144332 202157 144396
rect 202091 144331 202157 144332
rect 202278 144125 202338 156027
rect 202462 145893 202522 158339
rect 202646 146301 202706 158611
rect 202830 157725 202890 160515
rect 203198 159765 203258 162011
rect 203379 160852 203445 160853
rect 203379 160788 203380 160852
rect 203444 160788 203445 160852
rect 203379 160787 203445 160788
rect 203382 159765 203442 160787
rect 203566 159901 203626 163507
rect 203563 159900 203629 159901
rect 203563 159836 203564 159900
rect 203628 159836 203629 159900
rect 203563 159835 203629 159836
rect 203195 159764 203261 159765
rect 203195 159700 203196 159764
rect 203260 159700 203261 159764
rect 203195 159699 203261 159700
rect 203379 159764 203445 159765
rect 203379 159700 203380 159764
rect 203444 159700 203445 159764
rect 203379 159699 203445 159700
rect 202827 157724 202893 157725
rect 202827 157660 202828 157724
rect 202892 157660 202893 157724
rect 202827 157659 202893 157660
rect 203566 157350 203626 159835
rect 203934 159765 203994 165003
rect 204118 159901 204178 179963
rect 205403 177308 205469 177309
rect 205403 177244 205404 177308
rect 205468 177244 205469 177308
rect 205403 177243 205469 177244
rect 205219 169012 205285 169013
rect 205219 168948 205220 169012
rect 205284 168948 205285 169012
rect 205219 168947 205285 168948
rect 205222 167010 205282 168947
rect 205038 166950 205282 167010
rect 204667 166020 204733 166021
rect 204667 165956 204668 166020
rect 204732 165956 204733 166020
rect 204667 165955 204733 165956
rect 204115 159900 204181 159901
rect 204115 159836 204116 159900
rect 204180 159836 204181 159900
rect 204115 159835 204181 159836
rect 203931 159764 203997 159765
rect 203931 159700 203932 159764
rect 203996 159700 203997 159764
rect 203931 159699 203997 159700
rect 203747 158676 203813 158677
rect 203747 158612 203748 158676
rect 203812 158612 203813 158676
rect 203747 158611 203813 158612
rect 203931 158676 203997 158677
rect 203931 158612 203932 158676
rect 203996 158612 203997 158676
rect 203931 158611 203997 158612
rect 203198 157290 203626 157350
rect 202643 146300 202709 146301
rect 202643 146236 202644 146300
rect 202708 146236 202709 146300
rect 202643 146235 202709 146236
rect 202459 145892 202525 145893
rect 202459 145828 202460 145892
rect 202524 145828 202525 145892
rect 202459 145827 202525 145828
rect 202275 144124 202341 144125
rect 202275 144060 202276 144124
rect 202340 144060 202341 144124
rect 202275 144059 202341 144060
rect 202278 105501 202338 144059
rect 202275 105500 202341 105501
rect 202275 105436 202276 105500
rect 202340 105436 202341 105500
rect 202275 105435 202341 105436
rect 202462 104141 202522 145827
rect 202459 104140 202525 104141
rect 202459 104076 202460 104140
rect 202524 104076 202525 104140
rect 202459 104075 202525 104076
rect 202646 102781 202706 146235
rect 202643 102780 202709 102781
rect 202643 102716 202644 102780
rect 202708 102716 202709 102780
rect 202643 102715 202709 102716
rect 203198 98701 203258 157290
rect 203750 146029 203810 158611
rect 203934 153917 203994 158611
rect 203931 153916 203997 153917
rect 203931 153852 203932 153916
rect 203996 153852 203997 153916
rect 203931 153851 203997 153852
rect 203747 146028 203813 146029
rect 203747 145964 203748 146028
rect 203812 145964 203813 146028
rect 203747 145963 203813 145964
rect 203750 122093 203810 145963
rect 203747 122092 203813 122093
rect 203747 122028 203748 122092
rect 203812 122028 203813 122092
rect 203747 122027 203813 122028
rect 203195 98700 203261 98701
rect 203195 98636 203196 98700
rect 203260 98636 203261 98700
rect 203195 98635 203261 98636
rect 204118 97205 204178 159835
rect 204670 159085 204730 165955
rect 204851 163436 204917 163437
rect 204851 163372 204852 163436
rect 204916 163372 204917 163436
rect 204851 163371 204917 163372
rect 204854 159765 204914 163371
rect 205038 159901 205098 166950
rect 205406 159901 205466 177243
rect 205958 159901 206018 190979
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 207611 182884 207677 182885
rect 207611 182820 207612 182884
rect 207676 182820 207677 182884
rect 207611 182819 207677 182820
rect 206875 171732 206941 171733
rect 206875 171668 206876 171732
rect 206940 171668 206941 171732
rect 206875 171667 206941 171668
rect 206507 164932 206573 164933
rect 206507 164868 206508 164932
rect 206572 164868 206573 164932
rect 206507 164867 206573 164868
rect 206510 159901 206570 164867
rect 206691 162212 206757 162213
rect 206691 162148 206692 162212
rect 206756 162148 206757 162212
rect 206691 162147 206757 162148
rect 205035 159900 205101 159901
rect 205035 159836 205036 159900
rect 205100 159898 205101 159900
rect 205403 159900 205469 159901
rect 205100 159838 205282 159898
rect 205100 159836 205101 159838
rect 205035 159835 205101 159836
rect 204851 159764 204917 159765
rect 204851 159700 204852 159764
rect 204916 159700 204917 159764
rect 204851 159699 204917 159700
rect 204667 159084 204733 159085
rect 204667 159020 204668 159084
rect 204732 159020 204733 159084
rect 204667 159019 204733 159020
rect 204670 158405 204730 159019
rect 205035 158676 205101 158677
rect 205035 158612 205036 158676
rect 205100 158612 205101 158676
rect 205035 158611 205101 158612
rect 204667 158404 204733 158405
rect 204667 158340 204668 158404
rect 204732 158340 204733 158404
rect 204667 158339 204733 158340
rect 205038 145757 205098 158611
rect 205035 145756 205101 145757
rect 205035 145692 205036 145756
rect 205100 145692 205101 145756
rect 205035 145691 205101 145692
rect 205038 120733 205098 145691
rect 205035 120732 205101 120733
rect 205035 120668 205036 120732
rect 205100 120668 205101 120732
rect 205035 120667 205101 120668
rect 204115 97204 204181 97205
rect 204115 97140 204116 97204
rect 204180 97140 204181 97204
rect 204115 97139 204181 97140
rect 205222 95845 205282 159838
rect 205403 159836 205404 159900
rect 205468 159836 205469 159900
rect 205403 159835 205469 159836
rect 205955 159900 206021 159901
rect 205955 159836 205956 159900
rect 206020 159836 206021 159900
rect 205955 159835 206021 159836
rect 206507 159900 206573 159901
rect 206507 159836 206508 159900
rect 206572 159836 206573 159900
rect 206507 159835 206573 159836
rect 205219 95844 205285 95845
rect 205219 95780 205220 95844
rect 205284 95780 205285 95844
rect 205219 95779 205285 95780
rect 205406 93125 205466 159835
rect 206694 158269 206754 162147
rect 206878 159901 206938 171667
rect 206875 159900 206941 159901
rect 206875 159836 206876 159900
rect 206940 159836 206941 159900
rect 206875 159835 206941 159836
rect 207614 159765 207674 182819
rect 207979 178668 208045 178669
rect 207979 178604 207980 178668
rect 208044 178604 208045 178668
rect 207979 178603 208045 178604
rect 207795 173228 207861 173229
rect 207795 173164 207796 173228
rect 207860 173164 207861 173228
rect 207795 173163 207861 173164
rect 207798 159901 207858 173163
rect 207795 159900 207861 159901
rect 207795 159836 207796 159900
rect 207860 159836 207861 159900
rect 207795 159835 207861 159836
rect 207611 159764 207677 159765
rect 207611 159700 207612 159764
rect 207676 159700 207677 159764
rect 207611 159699 207677 159700
rect 206691 158268 206757 158269
rect 206691 158204 206692 158268
rect 206756 158204 206757 158268
rect 206691 158203 206757 158204
rect 207982 158133 208042 178603
rect 209083 173364 209149 173365
rect 209083 173300 209084 173364
rect 209148 173300 209149 173364
rect 209083 173299 209149 173300
rect 209086 158677 209146 173299
rect 209267 169148 209333 169149
rect 209267 169084 209268 169148
rect 209332 169084 209333 169148
rect 209267 169083 209333 169084
rect 209083 158676 209149 158677
rect 209083 158612 209084 158676
rect 209148 158612 209149 158676
rect 209083 158611 209149 158612
rect 207979 158132 208045 158133
rect 207979 158068 207980 158132
rect 208044 158068 208045 158132
rect 207979 158067 208045 158068
rect 209270 157725 209330 169083
rect 209267 157724 209333 157725
rect 209267 157660 209268 157724
rect 209332 157660 209333 157724
rect 209267 157659 209333 157660
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 205403 93124 205469 93125
rect 205403 93060 205404 93124
rect 205468 93060 205469 93124
rect 205403 93059 205469 93060
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 201355 39268 201421 39269
rect 201355 39204 201356 39268
rect 201420 39204 201421 39268
rect 201355 39203 201421 39204
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 199883 3364 199949 3365
rect 199883 3300 199884 3364
rect 199948 3300 199949 3364
rect 199883 3299 199949 3300
rect 185514 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 186134 -1306
rect 185514 -1626 186134 -1542
rect 185514 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 186134 -1626
rect 185514 -1894 186134 -1862
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 223174 222134 258618
rect 222702 241773 222762 306851
rect 223067 296172 223133 296173
rect 223067 296108 223068 296172
rect 223132 296108 223133 296172
rect 223067 296107 223133 296108
rect 222699 241772 222765 241773
rect 222699 241708 222700 241772
rect 222764 241708 222765 241772
rect 222699 241707 222765 241708
rect 222515 240412 222581 240413
rect 222515 240348 222516 240412
rect 222580 240348 222581 240412
rect 222515 240347 222581 240348
rect 222518 240005 222578 240347
rect 222515 240004 222581 240005
rect 222515 239940 222516 240004
rect 222580 239940 222581 240004
rect 222515 239939 222581 239940
rect 222702 239461 222762 241707
rect 223070 240005 223130 296107
rect 223067 240004 223133 240005
rect 223067 239940 223068 240004
rect 223132 239940 223133 240004
rect 223067 239939 223133 239940
rect 223254 239869 223314 314059
rect 223251 239868 223317 239869
rect 223251 239804 223252 239868
rect 223316 239804 223317 239868
rect 223251 239803 223317 239804
rect 223438 239733 223498 316915
rect 231715 316844 231781 316845
rect 231715 316780 231716 316844
rect 231780 316780 231781 316844
rect 231715 316779 231781 316780
rect 224723 315620 224789 315621
rect 224723 315556 224724 315620
rect 224788 315556 224789 315620
rect 224723 315555 224789 315556
rect 223987 314260 224053 314261
rect 223987 314196 223988 314260
rect 224052 314196 224053 314260
rect 223987 314195 224053 314196
rect 223803 301612 223869 301613
rect 223803 301548 223804 301612
rect 223868 301548 223869 301612
rect 223803 301547 223869 301548
rect 223619 295356 223685 295357
rect 223619 295292 223620 295356
rect 223684 295292 223685 295356
rect 223619 295291 223685 295292
rect 223622 239733 223682 295291
rect 223806 240005 223866 301547
rect 223990 240005 224050 314195
rect 224171 241364 224237 241365
rect 224171 241300 224172 241364
rect 224236 241300 224237 241364
rect 224171 241299 224237 241300
rect 224174 240549 224234 241299
rect 224171 240548 224237 240549
rect 224171 240484 224172 240548
rect 224236 240484 224237 240548
rect 224171 240483 224237 240484
rect 223803 240004 223869 240005
rect 223803 239940 223804 240004
rect 223868 239940 223869 240004
rect 223803 239939 223869 239940
rect 223987 240004 224053 240005
rect 223987 239940 223988 240004
rect 224052 239940 224053 240004
rect 223987 239939 224053 239940
rect 223435 239732 223501 239733
rect 223435 239668 223436 239732
rect 223500 239668 223501 239732
rect 223435 239667 223501 239668
rect 223619 239732 223685 239733
rect 223619 239668 223620 239732
rect 223684 239668 223685 239732
rect 223619 239667 223685 239668
rect 222699 239460 222765 239461
rect 222699 239396 222700 239460
rect 222764 239396 222765 239460
rect 222699 239395 222765 239396
rect 223806 239053 223866 239939
rect 223803 239052 223869 239053
rect 223803 238988 223804 239052
rect 223868 238988 223869 239052
rect 223803 238987 223869 238988
rect 223990 238237 224050 239939
rect 224174 239869 224234 240483
rect 224726 239869 224786 315555
rect 226195 312764 226261 312765
rect 226195 312700 226196 312764
rect 226260 312700 226261 312764
rect 226195 312699 226261 312700
rect 225459 309772 225525 309773
rect 225459 309708 225460 309772
rect 225524 309708 225525 309772
rect 225459 309707 225525 309708
rect 225275 294676 225341 294677
rect 225275 294612 225276 294676
rect 225340 294612 225341 294676
rect 225275 294611 225341 294612
rect 224171 239868 224237 239869
rect 224171 239804 224172 239868
rect 224236 239804 224237 239868
rect 224171 239803 224237 239804
rect 224723 239868 224789 239869
rect 224723 239804 224724 239868
rect 224788 239804 224789 239868
rect 224723 239803 224789 239804
rect 225091 239868 225157 239869
rect 225091 239804 225092 239868
rect 225156 239804 225157 239868
rect 225091 239803 225157 239804
rect 223987 238236 224053 238237
rect 223987 238172 223988 238236
rect 224052 238172 224053 238236
rect 223987 238171 224053 238172
rect 224723 236332 224789 236333
rect 224723 236268 224724 236332
rect 224788 236268 224789 236332
rect 224723 236267 224789 236268
rect 224726 224970 224786 236267
rect 225094 229805 225154 239803
rect 225278 239597 225338 294611
rect 225462 241637 225522 309707
rect 226011 296444 226077 296445
rect 226011 296380 226012 296444
rect 226076 296380 226077 296444
rect 226011 296379 226077 296380
rect 225459 241636 225525 241637
rect 225459 241572 225460 241636
rect 225524 241572 225525 241636
rect 225459 241571 225525 241572
rect 225275 239596 225341 239597
rect 225275 239532 225276 239596
rect 225340 239532 225341 239596
rect 225275 239531 225341 239532
rect 225462 239053 225522 241571
rect 225643 241500 225709 241501
rect 225643 241436 225644 241500
rect 225708 241436 225709 241500
rect 225643 241435 225709 241436
rect 225646 239325 225706 241435
rect 226014 239461 226074 296379
rect 226198 239869 226258 312699
rect 230059 311540 230125 311541
rect 230059 311476 230060 311540
rect 230124 311476 230125 311540
rect 230059 311475 230125 311476
rect 229323 311132 229389 311133
rect 229323 311068 229324 311132
rect 229388 311068 229389 311132
rect 229323 311067 229389 311068
rect 228955 310316 229021 310317
rect 228955 310252 228956 310316
rect 229020 310252 229021 310316
rect 228955 310251 229021 310252
rect 227483 310180 227549 310181
rect 227483 310116 227484 310180
rect 227548 310116 227549 310180
rect 227483 310115 227549 310116
rect 226379 296308 226445 296309
rect 226379 296244 226380 296308
rect 226444 296244 226445 296308
rect 226379 296243 226445 296244
rect 226382 240005 226442 296243
rect 226563 296036 226629 296037
rect 226563 295972 226564 296036
rect 226628 295972 226629 296036
rect 226563 295971 226629 295972
rect 226379 240004 226445 240005
rect 226379 239940 226380 240004
rect 226444 239940 226445 240004
rect 226379 239939 226445 239940
rect 226195 239868 226261 239869
rect 226195 239804 226196 239868
rect 226260 239804 226261 239868
rect 226195 239803 226261 239804
rect 226382 239597 226442 239939
rect 226379 239596 226445 239597
rect 226379 239532 226380 239596
rect 226444 239532 226445 239596
rect 226379 239531 226445 239532
rect 226566 239461 226626 295971
rect 227299 294812 227365 294813
rect 227299 294748 227300 294812
rect 227364 294748 227365 294812
rect 227299 294747 227365 294748
rect 227302 239869 227362 294747
rect 227299 239868 227365 239869
rect 227299 239804 227300 239868
rect 227364 239804 227365 239868
rect 227299 239803 227365 239804
rect 226747 239732 226813 239733
rect 226747 239668 226748 239732
rect 226812 239668 226813 239732
rect 226747 239667 226813 239668
rect 226011 239460 226077 239461
rect 226011 239396 226012 239460
rect 226076 239396 226077 239460
rect 226011 239395 226077 239396
rect 226563 239460 226629 239461
rect 226563 239396 226564 239460
rect 226628 239396 226629 239460
rect 226563 239395 226629 239396
rect 225643 239324 225709 239325
rect 225643 239260 225644 239324
rect 225708 239260 225709 239324
rect 225643 239259 225709 239260
rect 225459 239052 225525 239053
rect 225459 238988 225460 239052
rect 225524 238988 225525 239052
rect 225459 238987 225525 238988
rect 226750 235925 226810 239667
rect 227302 238237 227362 239803
rect 227486 239461 227546 310115
rect 228219 310044 228285 310045
rect 228219 309980 228220 310044
rect 228284 309980 228285 310044
rect 228219 309979 228285 309980
rect 227667 240956 227733 240957
rect 227667 240892 227668 240956
rect 227732 240892 227733 240956
rect 227667 240891 227733 240892
rect 227670 239733 227730 240891
rect 227667 239732 227733 239733
rect 227667 239668 227668 239732
rect 227732 239668 227733 239732
rect 227667 239667 227733 239668
rect 227483 239460 227549 239461
rect 227483 239396 227484 239460
rect 227548 239396 227549 239460
rect 227483 239395 227549 239396
rect 227299 238236 227365 238237
rect 227299 238172 227300 238236
rect 227364 238172 227365 238236
rect 227299 238171 227365 238172
rect 227115 238100 227181 238101
rect 227115 238036 227116 238100
rect 227180 238036 227181 238100
rect 227115 238035 227181 238036
rect 226747 235924 226813 235925
rect 226747 235860 226748 235924
rect 226812 235860 226813 235924
rect 226747 235859 226813 235860
rect 227118 234630 227178 238035
rect 226934 234570 227178 234630
rect 225091 229804 225157 229805
rect 225091 229740 225092 229804
rect 225156 229740 225157 229804
rect 225091 229739 225157 229740
rect 224726 224910 225154 224970
rect 225094 223549 225154 224910
rect 225091 223548 225157 223549
rect 225091 223484 225092 223548
rect 225156 223484 225157 223548
rect 225091 223483 225157 223484
rect 221514 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 222134 223174
rect 221514 222854 222134 222938
rect 221514 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 222134 222854
rect 221514 187174 222134 222618
rect 221514 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 222134 187174
rect 221514 186854 222134 186938
rect 221514 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 222134 186854
rect 221514 151174 222134 186618
rect 226934 151197 226994 234570
rect 227670 225997 227730 239667
rect 228222 239461 228282 309979
rect 228587 299028 228653 299029
rect 228587 298964 228588 299028
rect 228652 298964 228653 299028
rect 228587 298963 228653 298964
rect 228403 294540 228469 294541
rect 228403 294476 228404 294540
rect 228468 294476 228469 294540
rect 228403 294475 228469 294476
rect 227851 239460 227917 239461
rect 227851 239396 227852 239460
rect 227916 239396 227917 239460
rect 227851 239395 227917 239396
rect 228219 239460 228285 239461
rect 228219 239396 228220 239460
rect 228284 239396 228285 239460
rect 228219 239395 228285 239396
rect 227854 231709 227914 239395
rect 228406 238781 228466 294475
rect 228590 239733 228650 298963
rect 228587 239732 228653 239733
rect 228587 239668 228588 239732
rect 228652 239668 228653 239732
rect 228587 239667 228653 239668
rect 228958 239597 229018 310251
rect 229139 240820 229205 240821
rect 229139 240756 229140 240820
rect 229204 240756 229205 240820
rect 229139 240755 229205 240756
rect 229142 239733 229202 240755
rect 229139 239732 229205 239733
rect 229139 239668 229140 239732
rect 229204 239668 229205 239732
rect 229139 239667 229205 239668
rect 228955 239596 229021 239597
rect 228955 239532 228956 239596
rect 229020 239532 229021 239596
rect 228955 239531 229021 239532
rect 229326 239461 229386 311067
rect 229507 294948 229573 294949
rect 229507 294884 229508 294948
rect 229572 294884 229573 294948
rect 229507 294883 229573 294884
rect 229510 239869 229570 294883
rect 229875 294268 229941 294269
rect 229875 294204 229876 294268
rect 229940 294204 229941 294268
rect 229875 294203 229941 294204
rect 229507 239868 229573 239869
rect 229507 239804 229508 239868
rect 229572 239804 229573 239868
rect 229507 239803 229573 239804
rect 229510 239597 229570 239803
rect 229878 239733 229938 294203
rect 230062 239869 230122 311475
rect 231347 311404 231413 311405
rect 231347 311340 231348 311404
rect 231412 311340 231413 311404
rect 231347 311339 231413 311340
rect 231163 311268 231229 311269
rect 231163 311204 231164 311268
rect 231228 311204 231229 311268
rect 231163 311203 231229 311204
rect 230795 241228 230861 241229
rect 230795 241164 230796 241228
rect 230860 241164 230861 241228
rect 230795 241163 230861 241164
rect 230427 240548 230493 240549
rect 230427 240484 230428 240548
rect 230492 240484 230493 240548
rect 230427 240483 230493 240484
rect 230059 239868 230125 239869
rect 230059 239804 230060 239868
rect 230124 239804 230125 239868
rect 230059 239803 230125 239804
rect 229875 239732 229941 239733
rect 229875 239668 229876 239732
rect 229940 239668 229941 239732
rect 229875 239667 229941 239668
rect 229507 239596 229573 239597
rect 229507 239532 229508 239596
rect 229572 239532 229573 239596
rect 229507 239531 229573 239532
rect 229323 239460 229389 239461
rect 229323 239396 229324 239460
rect 229388 239396 229389 239460
rect 229323 239395 229389 239396
rect 228403 238780 228469 238781
rect 228403 238716 228404 238780
rect 228468 238716 228469 238780
rect 228403 238715 228469 238716
rect 229691 237828 229757 237829
rect 229691 237764 229692 237828
rect 229756 237764 229757 237828
rect 229691 237763 229757 237764
rect 229694 236469 229754 237763
rect 229691 236468 229757 236469
rect 229691 236404 229692 236468
rect 229756 236404 229757 236468
rect 229691 236403 229757 236404
rect 229878 236061 229938 239667
rect 230062 237557 230122 239803
rect 230430 239461 230490 240483
rect 230798 239733 230858 241163
rect 230979 240140 231045 240141
rect 230979 240076 230980 240140
rect 231044 240076 231045 240140
rect 230979 240075 231045 240076
rect 230982 239869 231042 240075
rect 230979 239868 231045 239869
rect 230979 239804 230980 239868
rect 231044 239804 231045 239868
rect 230979 239803 231045 239804
rect 230795 239732 230861 239733
rect 230795 239668 230796 239732
rect 230860 239668 230861 239732
rect 230795 239667 230861 239668
rect 231166 239597 231226 311203
rect 231350 239733 231410 311339
rect 231531 289916 231597 289917
rect 231531 289852 231532 289916
rect 231596 289852 231597 289916
rect 231531 289851 231597 289852
rect 231534 288421 231594 289851
rect 231531 288420 231597 288421
rect 231531 288356 231532 288420
rect 231596 288356 231597 288420
rect 231531 288355 231597 288356
rect 231534 287741 231594 288355
rect 231531 287740 231597 287741
rect 231531 287676 231532 287740
rect 231596 287676 231597 287740
rect 231531 287675 231597 287676
rect 231718 239869 231778 316779
rect 237235 315892 237301 315893
rect 237235 315828 237236 315892
rect 237300 315828 237301 315892
rect 237235 315827 237301 315828
rect 235211 315756 235277 315757
rect 235211 315692 235212 315756
rect 235276 315692 235277 315756
rect 235211 315691 235277 315692
rect 232267 314532 232333 314533
rect 232267 314468 232268 314532
rect 232332 314468 232333 314532
rect 232267 314467 232333 314468
rect 232083 241092 232149 241093
rect 232083 241028 232084 241092
rect 232148 241028 232149 241092
rect 232083 241027 232149 241028
rect 231715 239868 231781 239869
rect 231715 239804 231716 239868
rect 231780 239804 231781 239868
rect 231715 239803 231781 239804
rect 231347 239732 231413 239733
rect 231347 239668 231348 239732
rect 231412 239668 231413 239732
rect 231347 239667 231413 239668
rect 231531 239732 231597 239733
rect 231531 239668 231532 239732
rect 231596 239668 231597 239732
rect 231531 239667 231597 239668
rect 231163 239596 231229 239597
rect 231163 239532 231164 239596
rect 231228 239532 231229 239596
rect 231163 239531 231229 239532
rect 230427 239460 230493 239461
rect 230427 239396 230428 239460
rect 230492 239396 230493 239460
rect 230427 239395 230493 239396
rect 231163 238780 231229 238781
rect 231163 238716 231164 238780
rect 231228 238716 231229 238780
rect 231163 238715 231229 238716
rect 230611 237964 230677 237965
rect 230611 237900 230612 237964
rect 230676 237900 230677 237964
rect 230611 237899 230677 237900
rect 230059 237556 230125 237557
rect 230059 237492 230060 237556
rect 230124 237492 230125 237556
rect 230059 237491 230125 237492
rect 229875 236060 229941 236061
rect 229875 235996 229876 236060
rect 229940 235996 229941 236060
rect 229875 235995 229941 235996
rect 230614 235789 230674 237899
rect 230611 235788 230677 235789
rect 230611 235724 230612 235788
rect 230676 235724 230677 235788
rect 230611 235723 230677 235724
rect 227851 231708 227917 231709
rect 227851 231644 227852 231708
rect 227916 231644 227917 231708
rect 227851 231643 227917 231644
rect 227667 225996 227733 225997
rect 227667 225932 227668 225996
rect 227732 225932 227733 225996
rect 227667 225931 227733 225932
rect 231166 220693 231226 238715
rect 230427 220692 230493 220693
rect 230427 220628 230428 220692
rect 230492 220628 230493 220692
rect 230427 220627 230493 220628
rect 231163 220692 231229 220693
rect 231163 220628 231164 220692
rect 231228 220628 231229 220692
rect 231163 220627 231229 220628
rect 230430 220149 230490 220627
rect 231534 220557 231594 239667
rect 231718 238237 231778 239803
rect 232086 239733 232146 241027
rect 232083 239732 232149 239733
rect 232083 239668 232084 239732
rect 232148 239668 232149 239732
rect 232083 239667 232149 239668
rect 232270 239597 232330 314467
rect 232819 313988 232885 313989
rect 232819 313924 232820 313988
rect 232884 313924 232885 313988
rect 232819 313923 232885 313924
rect 232635 311676 232701 311677
rect 232635 311612 232636 311676
rect 232700 311612 232701 311676
rect 232635 311611 232701 311612
rect 232451 294404 232517 294405
rect 232451 294340 232452 294404
rect 232516 294340 232517 294404
rect 232451 294339 232517 294340
rect 232267 239596 232333 239597
rect 232267 239532 232268 239596
rect 232332 239532 232333 239596
rect 232267 239531 232333 239532
rect 232454 238781 232514 294339
rect 232638 239869 232698 311611
rect 232822 239869 232882 313923
rect 234291 312628 234357 312629
rect 234291 312564 234292 312628
rect 234356 312564 234357 312628
rect 234291 312563 234357 312564
rect 234107 308412 234173 308413
rect 234107 308348 234108 308412
rect 234172 308348 234173 308412
rect 234107 308347 234173 308348
rect 233923 298756 233989 298757
rect 233923 298692 233924 298756
rect 233988 298692 233989 298756
rect 233923 298691 233989 298692
rect 233371 241092 233437 241093
rect 233371 241028 233372 241092
rect 233436 241028 233437 241092
rect 233371 241027 233437 241028
rect 233187 240684 233253 240685
rect 233187 240620 233188 240684
rect 233252 240620 233253 240684
rect 233187 240619 233253 240620
rect 233003 240412 233069 240413
rect 233003 240348 233004 240412
rect 233068 240348 233069 240412
rect 233003 240347 233069 240348
rect 232635 239868 232701 239869
rect 232635 239804 232636 239868
rect 232700 239804 232701 239868
rect 232635 239803 232701 239804
rect 232819 239868 232885 239869
rect 232819 239804 232820 239868
rect 232884 239804 232885 239868
rect 232819 239803 232885 239804
rect 232451 238780 232517 238781
rect 232451 238716 232452 238780
rect 232516 238716 232517 238780
rect 232451 238715 232517 238716
rect 231715 238236 231781 238237
rect 231715 238172 231716 238236
rect 231780 238172 231781 238236
rect 231715 238171 231781 238172
rect 232451 236604 232517 236605
rect 232451 236540 232452 236604
rect 232516 236540 232517 236604
rect 232451 236539 232517 236540
rect 230979 220556 231045 220557
rect 230979 220492 230980 220556
rect 231044 220492 231045 220556
rect 230979 220491 231045 220492
rect 231531 220556 231597 220557
rect 231531 220492 231532 220556
rect 231596 220492 231597 220556
rect 231531 220491 231597 220492
rect 230427 220148 230493 220149
rect 230427 220084 230428 220148
rect 230492 220084 230493 220148
rect 230427 220083 230493 220084
rect 221514 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 222134 151174
rect 226931 151196 226997 151197
rect 226931 151132 226932 151196
rect 226996 151132 226997 151196
rect 226931 151131 226997 151132
rect 221514 150854 222134 150938
rect 221514 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 222134 150854
rect 221514 115174 222134 150618
rect 230982 144533 231042 220491
rect 232454 147117 232514 236539
rect 232638 235789 232698 239803
rect 233006 239597 233066 240347
rect 233190 239733 233250 240619
rect 233374 239869 233434 241027
rect 233739 240684 233805 240685
rect 233739 240620 233740 240684
rect 233804 240620 233805 240684
rect 233739 240619 233805 240620
rect 233371 239868 233437 239869
rect 233371 239804 233372 239868
rect 233436 239804 233437 239868
rect 233371 239803 233437 239804
rect 233187 239732 233253 239733
rect 233187 239668 233188 239732
rect 233252 239668 233253 239732
rect 233187 239667 233253 239668
rect 233003 239596 233069 239597
rect 233003 239532 233004 239596
rect 233068 239532 233069 239596
rect 233003 239531 233069 239532
rect 232635 235788 232701 235789
rect 232635 235724 232636 235788
rect 232700 235724 232701 235788
rect 232635 235723 232701 235724
rect 233374 234021 233434 239803
rect 233742 239733 233802 240619
rect 233926 239869 233986 298691
rect 233923 239868 233989 239869
rect 233923 239804 233924 239868
rect 233988 239804 233989 239868
rect 233923 239803 233989 239804
rect 233739 239732 233805 239733
rect 233739 239668 233740 239732
rect 233804 239668 233805 239732
rect 233739 239667 233805 239668
rect 233742 238781 233802 239667
rect 233739 238780 233805 238781
rect 233739 238716 233740 238780
rect 233804 238716 233805 238780
rect 233739 238715 233805 238716
rect 233926 238645 233986 239803
rect 234110 239733 234170 308347
rect 234107 239732 234173 239733
rect 234107 239668 234108 239732
rect 234172 239668 234173 239732
rect 234107 239667 234173 239668
rect 234294 239461 234354 312563
rect 234475 312356 234541 312357
rect 234475 312292 234476 312356
rect 234540 312292 234541 312356
rect 234475 312291 234541 312292
rect 234478 240685 234538 312291
rect 235027 298892 235093 298893
rect 235027 298828 235028 298892
rect 235092 298828 235093 298892
rect 235027 298827 235093 298828
rect 234843 240820 234909 240821
rect 234843 240756 234844 240820
rect 234908 240756 234909 240820
rect 234843 240755 234909 240756
rect 234475 240684 234541 240685
rect 234475 240620 234476 240684
rect 234540 240620 234541 240684
rect 234475 240619 234541 240620
rect 234846 239869 234906 240755
rect 234843 239868 234909 239869
rect 234843 239804 234844 239868
rect 234908 239804 234909 239868
rect 234843 239803 234909 239804
rect 235030 239733 235090 298827
rect 235027 239732 235093 239733
rect 235027 239668 235028 239732
rect 235092 239668 235093 239732
rect 235027 239667 235093 239668
rect 235214 239461 235274 315691
rect 237051 315620 237117 315621
rect 237051 315556 237052 315620
rect 237116 315556 237117 315620
rect 237051 315555 237117 315556
rect 236867 307732 236933 307733
rect 236867 307668 236868 307732
rect 236932 307668 236933 307732
rect 236867 307667 236933 307668
rect 235579 304468 235645 304469
rect 235579 304404 235580 304468
rect 235644 304404 235645 304468
rect 235579 304403 235645 304404
rect 235395 301476 235461 301477
rect 235395 301412 235396 301476
rect 235460 301412 235461 301476
rect 235395 301411 235461 301412
rect 235398 239733 235458 301411
rect 235395 239732 235461 239733
rect 235395 239668 235396 239732
rect 235460 239668 235461 239732
rect 235395 239667 235461 239668
rect 234291 239460 234357 239461
rect 234291 239396 234292 239460
rect 234356 239396 234357 239460
rect 235211 239460 235277 239461
rect 235211 239458 235212 239460
rect 234291 239395 234357 239396
rect 235030 239398 235212 239458
rect 233923 238644 233989 238645
rect 233923 238580 233924 238644
rect 233988 238580 233989 238644
rect 233923 238579 233989 238580
rect 234291 238508 234357 238509
rect 234291 238444 234292 238508
rect 234356 238444 234357 238508
rect 234291 238443 234357 238444
rect 233555 238236 233621 238237
rect 233555 238172 233556 238236
rect 233620 238172 233621 238236
rect 233555 238171 233621 238172
rect 233371 234020 233437 234021
rect 233371 233956 233372 234020
rect 233436 233956 233437 234020
rect 233371 233955 233437 233956
rect 233558 221917 233618 238171
rect 234294 238101 234354 238443
rect 234291 238100 234357 238101
rect 234291 238036 234292 238100
rect 234356 238036 234357 238100
rect 234291 238035 234357 238036
rect 233739 236060 233805 236061
rect 233739 235996 233740 236060
rect 233804 235996 233805 236060
rect 233739 235995 233805 235996
rect 234475 236060 234541 236061
rect 234475 235996 234476 236060
rect 234540 235996 234541 236060
rect 234475 235995 234541 235996
rect 233742 225861 233802 235995
rect 234478 231709 234538 235995
rect 235030 235517 235090 239398
rect 235211 239396 235212 239398
rect 235276 239396 235277 239460
rect 235211 239395 235277 239396
rect 235211 236332 235277 236333
rect 235211 236268 235212 236332
rect 235276 236268 235277 236332
rect 235211 236267 235277 236268
rect 235027 235516 235093 235517
rect 235027 235452 235028 235516
rect 235092 235452 235093 235516
rect 235027 235451 235093 235452
rect 234475 231708 234541 231709
rect 234475 231644 234476 231708
rect 234540 231644 234541 231708
rect 234475 231643 234541 231644
rect 233739 225860 233805 225861
rect 233739 225796 233740 225860
rect 233804 225796 233805 225860
rect 233739 225795 233805 225796
rect 233187 221916 233253 221917
rect 233187 221852 233188 221916
rect 233252 221852 233253 221916
rect 233187 221851 233253 221852
rect 233555 221916 233621 221917
rect 233555 221852 233556 221916
rect 233620 221852 233621 221916
rect 233555 221851 233621 221852
rect 233190 221509 233250 221851
rect 233187 221508 233253 221509
rect 233187 221444 233188 221508
rect 233252 221444 233253 221508
rect 233187 221443 233253 221444
rect 233742 147525 233802 225795
rect 234478 225589 234538 231643
rect 234475 225588 234541 225589
rect 234475 225524 234476 225588
rect 234540 225524 234541 225588
rect 234475 225523 234541 225524
rect 233739 147524 233805 147525
rect 233739 147460 233740 147524
rect 233804 147460 233805 147524
rect 233739 147459 233805 147460
rect 232451 147116 232517 147117
rect 232451 147052 232452 147116
rect 232516 147052 232517 147116
rect 232451 147051 232517 147052
rect 235214 144805 235274 236267
rect 235398 233749 235458 239667
rect 235582 238781 235642 304403
rect 235947 293180 236013 293181
rect 235947 293116 235948 293180
rect 236012 293116 236013 293180
rect 235947 293115 236013 293116
rect 235950 266370 236010 293115
rect 235950 266310 236378 266370
rect 236131 239732 236197 239733
rect 236131 239668 236132 239732
rect 236196 239668 236197 239732
rect 236131 239667 236197 239668
rect 235579 238780 235645 238781
rect 235579 238716 235580 238780
rect 235644 238716 235645 238780
rect 235579 238715 235645 238716
rect 236134 238237 236194 239667
rect 236318 239461 236378 266310
rect 236683 240004 236749 240005
rect 236683 239940 236684 240004
rect 236748 239940 236749 240004
rect 236683 239939 236749 239940
rect 236315 239460 236381 239461
rect 236315 239396 236316 239460
rect 236380 239396 236381 239460
rect 236315 239395 236381 239396
rect 236686 238237 236746 239939
rect 236870 239869 236930 307667
rect 236867 239868 236933 239869
rect 236867 239804 236868 239868
rect 236932 239804 236933 239868
rect 236867 239803 236933 239804
rect 236131 238236 236197 238237
rect 236131 238172 236132 238236
rect 236196 238172 236197 238236
rect 236131 238171 236197 238172
rect 236683 238236 236749 238237
rect 236683 238172 236684 238236
rect 236748 238172 236749 238236
rect 236683 238171 236749 238172
rect 236870 237557 236930 239803
rect 237054 239461 237114 315555
rect 237238 239733 237298 315827
rect 237974 253950 238034 318003
rect 241099 314396 241165 314397
rect 241099 314332 241100 314396
rect 241164 314332 241165 314396
rect 241099 314331 241165 314332
rect 239443 313852 239509 313853
rect 239443 313788 239444 313852
rect 239508 313788 239509 313852
rect 239443 313787 239509 313788
rect 238523 308548 238589 308549
rect 238523 308484 238524 308548
rect 238588 308484 238589 308548
rect 238523 308483 238589 308484
rect 238339 300116 238405 300117
rect 238339 300052 238340 300116
rect 238404 300052 238405 300116
rect 238339 300051 238405 300052
rect 238155 293452 238221 293453
rect 238155 293388 238156 293452
rect 238220 293388 238221 293452
rect 238155 293387 238221 293388
rect 237790 253890 238034 253950
rect 237790 240549 237850 253890
rect 237971 240684 238037 240685
rect 237971 240620 237972 240684
rect 238036 240620 238037 240684
rect 237971 240619 238037 240620
rect 237787 240548 237853 240549
rect 237787 240484 237788 240548
rect 237852 240484 237853 240548
rect 237787 240483 237853 240484
rect 237974 239869 238034 240619
rect 237971 239868 238037 239869
rect 237971 239804 237972 239868
rect 238036 239804 238037 239868
rect 237971 239803 238037 239804
rect 237235 239732 237301 239733
rect 237235 239668 237236 239732
rect 237300 239668 237301 239732
rect 237235 239667 237301 239668
rect 238158 239461 238218 293387
rect 238342 239733 238402 300051
rect 238339 239732 238405 239733
rect 238339 239668 238340 239732
rect 238404 239668 238405 239732
rect 238339 239667 238405 239668
rect 238526 239461 238586 308483
rect 238707 306508 238773 306509
rect 238707 306444 238708 306508
rect 238772 306444 238773 306508
rect 238707 306443 238773 306444
rect 238710 306237 238770 306443
rect 238707 306236 238773 306237
rect 238707 306172 238708 306236
rect 238772 306172 238773 306236
rect 238707 306171 238773 306172
rect 239259 302292 239325 302293
rect 239259 302228 239260 302292
rect 239324 302228 239325 302292
rect 239259 302227 239325 302228
rect 238891 296852 238957 296853
rect 238891 296850 238892 296852
rect 238710 296790 238892 296850
rect 238710 296581 238770 296790
rect 238891 296788 238892 296790
rect 238956 296788 238957 296852
rect 238891 296787 238957 296788
rect 238707 296580 238773 296581
rect 238707 296516 238708 296580
rect 238772 296516 238773 296580
rect 238707 296515 238773 296516
rect 239075 293316 239141 293317
rect 239075 293252 239076 293316
rect 239140 293252 239141 293316
rect 239075 293251 239141 293252
rect 238891 290188 238957 290189
rect 238891 290124 238892 290188
rect 238956 290124 238957 290188
rect 238891 290123 238957 290124
rect 238707 239732 238773 239733
rect 238707 239668 238708 239732
rect 238772 239668 238773 239732
rect 238707 239667 238773 239668
rect 237051 239460 237117 239461
rect 237051 239396 237052 239460
rect 237116 239396 237117 239460
rect 237051 239395 237117 239396
rect 238155 239460 238221 239461
rect 238155 239396 238156 239460
rect 238220 239396 238221 239460
rect 238155 239395 238221 239396
rect 238523 239460 238589 239461
rect 238523 239396 238524 239460
rect 238588 239396 238589 239460
rect 238523 239395 238589 239396
rect 236867 237556 236933 237557
rect 236867 237492 236868 237556
rect 236932 237492 236933 237556
rect 236867 237491 236933 237492
rect 236499 236876 236565 236877
rect 236499 236812 236500 236876
rect 236564 236812 236565 236876
rect 236499 236811 236565 236812
rect 235395 233748 235461 233749
rect 235395 233684 235396 233748
rect 235460 233684 235461 233748
rect 235395 233683 235461 233684
rect 236502 152693 236562 236811
rect 237054 236197 237114 239395
rect 237051 236196 237117 236197
rect 237051 236132 237052 236196
rect 237116 236132 237117 236196
rect 237051 236131 237117 236132
rect 238526 235789 238586 239395
rect 238523 235788 238589 235789
rect 238523 235724 238524 235788
rect 238588 235724 238589 235788
rect 238523 235723 238589 235724
rect 238710 234630 238770 239667
rect 238894 239461 238954 290123
rect 239078 239869 239138 293251
rect 239075 239868 239141 239869
rect 239075 239804 239076 239868
rect 239140 239804 239141 239868
rect 239075 239803 239141 239804
rect 238891 239460 238957 239461
rect 238891 239396 238892 239460
rect 238956 239396 238957 239460
rect 238891 239395 238957 239396
rect 238526 234570 238770 234630
rect 236499 152692 236565 152693
rect 236499 152628 236500 152692
rect 236564 152628 236565 152692
rect 236499 152627 236565 152628
rect 235211 144804 235277 144805
rect 235211 144740 235212 144804
rect 235276 144740 235277 144804
rect 235211 144739 235277 144740
rect 230979 144532 231045 144533
rect 230979 144468 230980 144532
rect 231044 144468 231045 144532
rect 230979 144467 231045 144468
rect 238526 142170 238586 234570
rect 238894 218653 238954 239395
rect 239078 236741 239138 239803
rect 239262 239461 239322 302227
rect 239259 239460 239325 239461
rect 239259 239396 239260 239460
rect 239324 239396 239325 239460
rect 239259 239395 239325 239396
rect 239262 238237 239322 239395
rect 239446 238781 239506 313787
rect 240915 301748 240981 301749
rect 240915 301684 240916 301748
rect 240980 301684 240981 301748
rect 240915 301683 240981 301684
rect 239811 240276 239877 240277
rect 239811 240212 239812 240276
rect 239876 240212 239877 240276
rect 239811 240211 239877 240212
rect 239627 240004 239693 240005
rect 239627 239940 239628 240004
rect 239692 239940 239693 240004
rect 239627 239939 239693 239940
rect 239443 238780 239509 238781
rect 239443 238716 239444 238780
rect 239508 238716 239509 238780
rect 239443 238715 239509 238716
rect 239259 238236 239325 238237
rect 239259 238172 239260 238236
rect 239324 238172 239325 238236
rect 239259 238171 239325 238172
rect 239075 236740 239141 236741
rect 239075 236676 239076 236740
rect 239140 236676 239141 236740
rect 239075 236675 239141 236676
rect 238891 218652 238957 218653
rect 238891 218588 238892 218652
rect 238956 218588 238957 218652
rect 238891 218587 238957 218588
rect 239446 211853 239506 238715
rect 239630 237557 239690 239939
rect 239814 239461 239874 240211
rect 240179 239868 240245 239869
rect 240179 239804 240180 239868
rect 240244 239804 240245 239868
rect 240179 239803 240245 239804
rect 240547 239868 240613 239869
rect 240547 239804 240548 239868
rect 240612 239804 240613 239868
rect 240547 239803 240613 239804
rect 239811 239460 239877 239461
rect 239811 239396 239812 239460
rect 239876 239396 239877 239460
rect 239811 239395 239877 239396
rect 239627 237556 239693 237557
rect 239627 237492 239628 237556
rect 239692 237492 239693 237556
rect 239627 237491 239693 237492
rect 239627 235516 239693 235517
rect 239627 235452 239628 235516
rect 239692 235452 239693 235516
rect 239627 235451 239693 235452
rect 239630 223005 239690 235451
rect 240182 224909 240242 239803
rect 240550 233205 240610 239803
rect 240918 238781 240978 301683
rect 241102 239869 241162 314331
rect 244595 314124 244661 314125
rect 244595 314060 244596 314124
rect 244660 314060 244661 314124
rect 244595 314059 244661 314060
rect 241283 313716 241349 313717
rect 241283 313652 241284 313716
rect 241348 313652 241349 313716
rect 241283 313651 241349 313652
rect 241099 239868 241165 239869
rect 241099 239804 241100 239868
rect 241164 239804 241165 239868
rect 241099 239803 241165 239804
rect 240915 238780 240981 238781
rect 240915 238716 240916 238780
rect 240980 238716 240981 238780
rect 240915 238715 240981 238716
rect 241102 238645 241162 239803
rect 241099 238644 241165 238645
rect 241099 238580 241100 238644
rect 241164 238580 241165 238644
rect 241099 238579 241165 238580
rect 241286 238237 241346 313651
rect 242939 293588 243005 293589
rect 242939 293524 242940 293588
rect 243004 293524 243005 293588
rect 242939 293523 243005 293524
rect 241835 241908 241901 241909
rect 241835 241844 241836 241908
rect 241900 241844 241901 241908
rect 241835 241843 241901 241844
rect 241838 240141 241898 241843
rect 241835 240140 241901 240141
rect 241835 240076 241836 240140
rect 241900 240076 241901 240140
rect 241835 240075 241901 240076
rect 242019 240140 242085 240141
rect 242019 240076 242020 240140
rect 242084 240076 242085 240140
rect 242019 240075 242085 240076
rect 241283 238236 241349 238237
rect 241283 238172 241284 238236
rect 241348 238172 241349 238236
rect 241283 238171 241349 238172
rect 240731 236740 240797 236741
rect 240731 236676 240732 236740
rect 240796 236676 240797 236740
rect 240731 236675 240797 236676
rect 241835 236740 241901 236741
rect 241835 236676 241836 236740
rect 241900 236676 241901 236740
rect 241835 236675 241901 236676
rect 240547 233204 240613 233205
rect 240547 233140 240548 233204
rect 240612 233140 240613 233204
rect 240547 233139 240613 233140
rect 240179 224908 240245 224909
rect 240179 224844 240180 224908
rect 240244 224844 240245 224908
rect 240179 224843 240245 224844
rect 239627 223004 239693 223005
rect 239627 222940 239628 223004
rect 239692 222940 239693 223004
rect 239627 222939 239693 222940
rect 240734 222869 240794 236675
rect 241838 230349 241898 236675
rect 241835 230348 241901 230349
rect 241835 230284 241836 230348
rect 241900 230284 241901 230348
rect 241835 230283 241901 230284
rect 240731 222868 240797 222869
rect 240731 222804 240732 222868
rect 240796 222804 240797 222868
rect 240731 222803 240797 222804
rect 239443 211852 239509 211853
rect 239443 211788 239444 211852
rect 239508 211788 239509 211852
rect 239443 211787 239509 211788
rect 238526 142110 238770 142170
rect 238710 141813 238770 142110
rect 240734 141949 240794 222803
rect 242022 143173 242082 240075
rect 242942 239733 243002 293523
rect 244227 290188 244293 290189
rect 244227 290124 244228 290188
rect 244292 290124 244293 290188
rect 244227 290123 244293 290124
rect 244230 289781 244290 290123
rect 244227 289780 244293 289781
rect 244227 289716 244228 289780
rect 244292 289716 244293 289780
rect 244227 289715 244293 289716
rect 244598 239733 244658 314059
rect 244779 309908 244845 309909
rect 244779 309844 244780 309908
rect 244844 309844 244845 309908
rect 244779 309843 244845 309844
rect 242939 239732 243005 239733
rect 242939 239668 242940 239732
rect 243004 239668 243005 239732
rect 242939 239667 243005 239668
rect 244595 239732 244661 239733
rect 244595 239668 244596 239732
rect 244660 239668 244661 239732
rect 244595 239667 244661 239668
rect 244782 239461 244842 309843
rect 246435 301612 246501 301613
rect 246435 301548 246436 301612
rect 246500 301548 246501 301612
rect 246435 301547 246501 301548
rect 245147 290868 245213 290869
rect 245147 290804 245148 290868
rect 245212 290804 245213 290868
rect 245147 290803 245213 290804
rect 244963 289780 245029 289781
rect 244963 289716 244964 289780
rect 245028 289716 245029 289780
rect 244963 289715 245029 289716
rect 244966 239869 245026 289715
rect 245150 239869 245210 290803
rect 246251 290460 246317 290461
rect 246251 290396 246252 290460
rect 246316 290396 246317 290460
rect 246251 290395 246317 290396
rect 245331 289508 245397 289509
rect 245331 289444 245332 289508
rect 245396 289444 245397 289508
rect 245331 289443 245397 289444
rect 245334 289101 245394 289443
rect 245331 289100 245397 289101
rect 245331 289036 245332 289100
rect 245396 289036 245397 289100
rect 245331 289035 245397 289036
rect 245699 242044 245765 242045
rect 245699 241980 245700 242044
rect 245764 241980 245765 242044
rect 245699 241979 245765 241980
rect 244963 239868 245029 239869
rect 244963 239804 244964 239868
rect 245028 239804 245029 239868
rect 244963 239803 245029 239804
rect 245147 239868 245213 239869
rect 245147 239804 245148 239868
rect 245212 239804 245213 239868
rect 245147 239803 245213 239804
rect 245331 239732 245397 239733
rect 245331 239668 245332 239732
rect 245396 239668 245397 239732
rect 245331 239667 245397 239668
rect 243123 239460 243189 239461
rect 243123 239396 243124 239460
rect 243188 239396 243189 239460
rect 243123 239395 243189 239396
rect 244779 239460 244845 239461
rect 244779 239396 244780 239460
rect 244844 239396 244845 239460
rect 244779 239395 244845 239396
rect 242387 238236 242453 238237
rect 242387 238172 242388 238236
rect 242452 238172 242453 238236
rect 242387 238171 242453 238172
rect 242390 228309 242450 238171
rect 243126 234701 243186 239395
rect 245334 238645 245394 239667
rect 245702 238781 245762 241979
rect 246254 240141 246314 290395
rect 246251 240140 246317 240141
rect 246251 240076 246252 240140
rect 246316 240076 246317 240140
rect 246251 240075 246317 240076
rect 246438 239869 246498 301547
rect 247542 241501 247602 318275
rect 247907 313172 247973 313173
rect 247907 313108 247908 313172
rect 247972 313108 247973 313172
rect 247907 313107 247973 313108
rect 247539 241500 247605 241501
rect 247539 241436 247540 241500
rect 247604 241436 247605 241500
rect 247539 241435 247605 241436
rect 245883 239868 245949 239869
rect 245883 239804 245884 239868
rect 245948 239804 245949 239868
rect 245883 239803 245949 239804
rect 246435 239868 246501 239869
rect 246435 239804 246436 239868
rect 246500 239804 246501 239868
rect 246435 239803 246501 239804
rect 245699 238780 245765 238781
rect 245699 238716 245700 238780
rect 245764 238716 245765 238780
rect 245699 238715 245765 238716
rect 245331 238644 245397 238645
rect 245331 238580 245332 238644
rect 245396 238580 245397 238644
rect 245331 238579 245397 238580
rect 244779 235380 244845 235381
rect 244779 235316 244780 235380
rect 244844 235316 244845 235380
rect 244779 235315 244845 235316
rect 243123 234700 243189 234701
rect 243123 234636 243124 234700
rect 243188 234636 243189 234700
rect 243123 234635 243189 234636
rect 242387 228308 242453 228309
rect 242387 228244 242388 228308
rect 242452 228244 242453 228308
rect 242387 228243 242453 228244
rect 243126 226133 243186 234635
rect 243123 226132 243189 226133
rect 243123 226068 243124 226132
rect 243188 226068 243189 226132
rect 243123 226067 243189 226068
rect 243126 225045 243186 226067
rect 243123 225044 243189 225045
rect 243123 224980 243124 225044
rect 243188 224980 243189 225044
rect 243123 224979 243189 224980
rect 244782 157997 244842 235315
rect 245886 226350 245946 239803
rect 247910 239733 247970 313107
rect 249563 313036 249629 313037
rect 249563 312972 249564 313036
rect 249628 312972 249629 313036
rect 249563 312971 249629 312972
rect 248091 291820 248157 291821
rect 248091 291756 248092 291820
rect 248156 291756 248157 291820
rect 248091 291755 248157 291756
rect 246803 239732 246869 239733
rect 246803 239668 246804 239732
rect 246868 239668 246869 239732
rect 246803 239667 246869 239668
rect 247907 239732 247973 239733
rect 247907 239668 247908 239732
rect 247972 239668 247973 239732
rect 247907 239667 247973 239668
rect 246435 233204 246501 233205
rect 246435 233140 246436 233204
rect 246500 233140 246501 233204
rect 246435 233139 246501 233140
rect 245702 226290 245946 226350
rect 245702 160581 245762 226290
rect 246438 224501 246498 233139
rect 246435 224500 246501 224501
rect 246435 224436 246436 224500
rect 246500 224436 246501 224500
rect 246435 224435 246501 224436
rect 246806 218653 246866 239667
rect 248094 239461 248154 291755
rect 249379 289236 249445 289237
rect 249379 289172 249380 289236
rect 249444 289172 249445 289236
rect 249379 289171 249445 289172
rect 249195 240004 249261 240005
rect 249195 239940 249196 240004
rect 249260 239940 249261 240004
rect 249195 239939 249261 239940
rect 248275 239868 248341 239869
rect 248275 239804 248276 239868
rect 248340 239804 248341 239868
rect 248275 239803 248341 239804
rect 248643 239868 248709 239869
rect 248643 239804 248644 239868
rect 248708 239804 248709 239868
rect 248643 239803 248709 239804
rect 247539 239460 247605 239461
rect 247539 239396 247540 239460
rect 247604 239396 247605 239460
rect 247539 239395 247605 239396
rect 248091 239460 248157 239461
rect 248091 239396 248092 239460
rect 248156 239396 248157 239460
rect 248091 239395 248157 239396
rect 246987 226268 247053 226269
rect 246987 226204 246988 226268
rect 247052 226204 247053 226268
rect 246987 226203 247053 226204
rect 246990 224229 247050 226203
rect 246987 224228 247053 224229
rect 246987 224164 246988 224228
rect 247052 224164 247053 224228
rect 246987 224163 247053 224164
rect 247542 218925 247602 239395
rect 248278 226269 248338 239803
rect 248459 239732 248525 239733
rect 248459 239668 248460 239732
rect 248524 239668 248525 239732
rect 248459 239667 248525 239668
rect 248275 226268 248341 226269
rect 248275 226204 248276 226268
rect 248340 226204 248341 226268
rect 248275 226203 248341 226204
rect 248278 225997 248338 226203
rect 248275 225996 248341 225997
rect 248275 225932 248276 225996
rect 248340 225932 248341 225996
rect 248275 225931 248341 225932
rect 247539 218924 247605 218925
rect 247539 218860 247540 218924
rect 247604 218860 247605 218924
rect 247539 218859 247605 218860
rect 246803 218652 246869 218653
rect 246803 218588 246804 218652
rect 246868 218588 246869 218652
rect 246803 218587 246869 218588
rect 245699 160580 245765 160581
rect 245699 160516 245700 160580
rect 245764 160516 245765 160580
rect 245699 160515 245765 160516
rect 244779 157996 244845 157997
rect 244779 157932 244780 157996
rect 244844 157932 244845 157996
rect 244779 157931 244845 157932
rect 248462 143445 248522 239667
rect 248646 236469 248706 239803
rect 248643 236468 248709 236469
rect 248643 236404 248644 236468
rect 248708 236404 248709 236468
rect 248643 236403 248709 236404
rect 249198 227221 249258 239939
rect 249382 239869 249442 289171
rect 249379 239868 249445 239869
rect 249379 239804 249380 239868
rect 249444 239804 249445 239868
rect 249379 239803 249445 239804
rect 249566 239461 249626 312971
rect 252323 312900 252389 312901
rect 252323 312836 252324 312900
rect 252388 312836 252389 312900
rect 252323 312835 252389 312836
rect 251771 312764 251837 312765
rect 251771 312700 251772 312764
rect 251836 312700 251837 312764
rect 251771 312699 251837 312700
rect 250851 239868 250917 239869
rect 250851 239804 250852 239868
rect 250916 239804 250917 239868
rect 250851 239803 250917 239804
rect 250115 239732 250181 239733
rect 250115 239668 250116 239732
rect 250180 239668 250181 239732
rect 250115 239667 250181 239668
rect 249563 239460 249629 239461
rect 249563 239396 249564 239460
rect 249628 239396 249629 239460
rect 249563 239395 249629 239396
rect 249931 238780 249997 238781
rect 249931 238716 249932 238780
rect 249996 238716 249997 238780
rect 249931 238715 249997 238716
rect 249934 236741 249994 238715
rect 249931 236740 249997 236741
rect 249931 236676 249932 236740
rect 249996 236676 249997 236740
rect 249931 236675 249997 236676
rect 250118 234293 250178 239667
rect 250299 238644 250365 238645
rect 250299 238580 250300 238644
rect 250364 238580 250365 238644
rect 250299 238579 250365 238580
rect 250115 234292 250181 234293
rect 250115 234228 250116 234292
rect 250180 234228 250181 234292
rect 250115 234227 250181 234228
rect 249747 228308 249813 228309
rect 249747 228244 249748 228308
rect 249812 228244 249813 228308
rect 249747 228243 249813 228244
rect 249750 227357 249810 228243
rect 249747 227356 249813 227357
rect 249747 227292 249748 227356
rect 249812 227292 249813 227356
rect 249747 227291 249813 227292
rect 249195 227220 249261 227221
rect 249195 227156 249196 227220
rect 249260 227156 249261 227220
rect 249195 227155 249261 227156
rect 249198 226949 249258 227155
rect 249195 226948 249261 226949
rect 249195 226884 249196 226948
rect 249260 226884 249261 226948
rect 249195 226883 249261 226884
rect 250302 219333 250362 238579
rect 250854 228309 250914 239803
rect 251774 239733 251834 312699
rect 251955 293724 252021 293725
rect 251955 293660 251956 293724
rect 252020 293660 252021 293724
rect 251955 293659 252021 293660
rect 251958 239869 252018 293659
rect 251955 239868 252021 239869
rect 251955 239804 251956 239868
rect 252020 239804 252021 239868
rect 251955 239803 252021 239804
rect 251771 239732 251837 239733
rect 251771 239668 251772 239732
rect 251836 239668 251837 239732
rect 251771 239667 251837 239668
rect 251035 237828 251101 237829
rect 251035 237764 251036 237828
rect 251100 237764 251101 237828
rect 251035 237763 251101 237764
rect 250851 228308 250917 228309
rect 250851 228244 250852 228308
rect 250916 228244 250917 228308
rect 250851 228243 250917 228244
rect 251038 222189 251098 237763
rect 251774 233250 251834 239667
rect 252326 239461 252386 312835
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253059 291004 253125 291005
rect 253059 290940 253060 291004
rect 253124 290940 253125 291004
rect 253059 290939 253125 290940
rect 252691 241772 252757 241773
rect 252691 241708 252692 241772
rect 252756 241708 252757 241772
rect 252691 241707 252757 241708
rect 252694 239869 252754 241707
rect 252691 239868 252757 239869
rect 252691 239804 252692 239868
rect 252756 239804 252757 239868
rect 252691 239803 252757 239804
rect 253062 239461 253122 290939
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253243 290732 253309 290733
rect 253243 290668 253244 290732
rect 253308 290668 253309 290732
rect 253243 290667 253309 290668
rect 253246 239461 253306 290667
rect 253794 255454 254414 290898
rect 257514 705798 258134 705830
rect 257514 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 258134 705798
rect 257514 705478 258134 705562
rect 257514 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 258134 705478
rect 257514 691174 258134 705242
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 475174 258134 510618
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 439174 258134 474618
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 279923 452708 279989 452709
rect 279923 452644 279924 452708
rect 279988 452644 279989 452708
rect 279923 452643 279989 452644
rect 278635 451892 278701 451893
rect 278635 451828 278636 451892
rect 278700 451828 278701 451892
rect 278635 451827 278701 451828
rect 257514 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 258134 439174
rect 257514 438854 258134 438938
rect 257514 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 258134 438854
rect 257514 403174 258134 438618
rect 257514 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 258134 403174
rect 257514 402854 258134 402938
rect 257514 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 258134 402854
rect 257514 367174 258134 402618
rect 277899 375460 277965 375461
rect 277899 375396 277900 375460
rect 277964 375396 277965 375460
rect 277899 375395 277965 375396
rect 276611 371516 276677 371517
rect 276611 371452 276612 371516
rect 276676 371452 276677 371516
rect 276611 371451 276677 371452
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 257514 331174 258134 366618
rect 257514 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 258134 331174
rect 257514 330854 258134 330938
rect 257514 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 258134 330854
rect 257514 295174 258134 330618
rect 276614 323645 276674 371451
rect 276611 323644 276677 323645
rect 276611 323580 276612 323644
rect 276676 323580 276677 323644
rect 276611 323579 276677 323580
rect 274587 301340 274653 301341
rect 274587 301276 274588 301340
rect 274652 301276 274653 301340
rect 274587 301275 274653 301276
rect 257514 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 258134 295174
rect 257514 294854 258134 294938
rect 257514 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 258134 294854
rect 255635 267068 255701 267069
rect 255635 267004 255636 267068
rect 255700 267004 255701 267068
rect 255635 267003 255701 267004
rect 255451 258772 255517 258773
rect 255451 258708 255452 258772
rect 255516 258708 255517 258772
rect 255451 258707 255517 258708
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253427 239732 253493 239733
rect 253427 239668 253428 239732
rect 253492 239668 253493 239732
rect 253427 239667 253493 239668
rect 252323 239460 252389 239461
rect 252323 239396 252324 239460
rect 252388 239396 252389 239460
rect 252323 239395 252389 239396
rect 253059 239460 253125 239461
rect 253059 239396 253060 239460
rect 253124 239396 253125 239460
rect 253059 239395 253125 239396
rect 253243 239460 253309 239461
rect 253243 239396 253244 239460
rect 253308 239396 253309 239460
rect 253243 239395 253309 239396
rect 252326 233250 252386 239395
rect 252507 236740 252573 236741
rect 252507 236676 252508 236740
rect 252572 236676 252573 236740
rect 252507 236675 252573 236676
rect 251590 233190 251834 233250
rect 252142 233190 252386 233250
rect 251590 224365 251650 233190
rect 252142 232253 252202 233190
rect 252139 232252 252205 232253
rect 252139 232188 252140 232252
rect 252204 232188 252205 232252
rect 252139 232187 252205 232188
rect 252510 230077 252570 236675
rect 252875 236468 252941 236469
rect 252875 236404 252876 236468
rect 252940 236404 252941 236468
rect 252875 236403 252941 236404
rect 252507 230076 252573 230077
rect 252507 230012 252508 230076
rect 252572 230012 252573 230076
rect 252507 230011 252573 230012
rect 252878 228445 252938 236403
rect 253246 235789 253306 239395
rect 253243 235788 253309 235789
rect 253243 235724 253244 235788
rect 253308 235724 253309 235788
rect 253243 235723 253309 235724
rect 252875 228444 252941 228445
rect 252875 228380 252876 228444
rect 252940 228380 252941 228444
rect 252875 228379 252941 228380
rect 251587 224364 251653 224365
rect 251587 224300 251588 224364
rect 251652 224300 251653 224364
rect 251587 224299 251653 224300
rect 251035 222188 251101 222189
rect 251035 222124 251036 222188
rect 251100 222124 251101 222188
rect 251035 222123 251101 222124
rect 250299 219332 250365 219333
rect 250299 219268 250300 219332
rect 250364 219268 250365 219332
rect 250299 219267 250365 219268
rect 250302 218789 250362 219267
rect 253430 218925 253490 239667
rect 253794 219454 254414 254898
rect 254899 239868 254965 239869
rect 254899 239804 254900 239868
rect 254964 239804 254965 239868
rect 254899 239803 254965 239804
rect 254902 234429 254962 239803
rect 255454 239733 255514 258707
rect 255451 239732 255517 239733
rect 255451 239668 255452 239732
rect 255516 239668 255517 239732
rect 255451 239667 255517 239668
rect 255454 237965 255514 239667
rect 255638 238645 255698 267003
rect 257107 264484 257173 264485
rect 257107 264420 257108 264484
rect 257172 264420 257173 264484
rect 257107 264419 257173 264420
rect 256371 264212 256437 264213
rect 256371 264148 256372 264212
rect 256436 264148 256437 264212
rect 256371 264147 256437 264148
rect 256003 251836 256069 251837
rect 256003 251772 256004 251836
rect 256068 251772 256069 251836
rect 256003 251771 256069 251772
rect 256006 239869 256066 251771
rect 256003 239868 256069 239869
rect 256003 239804 256004 239868
rect 256068 239804 256069 239868
rect 256003 239803 256069 239804
rect 255635 238644 255701 238645
rect 255635 238580 255636 238644
rect 255700 238580 255701 238644
rect 255635 238579 255701 238580
rect 255451 237964 255517 237965
rect 255451 237900 255452 237964
rect 255516 237900 255517 237964
rect 255451 237899 255517 237900
rect 254899 234428 254965 234429
rect 254899 234364 254900 234428
rect 254964 234364 254965 234428
rect 254899 234363 254965 234364
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253427 218924 253493 218925
rect 253427 218860 253428 218924
rect 253492 218860 253493 218924
rect 253427 218859 253493 218860
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 250299 218788 250365 218789
rect 250299 218724 250300 218788
rect 250364 218724 250365 218788
rect 250299 218723 250365 218724
rect 253430 218109 253490 218859
rect 253427 218108 253493 218109
rect 253427 218044 253428 218108
rect 253492 218044 253493 218108
rect 253427 218043 253493 218044
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 248459 143444 248525 143445
rect 248459 143380 248460 143444
rect 248524 143380 248525 143444
rect 248459 143379 248525 143380
rect 242019 143172 242085 143173
rect 242019 143108 242020 143172
rect 242084 143108 242085 143172
rect 242019 143107 242085 143108
rect 240731 141948 240797 141949
rect 240731 141884 240732 141948
rect 240796 141884 240797 141948
rect 240731 141883 240797 141884
rect 238707 141812 238773 141813
rect 238707 141748 238708 141812
rect 238772 141748 238773 141812
rect 238707 141747 238773 141748
rect 221514 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 222134 115174
rect 221514 114854 222134 114938
rect 221514 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 222134 114854
rect 221514 79174 222134 114618
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -1306 222134 6618
rect 221514 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 222134 -1306
rect 221514 -1626 222134 -1542
rect 221514 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 222134 -1626
rect 221514 -1894 222134 -1862
rect 253794 111454 254414 146898
rect 254902 139093 254962 234363
rect 256006 233250 256066 239803
rect 256374 239461 256434 264147
rect 256923 244900 256989 244901
rect 256923 244836 256924 244900
rect 256988 244836 256989 244900
rect 256923 244835 256989 244836
rect 256371 239460 256437 239461
rect 256371 239396 256372 239460
rect 256436 239396 256437 239460
rect 256371 239395 256437 239396
rect 256926 238781 256986 244835
rect 257110 239733 257170 264419
rect 257514 259174 258134 294618
rect 262075 290596 262141 290597
rect 262075 290532 262076 290596
rect 262140 290532 262141 290596
rect 262075 290531 262141 290532
rect 260603 272508 260669 272509
rect 260603 272444 260604 272508
rect 260668 272444 260669 272508
rect 260603 272443 260669 272444
rect 259315 268428 259381 268429
rect 259315 268364 259316 268428
rect 259380 268364 259381 268428
rect 259315 268363 259381 268364
rect 259318 267750 259378 268363
rect 257514 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 258134 259174
rect 257514 258854 258134 258938
rect 257514 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 258134 258854
rect 257291 241636 257357 241637
rect 257291 241572 257292 241636
rect 257356 241572 257357 241636
rect 257291 241571 257357 241572
rect 257107 239732 257173 239733
rect 257107 239668 257108 239732
rect 257172 239668 257173 239732
rect 257107 239667 257173 239668
rect 257294 239461 257354 241571
rect 257291 239460 257357 239461
rect 257291 239396 257292 239460
rect 257356 239396 257357 239460
rect 257291 239395 257357 239396
rect 256923 238780 256989 238781
rect 256923 238716 256924 238780
rect 256988 238716 256989 238780
rect 256923 238715 256989 238716
rect 256371 236740 256437 236741
rect 256371 236676 256372 236740
rect 256436 236676 256437 236740
rect 256371 236675 256437 236676
rect 255822 233190 256066 233250
rect 255822 142901 255882 233190
rect 256374 222053 256434 236675
rect 256926 223590 256986 238715
rect 257107 235108 257173 235109
rect 257107 235044 257108 235108
rect 257172 235044 257173 235108
rect 257107 235043 257173 235044
rect 256742 223530 256986 223590
rect 256371 222052 256437 222053
rect 256371 221988 256372 222052
rect 256436 221988 256437 222052
rect 256371 221987 256437 221988
rect 256742 207637 256802 223530
rect 256739 207636 256805 207637
rect 256739 207572 256740 207636
rect 256804 207572 256805 207636
rect 256739 207571 256805 207572
rect 255819 142900 255885 142901
rect 255819 142836 255820 142900
rect 255884 142836 255885 142900
rect 255819 142835 255885 142836
rect 257110 139229 257170 235043
rect 257514 223174 258134 258618
rect 258766 267690 259378 267750
rect 258579 241500 258645 241501
rect 258579 241436 258580 241500
rect 258644 241436 258645 241500
rect 258579 241435 258645 241436
rect 258395 240684 258461 240685
rect 258395 240620 258396 240684
rect 258460 240620 258461 240684
rect 258395 240619 258461 240620
rect 258398 240277 258458 240619
rect 258395 240276 258461 240277
rect 258395 240212 258396 240276
rect 258460 240212 258461 240276
rect 258395 240211 258461 240212
rect 258395 240004 258461 240005
rect 258395 239940 258396 240004
rect 258460 239940 258461 240004
rect 258395 239939 258461 239940
rect 258398 238373 258458 239939
rect 258582 239461 258642 241435
rect 258579 239460 258645 239461
rect 258579 239396 258580 239460
rect 258644 239396 258645 239460
rect 258579 239395 258645 239396
rect 258395 238372 258461 238373
rect 258395 238308 258396 238372
rect 258460 238308 258461 238372
rect 258395 238307 258461 238308
rect 258582 236741 258642 239395
rect 258766 238101 258826 267690
rect 259131 262852 259197 262853
rect 259131 262788 259132 262852
rect 259196 262788 259197 262852
rect 259131 262787 259197 262788
rect 258947 248028 259013 248029
rect 258947 247964 258948 248028
rect 259012 247964 259013 248028
rect 258947 247963 259013 247964
rect 258950 238237 259010 247963
rect 259134 239461 259194 262787
rect 260419 257276 260485 257277
rect 260419 257212 260420 257276
rect 260484 257212 260485 257276
rect 260419 257211 260485 257212
rect 259499 242180 259565 242181
rect 259499 242116 259500 242180
rect 259564 242116 259565 242180
rect 259499 242115 259565 242116
rect 259502 239733 259562 242115
rect 259867 240684 259933 240685
rect 259867 240620 259868 240684
rect 259932 240620 259933 240684
rect 259867 240619 259933 240620
rect 259499 239732 259565 239733
rect 259499 239668 259500 239732
rect 259564 239668 259565 239732
rect 259499 239667 259565 239668
rect 259683 239732 259749 239733
rect 259683 239668 259684 239732
rect 259748 239668 259749 239732
rect 259683 239667 259749 239668
rect 259131 239460 259197 239461
rect 259131 239396 259132 239460
rect 259196 239396 259197 239460
rect 259131 239395 259197 239396
rect 259315 239460 259381 239461
rect 259315 239396 259316 239460
rect 259380 239396 259381 239460
rect 259315 239395 259381 239396
rect 259318 238509 259378 239395
rect 259499 238780 259565 238781
rect 259499 238716 259500 238780
rect 259564 238716 259565 238780
rect 259499 238715 259565 238716
rect 259315 238508 259381 238509
rect 259315 238444 259316 238508
rect 259380 238444 259381 238508
rect 259315 238443 259381 238444
rect 258947 238236 259013 238237
rect 258947 238172 258948 238236
rect 259012 238172 259013 238236
rect 258947 238171 259013 238172
rect 258763 238100 258829 238101
rect 258763 238036 258764 238100
rect 258828 238036 258829 238100
rect 258763 238035 258829 238036
rect 258579 236740 258645 236741
rect 258579 236676 258580 236740
rect 258644 236676 258645 236740
rect 258579 236675 258645 236676
rect 258579 233340 258645 233341
rect 258579 233276 258580 233340
rect 258644 233276 258645 233340
rect 258579 233275 258645 233276
rect 258582 227629 258642 233275
rect 259502 232389 259562 238715
rect 259499 232388 259565 232389
rect 259499 232324 259500 232388
rect 259564 232324 259565 232388
rect 259499 232323 259565 232324
rect 258579 227628 258645 227629
rect 258579 227564 258580 227628
rect 258644 227564 258645 227628
rect 258579 227563 258645 227564
rect 257514 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 258134 223174
rect 257514 222854 258134 222938
rect 257514 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 258134 222854
rect 257514 187174 258134 222618
rect 257514 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 258134 187174
rect 257514 186854 258134 186938
rect 257514 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 258134 186854
rect 257514 151174 258134 186618
rect 258582 152965 258642 227563
rect 258579 152964 258645 152965
rect 258579 152900 258580 152964
rect 258644 152900 258645 152964
rect 258579 152899 258645 152900
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 257107 139228 257173 139229
rect 257107 139164 257108 139228
rect 257172 139164 257173 139228
rect 257107 139163 257173 139164
rect 254899 139092 254965 139093
rect 254899 139028 254900 139092
rect 254964 139028 254965 139092
rect 254899 139027 254965 139028
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 115174 258134 150618
rect 259686 144397 259746 239667
rect 259870 238373 259930 240619
rect 260422 239733 260482 257211
rect 260419 239732 260485 239733
rect 260419 239668 260420 239732
rect 260484 239668 260485 239732
rect 260419 239667 260485 239668
rect 260606 238781 260666 272443
rect 261891 261492 261957 261493
rect 261891 261428 261892 261492
rect 261956 261428 261957 261492
rect 261891 261427 261957 261428
rect 261707 253196 261773 253197
rect 261707 253132 261708 253196
rect 261772 253132 261773 253196
rect 261707 253131 261773 253132
rect 261710 247050 261770 253131
rect 261158 246990 261770 247050
rect 261158 239461 261218 246990
rect 261894 240002 261954 261427
rect 261526 239942 261954 240002
rect 261526 239733 261586 239942
rect 261707 239868 261773 239869
rect 261707 239804 261708 239868
rect 261772 239804 261773 239868
rect 261707 239803 261773 239804
rect 261523 239732 261589 239733
rect 261523 239668 261524 239732
rect 261588 239668 261589 239732
rect 261523 239667 261589 239668
rect 261155 239460 261221 239461
rect 261155 239396 261156 239460
rect 261220 239396 261221 239460
rect 261155 239395 261221 239396
rect 261158 239050 261218 239395
rect 260974 238990 261218 239050
rect 260419 238780 260485 238781
rect 260419 238716 260420 238780
rect 260484 238716 260485 238780
rect 260419 238715 260485 238716
rect 260603 238780 260669 238781
rect 260603 238716 260604 238780
rect 260668 238716 260669 238780
rect 260603 238715 260669 238716
rect 259867 238372 259933 238373
rect 259867 238308 259868 238372
rect 259932 238308 259933 238372
rect 259867 238307 259933 238308
rect 260422 226269 260482 238715
rect 260606 238373 260666 238715
rect 260603 238372 260669 238373
rect 260603 238308 260604 238372
rect 260668 238308 260669 238372
rect 260603 238307 260669 238308
rect 260419 226268 260485 226269
rect 260419 226204 260420 226268
rect 260484 226204 260485 226268
rect 260419 226203 260485 226204
rect 260974 221509 261034 238990
rect 261339 236196 261405 236197
rect 261339 236132 261340 236196
rect 261404 236132 261405 236196
rect 261339 236131 261405 236132
rect 261155 234564 261221 234565
rect 261155 234500 261156 234564
rect 261220 234500 261221 234564
rect 261155 234499 261221 234500
rect 260971 221508 261037 221509
rect 260971 221444 260972 221508
rect 261036 221444 261037 221508
rect 260971 221443 261037 221444
rect 261158 145893 261218 234499
rect 261342 224773 261402 236131
rect 261526 235109 261586 239667
rect 261710 235653 261770 239803
rect 262078 239733 262138 290531
rect 269619 287740 269685 287741
rect 269619 287676 269620 287740
rect 269684 287676 269685 287740
rect 269619 287675 269685 287676
rect 266675 271148 266741 271149
rect 266675 271084 266676 271148
rect 266740 271084 266741 271148
rect 266675 271083 266741 271084
rect 264835 264348 264901 264349
rect 264835 264284 264836 264348
rect 264900 264284 264901 264348
rect 264835 264283 264901 264284
rect 263547 258908 263613 258909
rect 263547 258844 263548 258908
rect 263612 258844 263613 258908
rect 263547 258843 263613 258844
rect 263550 251190 263610 258843
rect 263550 251130 263978 251190
rect 263547 250612 263613 250613
rect 263547 250548 263548 250612
rect 263612 250548 263613 250612
rect 263547 250547 263613 250548
rect 263550 249810 263610 250547
rect 263550 249750 263794 249810
rect 263363 247756 263429 247757
rect 263363 247692 263364 247756
rect 263428 247692 263429 247756
rect 263363 247691 263429 247692
rect 262443 239868 262509 239869
rect 262443 239804 262444 239868
rect 262508 239804 262509 239868
rect 262443 239803 262509 239804
rect 262995 239868 263061 239869
rect 262995 239804 262996 239868
rect 263060 239804 263061 239868
rect 262995 239803 263061 239804
rect 262075 239732 262141 239733
rect 262075 239668 262076 239732
rect 262140 239668 262141 239732
rect 262075 239667 262141 239668
rect 262259 239732 262325 239733
rect 262259 239668 262260 239732
rect 262324 239668 262325 239732
rect 262259 239667 262325 239668
rect 261707 235652 261773 235653
rect 261707 235588 261708 235652
rect 261772 235588 261773 235652
rect 261707 235587 261773 235588
rect 261523 235108 261589 235109
rect 261523 235044 261524 235108
rect 261588 235044 261589 235108
rect 261523 235043 261589 235044
rect 261339 224772 261405 224773
rect 261339 224708 261340 224772
rect 261404 224708 261405 224772
rect 261339 224707 261405 224708
rect 261155 145892 261221 145893
rect 261155 145828 261156 145892
rect 261220 145828 261221 145892
rect 261155 145827 261221 145828
rect 259683 144396 259749 144397
rect 259683 144332 259684 144396
rect 259748 144332 259749 144396
rect 259683 144331 259749 144332
rect 261342 143853 261402 224707
rect 262262 146029 262322 239667
rect 262446 232253 262506 239803
rect 262811 237964 262877 237965
rect 262811 237900 262812 237964
rect 262876 237900 262877 237964
rect 262811 237899 262877 237900
rect 262443 232252 262509 232253
rect 262443 232188 262444 232252
rect 262508 232188 262509 232252
rect 262443 232187 262509 232188
rect 262446 229805 262506 232187
rect 262814 230213 262874 237899
rect 262998 230893 263058 239803
rect 263366 239733 263426 247691
rect 263547 239868 263613 239869
rect 263547 239804 263548 239868
rect 263612 239804 263613 239868
rect 263547 239803 263613 239804
rect 263363 239732 263429 239733
rect 263363 239668 263364 239732
rect 263428 239668 263429 239732
rect 263363 239667 263429 239668
rect 263363 239460 263429 239461
rect 263363 239396 263364 239460
rect 263428 239396 263429 239460
rect 263363 239395 263429 239396
rect 263179 237692 263245 237693
rect 263179 237628 263180 237692
rect 263244 237628 263245 237692
rect 263179 237627 263245 237628
rect 262995 230892 263061 230893
rect 262995 230828 262996 230892
rect 263060 230828 263061 230892
rect 262995 230827 263061 230828
rect 262811 230212 262877 230213
rect 262811 230148 262812 230212
rect 262876 230148 262877 230212
rect 262811 230147 262877 230148
rect 262443 229804 262509 229805
rect 262443 229740 262444 229804
rect 262508 229740 262509 229804
rect 262443 229739 262509 229740
rect 263182 223549 263242 237627
rect 263179 223548 263245 223549
rect 263179 223484 263180 223548
rect 263244 223484 263245 223548
rect 263179 223483 263245 223484
rect 263366 221781 263426 239395
rect 263550 238237 263610 239803
rect 263734 239461 263794 249750
rect 263918 239869 263978 251130
rect 264283 245036 264349 245037
rect 264283 244972 264284 245036
rect 264348 244972 264349 245036
rect 264283 244971 264349 244972
rect 263915 239868 263981 239869
rect 263915 239804 263916 239868
rect 263980 239804 263981 239868
rect 263915 239803 263981 239804
rect 264099 239732 264165 239733
rect 264099 239730 264100 239732
rect 263918 239670 264100 239730
rect 263731 239460 263797 239461
rect 263731 239396 263732 239460
rect 263796 239396 263797 239460
rect 263731 239395 263797 239396
rect 263547 238236 263613 238237
rect 263547 238172 263548 238236
rect 263612 238172 263613 238236
rect 263547 238171 263613 238172
rect 263363 221780 263429 221781
rect 263363 221716 263364 221780
rect 263428 221716 263429 221780
rect 263363 221715 263429 221716
rect 263366 219450 263426 221715
rect 262814 219390 263426 219450
rect 262814 146301 262874 219390
rect 263918 169013 263978 239670
rect 264099 239668 264100 239670
rect 264164 239668 264165 239732
rect 264099 239667 264165 239668
rect 264099 238780 264165 238781
rect 264099 238716 264100 238780
rect 264164 238778 264165 238780
rect 264286 238778 264346 244971
rect 264838 239869 264898 264283
rect 266123 255916 266189 255917
rect 266123 255852 266124 255916
rect 266188 255852 266189 255916
rect 266123 255851 266189 255852
rect 266126 251190 266186 255851
rect 265758 251130 266186 251190
rect 265387 246668 265453 246669
rect 265387 246604 265388 246668
rect 265452 246604 265453 246668
rect 265387 246603 265453 246604
rect 265203 240412 265269 240413
rect 265203 240348 265204 240412
rect 265268 240348 265269 240412
rect 265203 240347 265269 240348
rect 264835 239868 264901 239869
rect 264835 239804 264836 239868
rect 264900 239804 264901 239868
rect 264835 239803 264901 239804
rect 265206 239733 265266 240347
rect 265390 239869 265450 246603
rect 265387 239868 265453 239869
rect 265387 239804 265388 239868
rect 265452 239804 265453 239868
rect 265387 239803 265453 239804
rect 265203 239732 265269 239733
rect 265203 239668 265204 239732
rect 265268 239668 265269 239732
rect 265203 239667 265269 239668
rect 265390 238781 265450 239803
rect 265758 239733 265818 251130
rect 266123 249116 266189 249117
rect 266123 249052 266124 249116
rect 266188 249052 266189 249116
rect 266123 249051 266189 249052
rect 266126 248430 266186 249051
rect 266126 248370 266370 248430
rect 266123 246260 266189 246261
rect 266123 246196 266124 246260
rect 266188 246196 266189 246260
rect 266123 246195 266189 246196
rect 266126 239733 266186 246195
rect 266310 239869 266370 248370
rect 266307 239868 266373 239869
rect 266307 239804 266308 239868
rect 266372 239804 266373 239868
rect 266307 239803 266373 239804
rect 266678 239733 266738 271083
rect 267411 253332 267477 253333
rect 267411 253268 267412 253332
rect 267476 253268 267477 253332
rect 267411 253267 267477 253268
rect 267414 242317 267474 253267
rect 267411 242316 267477 242317
rect 267411 242252 267412 242316
rect 267476 242252 267477 242316
rect 267411 242251 267477 242252
rect 269622 241637 269682 287675
rect 271091 273868 271157 273869
rect 271091 273804 271092 273868
rect 271156 273804 271157 273868
rect 271091 273803 271157 273804
rect 269619 241636 269685 241637
rect 269619 241572 269620 241636
rect 269684 241572 269685 241636
rect 269619 241571 269685 241572
rect 265755 239732 265821 239733
rect 265755 239668 265756 239732
rect 265820 239668 265821 239732
rect 265755 239667 265821 239668
rect 266123 239732 266189 239733
rect 266123 239668 266124 239732
rect 266188 239668 266189 239732
rect 266123 239667 266189 239668
rect 266675 239732 266741 239733
rect 266675 239668 266676 239732
rect 266740 239668 266741 239732
rect 266675 239667 266741 239668
rect 264164 238718 264346 238778
rect 265387 238780 265453 238781
rect 264164 238716 264165 238718
rect 264099 238715 264165 238716
rect 265387 238716 265388 238780
rect 265452 238716 265453 238780
rect 265387 238715 265453 238716
rect 264102 221373 264162 238715
rect 265755 237148 265821 237149
rect 265755 237084 265756 237148
rect 265820 237084 265821 237148
rect 265755 237083 265821 237084
rect 265758 232661 265818 237083
rect 266126 236741 266186 239667
rect 268331 237964 268397 237965
rect 268331 237900 268332 237964
rect 268396 237900 268397 237964
rect 268331 237899 268397 237900
rect 268334 237149 268394 237899
rect 271094 237693 271154 273803
rect 274590 240685 274650 301275
rect 277902 291957 277962 375395
rect 278451 373012 278517 373013
rect 278451 372948 278452 373012
rect 278516 372948 278517 373012
rect 278451 372947 278517 372948
rect 278454 358869 278514 372947
rect 278638 369205 278698 451827
rect 279371 371652 279437 371653
rect 279371 371588 279372 371652
rect 279436 371588 279437 371652
rect 279371 371587 279437 371588
rect 278635 369204 278701 369205
rect 278635 369140 278636 369204
rect 278700 369140 278701 369204
rect 278635 369139 278701 369140
rect 278451 358868 278517 358869
rect 278451 358804 278452 358868
rect 278516 358804 278517 358868
rect 278451 358803 278517 358804
rect 279374 321197 279434 371587
rect 279926 369341 279986 452643
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 287651 398988 287717 398989
rect 287651 398924 287652 398988
rect 287716 398924 287717 398988
rect 287651 398923 287717 398924
rect 283419 395996 283485 395997
rect 283419 395932 283420 395996
rect 283484 395932 283485 395996
rect 283419 395931 283485 395932
rect 282315 371924 282381 371925
rect 282315 371860 282316 371924
rect 282380 371860 282381 371924
rect 282315 371859 282381 371860
rect 281027 371788 281093 371789
rect 281027 371724 281028 371788
rect 281092 371724 281093 371788
rect 281027 371723 281093 371724
rect 280843 371652 280909 371653
rect 280843 371588 280844 371652
rect 280908 371588 280909 371652
rect 280843 371587 280909 371588
rect 280659 370292 280725 370293
rect 280659 370228 280660 370292
rect 280724 370228 280725 370292
rect 280659 370227 280725 370228
rect 279923 369340 279989 369341
rect 279923 369276 279924 369340
rect 279988 369276 279989 369340
rect 279923 369275 279989 369276
rect 279371 321196 279437 321197
rect 279371 321132 279372 321196
rect 279436 321132 279437 321196
rect 279371 321131 279437 321132
rect 280662 292365 280722 370227
rect 280846 362269 280906 371587
rect 281030 363629 281090 371723
rect 282131 369884 282197 369885
rect 282131 369820 282132 369884
rect 282196 369820 282197 369884
rect 282131 369819 282197 369820
rect 281395 369204 281461 369205
rect 281395 369140 281396 369204
rect 281460 369140 281461 369204
rect 281395 369139 281461 369140
rect 281027 363628 281093 363629
rect 281027 363564 281028 363628
rect 281092 363564 281093 363628
rect 281027 363563 281093 363564
rect 280843 362268 280909 362269
rect 280843 362204 280844 362268
rect 280908 362204 280909 362268
rect 280843 362203 280909 362204
rect 280659 292364 280725 292365
rect 280659 292300 280660 292364
rect 280724 292300 280725 292364
rect 280659 292299 280725 292300
rect 277899 291956 277965 291957
rect 277899 291892 277900 291956
rect 277964 291892 277965 291956
rect 277899 291891 277965 291892
rect 274587 240684 274653 240685
rect 274587 240620 274588 240684
rect 274652 240620 274653 240684
rect 274587 240619 274653 240620
rect 271827 238780 271893 238781
rect 271827 238716 271828 238780
rect 271892 238716 271893 238780
rect 271827 238715 271893 238716
rect 271091 237692 271157 237693
rect 271091 237628 271092 237692
rect 271156 237628 271157 237692
rect 271091 237627 271157 237628
rect 268331 237148 268397 237149
rect 268331 237084 268332 237148
rect 268396 237084 268397 237148
rect 268331 237083 268397 237084
rect 266123 236740 266189 236741
rect 266123 236676 266124 236740
rect 266188 236676 266189 236740
rect 266123 236675 266189 236676
rect 265755 232660 265821 232661
rect 265755 232596 265756 232660
rect 265820 232596 265821 232660
rect 265755 232595 265821 232596
rect 264099 221372 264165 221373
rect 264099 221308 264100 221372
rect 264164 221308 264165 221372
rect 264099 221307 264165 221308
rect 265758 219450 265818 232595
rect 265574 219390 265818 219450
rect 263915 169012 263981 169013
rect 263915 168948 263916 169012
rect 263980 168948 263981 169012
rect 263915 168947 263981 168948
rect 265574 147661 265634 219390
rect 265571 147660 265637 147661
rect 265571 147596 265572 147660
rect 265636 147596 265637 147660
rect 265571 147595 265637 147596
rect 262811 146300 262877 146301
rect 262811 146236 262812 146300
rect 262876 146236 262877 146300
rect 262811 146235 262877 146236
rect 262259 146028 262325 146029
rect 262259 145964 262260 146028
rect 262324 145964 262325 146028
rect 262259 145963 262325 145964
rect 261339 143852 261405 143853
rect 261339 143788 261340 143852
rect 261404 143788 261405 143852
rect 261339 143787 261405 143788
rect 268334 141813 268394 237083
rect 268331 141812 268397 141813
rect 268331 141748 268332 141812
rect 268396 141748 268397 141812
rect 268331 141747 268397 141748
rect 271830 138005 271890 238715
rect 274590 235925 274650 240619
rect 274587 235924 274653 235925
rect 274587 235860 274588 235924
rect 274652 235860 274653 235924
rect 274587 235859 274653 235860
rect 271827 138004 271893 138005
rect 271827 137940 271828 138004
rect 271892 137940 271893 138004
rect 271827 137939 271893 137940
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 257514 79174 258134 114618
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 281398 71909 281458 369139
rect 282134 292501 282194 369819
rect 282318 358053 282378 371859
rect 282315 358052 282381 358053
rect 282315 357988 282316 358052
rect 282380 357988 282381 358052
rect 282315 357987 282381 357988
rect 283422 320517 283482 395931
rect 283603 395180 283669 395181
rect 283603 395116 283604 395180
rect 283668 395116 283669 395180
rect 283603 395115 283669 395116
rect 283606 320653 283666 395115
rect 286915 394364 286981 394365
rect 286915 394300 286916 394364
rect 286980 394300 286981 394364
rect 286915 394299 286981 394300
rect 285075 391916 285141 391917
rect 285075 391852 285076 391916
rect 285140 391852 285141 391916
rect 285075 391851 285141 391852
rect 283787 387428 283853 387429
rect 283787 387364 283788 387428
rect 283852 387364 283853 387428
rect 283787 387363 283853 387364
rect 283790 320789 283850 387363
rect 283971 377636 284037 377637
rect 283971 377572 283972 377636
rect 284036 377572 284037 377636
rect 283971 377571 284037 377572
rect 283974 321605 284034 377571
rect 283971 321604 284037 321605
rect 283971 321540 283972 321604
rect 284036 321540 284037 321604
rect 283971 321539 284037 321540
rect 283974 320789 284034 321539
rect 283787 320788 283853 320789
rect 283787 320724 283788 320788
rect 283852 320724 283853 320788
rect 283787 320723 283853 320724
rect 283971 320788 284037 320789
rect 283971 320724 283972 320788
rect 284036 320724 284037 320788
rect 283971 320723 284037 320724
rect 283603 320652 283669 320653
rect 283603 320588 283604 320652
rect 283668 320588 283669 320652
rect 283603 320587 283669 320588
rect 283419 320516 283485 320517
rect 283419 320452 283420 320516
rect 283484 320452 283485 320516
rect 283419 320451 283485 320452
rect 283422 318613 283482 320451
rect 283606 319429 283666 320587
rect 283603 319428 283669 319429
rect 283603 319364 283604 319428
rect 283668 319364 283669 319428
rect 283603 319363 283669 319364
rect 283790 318749 283850 320723
rect 283971 320652 284037 320653
rect 283971 320588 283972 320652
rect 284036 320588 284037 320652
rect 283971 320587 284037 320588
rect 283974 320381 284034 320587
rect 285078 320381 285138 391851
rect 286363 388924 286429 388925
rect 286363 388860 286364 388924
rect 286428 388860 286429 388924
rect 286363 388859 286429 388860
rect 285443 387020 285509 387021
rect 285443 386956 285444 387020
rect 285508 386956 285509 387020
rect 285443 386955 285509 386956
rect 285259 381852 285325 381853
rect 285259 381788 285260 381852
rect 285324 381788 285325 381852
rect 285259 381787 285325 381788
rect 285262 320517 285322 381787
rect 285259 320516 285325 320517
rect 285259 320452 285260 320516
rect 285324 320452 285325 320516
rect 285259 320451 285325 320452
rect 283971 320380 284037 320381
rect 283971 320316 283972 320380
rect 284036 320316 284037 320380
rect 283971 320315 284037 320316
rect 284339 320380 284405 320381
rect 284339 320316 284340 320380
rect 284404 320316 284405 320380
rect 284339 320315 284405 320316
rect 285075 320380 285141 320381
rect 285075 320316 285076 320380
rect 285140 320316 285141 320380
rect 285075 320315 285141 320316
rect 283971 320108 284037 320109
rect 283971 320044 283972 320108
rect 284036 320044 284037 320108
rect 283971 320043 284037 320044
rect 283974 318885 284034 320043
rect 283971 318884 284037 318885
rect 283971 318820 283972 318884
rect 284036 318820 284037 318884
rect 283971 318819 284037 318820
rect 283787 318748 283853 318749
rect 283787 318684 283788 318748
rect 283852 318684 283853 318748
rect 283787 318683 283853 318684
rect 283419 318612 283485 318613
rect 283419 318548 283420 318612
rect 283484 318548 283485 318612
rect 283419 318547 283485 318548
rect 284342 318477 284402 320315
rect 284891 320108 284957 320109
rect 284891 320044 284892 320108
rect 284956 320044 284957 320108
rect 284891 320043 284957 320044
rect 284339 318476 284405 318477
rect 284339 318412 284340 318476
rect 284404 318412 284405 318476
rect 284339 318411 284405 318412
rect 283235 317796 283301 317797
rect 283235 317732 283236 317796
rect 283300 317732 283301 317796
rect 283235 317731 283301 317732
rect 283051 317524 283117 317525
rect 283051 317460 283052 317524
rect 283116 317460 283117 317524
rect 283051 317459 283117 317460
rect 282867 311948 282933 311949
rect 282867 311884 282868 311948
rect 282932 311884 282933 311948
rect 282867 311883 282933 311884
rect 282870 304877 282930 311883
rect 283054 307597 283114 317459
rect 283238 311949 283298 317731
rect 283235 311948 283301 311949
rect 283235 311884 283236 311948
rect 283300 311884 283301 311948
rect 284894 311910 284954 320043
rect 285078 318810 285138 320315
rect 285446 320109 285506 386955
rect 285627 369612 285693 369613
rect 285627 369548 285628 369612
rect 285692 369548 285693 369612
rect 285627 369547 285693 369548
rect 285630 368797 285690 369547
rect 285627 368796 285693 368797
rect 285627 368732 285628 368796
rect 285692 368732 285693 368796
rect 285627 368731 285693 368732
rect 286366 325710 286426 388859
rect 286547 385796 286613 385797
rect 286547 385732 286548 385796
rect 286612 385732 286613 385796
rect 286547 385731 286613 385732
rect 285998 325650 286426 325710
rect 285998 321570 286058 325650
rect 285630 321510 286058 321570
rect 285630 320109 285690 321510
rect 286363 320652 286429 320653
rect 286363 320588 286364 320652
rect 286428 320588 286429 320652
rect 286363 320587 286429 320588
rect 285811 320516 285877 320517
rect 285811 320452 285812 320516
rect 285876 320452 285877 320516
rect 285811 320451 285877 320452
rect 285443 320108 285509 320109
rect 285443 320044 285444 320108
rect 285508 320044 285509 320108
rect 285443 320043 285509 320044
rect 285627 320108 285693 320109
rect 285627 320044 285628 320108
rect 285692 320044 285693 320108
rect 285627 320043 285693 320044
rect 285078 318750 285506 318810
rect 285446 318341 285506 318750
rect 285443 318340 285509 318341
rect 285443 318276 285444 318340
rect 285508 318276 285509 318340
rect 285443 318275 285509 318276
rect 283235 311883 283301 311884
rect 284342 311850 284954 311910
rect 283051 307596 283117 307597
rect 283051 307532 283052 307596
rect 283116 307532 283117 307596
rect 283051 307531 283117 307532
rect 282867 304876 282933 304877
rect 282867 304812 282868 304876
rect 282932 304812 282933 304876
rect 282867 304811 282933 304812
rect 284342 296445 284402 311850
rect 284339 296444 284405 296445
rect 284339 296380 284340 296444
rect 284404 296380 284405 296444
rect 284339 296379 284405 296380
rect 285630 294677 285690 320043
rect 285814 294813 285874 320451
rect 286366 319701 286426 320587
rect 286550 320381 286610 385731
rect 286918 320517 286978 394299
rect 287283 369612 287349 369613
rect 287283 369548 287284 369612
rect 287348 369548 287349 369612
rect 287283 369547 287349 369548
rect 287286 369341 287346 369547
rect 287283 369340 287349 369341
rect 287283 369276 287284 369340
rect 287348 369276 287349 369340
rect 287283 369275 287349 369276
rect 287286 368661 287346 369275
rect 287283 368660 287349 368661
rect 287283 368596 287284 368660
rect 287348 368596 287349 368660
rect 287283 368595 287349 368596
rect 287099 320924 287165 320925
rect 287099 320860 287100 320924
rect 287164 320860 287165 320924
rect 287099 320859 287165 320860
rect 286915 320516 286981 320517
rect 286915 320452 286916 320516
rect 286980 320452 286981 320516
rect 286915 320451 286981 320452
rect 286547 320380 286613 320381
rect 286547 320316 286548 320380
rect 286612 320316 286613 320380
rect 286547 320315 286613 320316
rect 286363 319700 286429 319701
rect 286363 319636 286364 319700
rect 286428 319636 286429 319700
rect 286363 319635 286429 319636
rect 286363 309772 286429 309773
rect 286363 309708 286364 309772
rect 286428 309770 286429 309772
rect 286550 309770 286610 320315
rect 287102 320109 287162 320859
rect 287467 320380 287533 320381
rect 287467 320316 287468 320380
rect 287532 320316 287533 320380
rect 287467 320315 287533 320316
rect 287099 320108 287165 320109
rect 287099 320044 287100 320108
rect 287164 320044 287165 320108
rect 287099 320043 287165 320044
rect 287470 319293 287530 320315
rect 287467 319292 287533 319293
rect 287467 319228 287468 319292
rect 287532 319228 287533 319292
rect 287467 319227 287533 319228
rect 287654 318749 287714 398923
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 288939 391100 289005 391101
rect 288939 391036 288940 391100
rect 289004 391036 289005 391100
rect 288939 391035 289005 391036
rect 288203 388788 288269 388789
rect 288203 388724 288204 388788
rect 288268 388724 288269 388788
rect 288203 388723 288269 388724
rect 288206 320789 288266 388723
rect 288203 320788 288269 320789
rect 288203 320724 288204 320788
rect 288268 320724 288269 320788
rect 288203 320723 288269 320724
rect 287651 318748 287717 318749
rect 287651 318684 287652 318748
rect 287716 318684 287717 318748
rect 287651 318683 287717 318684
rect 287651 310996 287717 310997
rect 287651 310932 287652 310996
rect 287716 310932 287717 310996
rect 287651 310931 287717 310932
rect 286428 309710 286610 309770
rect 286428 309708 286429 309710
rect 286363 309707 286429 309708
rect 285811 294812 285877 294813
rect 285811 294748 285812 294812
rect 285876 294748 285877 294812
rect 285811 294747 285877 294748
rect 285627 294676 285693 294677
rect 285627 294612 285628 294676
rect 285692 294612 285693 294676
rect 285627 294611 285693 294612
rect 282131 292500 282197 292501
rect 282131 292436 282132 292500
rect 282196 292436 282197 292500
rect 282131 292435 282197 292436
rect 287654 237421 287714 310931
rect 288206 310045 288266 320723
rect 288387 320516 288453 320517
rect 288387 320452 288388 320516
rect 288452 320514 288453 320516
rect 288452 320454 288634 320514
rect 288452 320452 288453 320454
rect 288387 320451 288453 320452
rect 288387 320380 288453 320381
rect 288387 320316 288388 320380
rect 288452 320316 288453 320380
rect 288387 320315 288453 320316
rect 288203 310044 288269 310045
rect 288203 309980 288204 310044
rect 288268 309980 288269 310044
rect 288203 309979 288269 309980
rect 288390 294269 288450 320315
rect 288574 319293 288634 320454
rect 288755 320108 288821 320109
rect 288755 320044 288756 320108
rect 288820 320044 288821 320108
rect 288755 320043 288821 320044
rect 288571 319292 288637 319293
rect 288571 319228 288572 319292
rect 288636 319228 288637 319292
rect 288571 319227 288637 319228
rect 288758 319157 288818 320043
rect 288755 319156 288821 319157
rect 288755 319092 288756 319156
rect 288820 319092 288821 319156
rect 288755 319091 288821 319092
rect 288942 318613 289002 391035
rect 289491 388652 289557 388653
rect 289491 388588 289492 388652
rect 289556 388588 289557 388652
rect 289491 388587 289557 388588
rect 289307 378860 289373 378861
rect 289307 378796 289308 378860
rect 289372 378796 289373 378860
rect 289307 378795 289373 378796
rect 289123 378724 289189 378725
rect 289123 378660 289124 378724
rect 289188 378660 289189 378724
rect 289123 378659 289189 378660
rect 289126 320109 289186 378659
rect 289123 320108 289189 320109
rect 289123 320044 289124 320108
rect 289188 320044 289189 320108
rect 289123 320043 289189 320044
rect 288939 318612 289005 318613
rect 288939 318548 288940 318612
rect 289004 318548 289005 318612
rect 288939 318547 289005 318548
rect 289126 307461 289186 320043
rect 289310 318341 289370 378795
rect 289494 320381 289554 388587
rect 289794 363454 290414 398898
rect 293514 705798 294134 705830
rect 293514 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 294134 705798
rect 293514 705478 294134 705562
rect 293514 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 294134 705478
rect 293514 691174 294134 705242
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 475174 294134 510618
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 439174 294134 474618
rect 293514 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 294134 439174
rect 293514 438854 294134 438938
rect 293514 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 294134 438854
rect 293514 403174 294134 438618
rect 293514 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 294134 403174
rect 293514 402854 294134 402938
rect 293514 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 294134 402854
rect 293171 398852 293237 398853
rect 293171 398788 293172 398852
rect 293236 398788 293237 398852
rect 293171 398787 293237 398788
rect 292987 392324 293053 392325
rect 292987 392260 292988 392324
rect 293052 392260 293053 392324
rect 292987 392259 293053 392260
rect 292803 391508 292869 391509
rect 292803 391444 292804 391508
rect 292868 391444 292869 391508
rect 292803 391443 292869 391444
rect 290963 381716 291029 381717
rect 290963 381652 290964 381716
rect 291028 381652 291029 381716
rect 290963 381651 291029 381652
rect 290779 379404 290845 379405
rect 290779 379340 290780 379404
rect 290844 379340 290845 379404
rect 290779 379339 290845 379340
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289491 320380 289557 320381
rect 289491 320316 289492 320380
rect 289556 320316 289557 320380
rect 289491 320315 289557 320316
rect 289307 318340 289373 318341
rect 289307 318276 289308 318340
rect 289372 318276 289373 318340
rect 289307 318275 289373 318276
rect 289123 307460 289189 307461
rect 289123 307396 289124 307460
rect 289188 307396 289189 307460
rect 289123 307395 289189 307396
rect 288387 294268 288453 294269
rect 288387 294204 288388 294268
rect 288452 294204 288453 294268
rect 288387 294203 288453 294204
rect 289794 291454 290414 326898
rect 290782 320381 290842 379339
rect 290966 320789 291026 381651
rect 291883 379268 291949 379269
rect 291883 379204 291884 379268
rect 291948 379204 291949 379268
rect 291883 379203 291949 379204
rect 291699 373420 291765 373421
rect 291699 373356 291700 373420
rect 291764 373356 291765 373420
rect 291699 373355 291765 373356
rect 291702 320789 291762 373355
rect 290963 320788 291029 320789
rect 290963 320724 290964 320788
rect 291028 320724 291029 320788
rect 290963 320723 291029 320724
rect 291699 320788 291765 320789
rect 291699 320724 291700 320788
rect 291764 320724 291765 320788
rect 291699 320723 291765 320724
rect 290779 320380 290845 320381
rect 290779 320316 290780 320380
rect 290844 320316 290845 320380
rect 290779 320315 290845 320316
rect 290595 320108 290661 320109
rect 290595 320044 290596 320108
rect 290660 320044 290661 320108
rect 290595 320043 290661 320044
rect 290598 318885 290658 320043
rect 290595 318884 290661 318885
rect 290595 318820 290596 318884
rect 290660 318820 290661 318884
rect 290595 318819 290661 318820
rect 290782 311133 290842 320315
rect 290779 311132 290845 311133
rect 290779 311068 290780 311132
rect 290844 311068 290845 311132
rect 290779 311067 290845 311068
rect 290966 296730 291026 320723
rect 291147 319700 291213 319701
rect 291147 319636 291148 319700
rect 291212 319636 291213 319700
rect 291147 319635 291213 319636
rect 291150 318885 291210 319635
rect 291702 319157 291762 320723
rect 291886 320109 291946 379203
rect 292251 379132 292317 379133
rect 292251 379068 292252 379132
rect 292316 379068 292317 379132
rect 292251 379067 292317 379068
rect 292067 377364 292133 377365
rect 292067 377300 292068 377364
rect 292132 377300 292133 377364
rect 292067 377299 292133 377300
rect 292070 320789 292130 377299
rect 292067 320788 292133 320789
rect 292067 320724 292068 320788
rect 292132 320724 292133 320788
rect 292067 320723 292133 320724
rect 292067 320516 292133 320517
rect 292067 320452 292068 320516
rect 292132 320452 292133 320516
rect 292067 320451 292133 320452
rect 291883 320108 291949 320109
rect 291883 320044 291884 320108
rect 291948 320044 291949 320108
rect 291883 320043 291949 320044
rect 291699 319156 291765 319157
rect 291699 319092 291700 319156
rect 291764 319092 291765 319156
rect 291699 319091 291765 319092
rect 291147 318884 291213 318885
rect 291147 318820 291148 318884
rect 291212 318820 291213 318884
rect 291147 318819 291213 318820
rect 291331 318068 291397 318069
rect 291331 318004 291332 318068
rect 291396 318004 291397 318068
rect 291331 318003 291397 318004
rect 291147 317796 291213 317797
rect 291147 317732 291148 317796
rect 291212 317732 291213 317796
rect 291147 317731 291213 317732
rect 291150 311677 291210 317731
rect 291334 315757 291394 318003
rect 291331 315756 291397 315757
rect 291331 315692 291332 315756
rect 291396 315692 291397 315756
rect 291331 315691 291397 315692
rect 291147 311676 291213 311677
rect 291147 311612 291148 311676
rect 291212 311612 291213 311676
rect 291147 311611 291213 311612
rect 291886 311405 291946 320043
rect 292070 318205 292130 320451
rect 292254 320381 292314 379067
rect 292435 320788 292501 320789
rect 292435 320724 292436 320788
rect 292500 320724 292501 320788
rect 292435 320723 292501 320724
rect 292251 320380 292317 320381
rect 292251 320316 292252 320380
rect 292316 320316 292317 320380
rect 292251 320315 292317 320316
rect 292067 318204 292133 318205
rect 292067 318140 292068 318204
rect 292132 318140 292133 318204
rect 292067 318139 292133 318140
rect 291883 311404 291949 311405
rect 291883 311340 291884 311404
rect 291948 311340 291949 311404
rect 291883 311339 291949 311340
rect 292254 311269 292314 320315
rect 292438 319293 292498 320723
rect 292806 320517 292866 391443
rect 292803 320516 292869 320517
rect 292803 320452 292804 320516
rect 292868 320452 292869 320516
rect 292803 320451 292869 320452
rect 292619 320380 292685 320381
rect 292619 320316 292620 320380
rect 292684 320316 292685 320380
rect 292619 320315 292685 320316
rect 292435 319292 292501 319293
rect 292435 319228 292436 319292
rect 292500 319228 292501 319292
rect 292435 319227 292501 319228
rect 292622 312629 292682 320315
rect 292990 320245 293050 392259
rect 292803 320244 292869 320245
rect 292803 320180 292804 320244
rect 292868 320180 292869 320244
rect 292803 320179 292869 320180
rect 292987 320244 293053 320245
rect 292987 320180 292988 320244
rect 293052 320180 293053 320244
rect 292987 320179 293053 320180
rect 292806 319565 292866 320179
rect 292803 319564 292869 319565
rect 292803 319500 292804 319564
rect 292868 319500 292869 319564
rect 292803 319499 292869 319500
rect 292990 313989 293050 320179
rect 293174 320109 293234 398787
rect 293514 367174 294134 402618
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 318563 397084 318629 397085
rect 318563 397020 318564 397084
rect 318628 397020 318629 397084
rect 318563 397019 318629 397020
rect 315803 396948 315869 396949
rect 315803 396884 315804 396948
rect 315868 396884 315869 396948
rect 315803 396883 315869 396884
rect 313043 395996 313109 395997
rect 313043 395932 313044 395996
rect 313108 395932 313109 395996
rect 313043 395931 313109 395932
rect 295563 394500 295629 394501
rect 295563 394436 295564 394500
rect 295628 394436 295629 394500
rect 295563 394435 295629 394436
rect 295195 391780 295261 391781
rect 295195 391716 295196 391780
rect 295260 391716 295261 391780
rect 295195 391715 295261 391716
rect 295011 391644 295077 391645
rect 295011 391580 295012 391644
rect 295076 391580 295077 391644
rect 295011 391579 295077 391580
rect 294643 390284 294709 390285
rect 294643 390220 294644 390284
rect 294708 390220 294709 390284
rect 294643 390219 294709 390220
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 293514 331174 294134 366618
rect 293514 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 294134 331174
rect 293514 330854 294134 330938
rect 293514 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 294134 330854
rect 293355 320516 293421 320517
rect 293355 320452 293356 320516
rect 293420 320452 293421 320516
rect 293355 320451 293421 320452
rect 293171 320108 293237 320109
rect 293171 320044 293172 320108
rect 293236 320044 293237 320108
rect 293171 320043 293237 320044
rect 292987 313988 293053 313989
rect 292987 313924 292988 313988
rect 293052 313924 293053 313988
rect 292987 313923 293053 313924
rect 292619 312628 292685 312629
rect 292619 312564 292620 312628
rect 292684 312564 292685 312628
rect 292619 312563 292685 312564
rect 292251 311268 292317 311269
rect 292251 311204 292252 311268
rect 292316 311204 292317 311268
rect 292251 311203 292317 311204
rect 293174 296730 293234 320043
rect 293358 312357 293418 320451
rect 293355 312356 293421 312357
rect 293355 312292 293356 312356
rect 293420 312292 293421 312356
rect 293355 312291 293421 312292
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 287651 237420 287717 237421
rect 287651 237356 287652 237420
rect 287716 237356 287717 237420
rect 287651 237355 287717 237356
rect 289794 219454 290414 254898
rect 290598 296670 291026 296730
rect 292622 296670 293234 296730
rect 290598 220421 290658 296670
rect 292622 241093 292682 296670
rect 293514 295174 294134 330618
rect 294459 321332 294525 321333
rect 294459 321268 294460 321332
rect 294524 321268 294525 321332
rect 294459 321267 294525 321268
rect 294275 321196 294341 321197
rect 294275 321132 294276 321196
rect 294340 321132 294341 321196
rect 294275 321131 294341 321132
rect 294278 320517 294338 321131
rect 294275 320516 294341 320517
rect 294275 320452 294276 320516
rect 294340 320452 294341 320516
rect 294275 320451 294341 320452
rect 294462 320381 294522 321267
rect 294646 320517 294706 390219
rect 294827 389740 294893 389741
rect 294827 389676 294828 389740
rect 294892 389676 294893 389740
rect 294827 389675 294893 389676
rect 294643 320516 294709 320517
rect 294643 320452 294644 320516
rect 294708 320452 294709 320516
rect 294643 320451 294709 320452
rect 294459 320380 294525 320381
rect 294459 320316 294460 320380
rect 294524 320316 294525 320380
rect 294459 320315 294525 320316
rect 294459 320108 294525 320109
rect 294459 320044 294460 320108
rect 294524 320044 294525 320108
rect 294459 320043 294525 320044
rect 294462 318477 294522 320043
rect 294459 318476 294525 318477
rect 294459 318412 294460 318476
rect 294524 318412 294525 318476
rect 294459 318411 294525 318412
rect 294646 313290 294706 320451
rect 294830 320245 294890 389675
rect 294827 320244 294893 320245
rect 294827 320180 294828 320244
rect 294892 320180 294893 320244
rect 294827 320179 294893 320180
rect 293514 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 294134 295174
rect 293514 294854 294134 294938
rect 293514 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 294134 294854
rect 293514 259174 294134 294618
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 292619 241092 292685 241093
rect 292619 241028 292620 241092
rect 292684 241028 292685 241092
rect 292619 241027 292685 241028
rect 293514 223174 294134 258618
rect 294462 313230 294706 313290
rect 294462 240821 294522 313230
rect 294830 308413 294890 320179
rect 295014 319973 295074 391579
rect 295198 321197 295258 391715
rect 295195 321196 295261 321197
rect 295195 321132 295196 321196
rect 295260 321132 295261 321196
rect 295195 321131 295261 321132
rect 295566 320653 295626 394435
rect 296115 394228 296181 394229
rect 296115 394164 296116 394228
rect 296180 394164 296181 394228
rect 296115 394163 296181 394164
rect 295931 384436 295997 384437
rect 295931 384372 295932 384436
rect 295996 384372 295997 384436
rect 295931 384371 295997 384372
rect 295934 320789 295994 384371
rect 295931 320788 295997 320789
rect 295931 320724 295932 320788
rect 295996 320724 295997 320788
rect 295931 320723 295997 320724
rect 295563 320652 295629 320653
rect 295563 320588 295564 320652
rect 295628 320588 295629 320652
rect 295563 320587 295629 320588
rect 295747 320244 295813 320245
rect 295747 320180 295748 320244
rect 295812 320180 295813 320244
rect 295747 320179 295813 320180
rect 295195 320108 295261 320109
rect 295195 320044 295196 320108
rect 295260 320044 295261 320108
rect 295195 320043 295261 320044
rect 295011 319972 295077 319973
rect 295011 319908 295012 319972
rect 295076 319908 295077 319972
rect 295011 319907 295077 319908
rect 294827 308412 294893 308413
rect 294827 308348 294828 308412
rect 294892 308348 294893 308412
rect 294827 308347 294893 308348
rect 295014 298757 295074 319907
rect 295198 316029 295258 320043
rect 295195 316028 295261 316029
rect 295195 315964 295196 316028
rect 295260 315964 295261 316028
rect 295195 315963 295261 315964
rect 295750 314941 295810 320179
rect 295934 317525 295994 320723
rect 296118 319837 296178 394163
rect 297955 393820 298021 393821
rect 297955 393756 297956 393820
rect 298020 393756 298021 393820
rect 297955 393755 298021 393756
rect 296483 393684 296549 393685
rect 296483 393620 296484 393684
rect 296548 393620 296549 393684
rect 296483 393619 296549 393620
rect 296299 320788 296365 320789
rect 296299 320724 296300 320788
rect 296364 320724 296365 320788
rect 296299 320723 296365 320724
rect 296115 319836 296181 319837
rect 296115 319772 296116 319836
rect 296180 319772 296181 319836
rect 296115 319771 296181 319772
rect 295931 317524 295997 317525
rect 295931 317460 295932 317524
rect 295996 317460 295997 317524
rect 295931 317459 295997 317460
rect 296118 315485 296178 319771
rect 296302 318810 296362 320723
rect 296486 320245 296546 393619
rect 297035 392868 297101 392869
rect 297035 392804 297036 392868
rect 297100 392804 297101 392868
rect 297035 392803 297101 392804
rect 297038 321570 297098 392803
rect 297587 387292 297653 387293
rect 297587 387228 297588 387292
rect 297652 387228 297653 387292
rect 297587 387227 297653 387228
rect 297403 380220 297469 380221
rect 297403 380156 297404 380220
rect 297468 380156 297469 380220
rect 297403 380155 297469 380156
rect 297406 325710 297466 380155
rect 296854 321510 297098 321570
rect 297222 325650 297466 325710
rect 296667 320788 296733 320789
rect 296667 320724 296668 320788
rect 296732 320724 296733 320788
rect 296667 320723 296733 320724
rect 296483 320244 296549 320245
rect 296483 320180 296484 320244
rect 296548 320180 296549 320244
rect 296483 320179 296549 320180
rect 296302 318750 296546 318810
rect 296486 315893 296546 318750
rect 296483 315892 296549 315893
rect 296483 315828 296484 315892
rect 296548 315828 296549 315892
rect 296483 315827 296549 315828
rect 296115 315484 296181 315485
rect 296115 315420 296116 315484
rect 296180 315420 296181 315484
rect 296115 315419 296181 315420
rect 295931 315348 295997 315349
rect 295931 315284 295932 315348
rect 295996 315284 295997 315348
rect 295931 315283 295997 315284
rect 295747 314940 295813 314941
rect 295747 314876 295748 314940
rect 295812 314876 295813 314940
rect 295747 314875 295813 314876
rect 295011 298756 295077 298757
rect 295011 298692 295012 298756
rect 295076 298692 295077 298756
rect 295011 298691 295077 298692
rect 294459 240820 294525 240821
rect 294459 240756 294460 240820
rect 294524 240756 294525 240820
rect 294459 240755 294525 240756
rect 295934 231573 295994 315283
rect 296670 311910 296730 320723
rect 296854 320517 296914 321510
rect 296851 320516 296917 320517
rect 296851 320452 296852 320516
rect 296916 320452 296917 320516
rect 297222 320514 297282 325650
rect 296851 320451 296917 320452
rect 297038 320454 297282 320514
rect 296854 315757 296914 320451
rect 297038 320245 297098 320454
rect 297035 320244 297101 320245
rect 297035 320180 297036 320244
rect 297100 320180 297101 320244
rect 297035 320179 297101 320180
rect 296851 315756 296917 315757
rect 296851 315692 296852 315756
rect 296916 315692 296917 315756
rect 296851 315691 296917 315692
rect 297038 315621 297098 320179
rect 297590 320109 297650 387227
rect 297958 320789 298018 393755
rect 302187 393140 302253 393141
rect 302187 393076 302188 393140
rect 302252 393076 302253 393140
rect 302187 393075 302253 393076
rect 302003 393004 302069 393005
rect 302003 392940 302004 393004
rect 302068 392940 302069 393004
rect 302003 392939 302069 392940
rect 298507 392460 298573 392461
rect 298507 392396 298508 392460
rect 298572 392396 298573 392460
rect 298507 392395 298573 392396
rect 298510 320789 298570 392395
rect 299979 381580 300045 381581
rect 299979 381516 299980 381580
rect 300044 381516 300045 381580
rect 299979 381515 300045 381516
rect 299982 321570 300042 381515
rect 301451 369476 301517 369477
rect 301451 369412 301452 369476
rect 301516 369412 301517 369476
rect 301451 369411 301517 369412
rect 301454 321570 301514 369411
rect 299430 321510 300042 321570
rect 301270 321510 301514 321570
rect 297955 320788 298021 320789
rect 297955 320724 297956 320788
rect 298020 320724 298021 320788
rect 297955 320723 298021 320724
rect 298507 320788 298573 320789
rect 298507 320724 298508 320788
rect 298572 320724 298573 320788
rect 298507 320723 298573 320724
rect 299059 320788 299125 320789
rect 299059 320724 299060 320788
rect 299124 320724 299125 320788
rect 299059 320723 299125 320724
rect 298323 320516 298389 320517
rect 298323 320452 298324 320516
rect 298388 320452 298389 320516
rect 298323 320451 298389 320452
rect 297587 320108 297653 320109
rect 297587 320044 297588 320108
rect 297652 320044 297653 320108
rect 297587 320043 297653 320044
rect 297955 319972 298021 319973
rect 297955 319908 297956 319972
rect 298020 319908 298021 319972
rect 297955 319907 298021 319908
rect 297587 319836 297653 319837
rect 297587 319772 297588 319836
rect 297652 319772 297653 319836
rect 297587 319771 297653 319772
rect 297035 315620 297101 315621
rect 297035 315556 297036 315620
rect 297100 315556 297101 315620
rect 297035 315555 297101 315556
rect 296486 311850 296730 311910
rect 296486 307733 296546 311850
rect 296483 307732 296549 307733
rect 296483 307668 296484 307732
rect 296548 307668 296549 307732
rect 296483 307667 296549 307668
rect 297590 307325 297650 319771
rect 297958 316709 298018 319907
rect 298326 319293 298386 320451
rect 298510 319701 298570 320723
rect 298875 320516 298941 320517
rect 298875 320452 298876 320516
rect 298940 320452 298941 320516
rect 298875 320451 298941 320452
rect 298507 319700 298573 319701
rect 298507 319636 298508 319700
rect 298572 319636 298573 319700
rect 298507 319635 298573 319636
rect 298323 319292 298389 319293
rect 298323 319228 298324 319292
rect 298388 319228 298389 319292
rect 298323 319227 298389 319228
rect 298691 319292 298757 319293
rect 298691 319228 298692 319292
rect 298756 319228 298757 319292
rect 298691 319227 298757 319228
rect 298139 317932 298205 317933
rect 298139 317868 298140 317932
rect 298204 317868 298205 317932
rect 298139 317867 298205 317868
rect 297955 316708 298021 316709
rect 297955 316644 297956 316708
rect 298020 316644 298021 316708
rect 297955 316643 298021 316644
rect 297587 307324 297653 307325
rect 297587 307260 297588 307324
rect 297652 307260 297653 307324
rect 297587 307259 297653 307260
rect 298142 300117 298202 317867
rect 298694 310453 298754 319227
rect 298878 314261 298938 320451
rect 299062 319701 299122 320723
rect 299430 320245 299490 321510
rect 299427 320244 299493 320245
rect 299427 320180 299428 320244
rect 299492 320180 299493 320244
rect 299427 320179 299493 320180
rect 300899 320244 300965 320245
rect 300899 320180 300900 320244
rect 300964 320180 300965 320244
rect 300899 320179 300965 320180
rect 299243 320108 299309 320109
rect 299243 320044 299244 320108
rect 299308 320044 299309 320108
rect 299243 320043 299309 320044
rect 299059 319700 299125 319701
rect 299059 319636 299060 319700
rect 299124 319636 299125 319700
rect 299059 319635 299125 319636
rect 299246 315077 299306 320043
rect 299430 318069 299490 320179
rect 299795 320108 299861 320109
rect 299795 320044 299796 320108
rect 299860 320044 299861 320108
rect 299795 320043 299861 320044
rect 299427 318068 299493 318069
rect 299427 318004 299428 318068
rect 299492 318004 299493 318068
rect 299427 318003 299493 318004
rect 299611 317932 299677 317933
rect 299611 317868 299612 317932
rect 299676 317868 299677 317932
rect 299611 317867 299677 317868
rect 299427 317524 299493 317525
rect 299427 317460 299428 317524
rect 299492 317460 299493 317524
rect 299427 317459 299493 317460
rect 299243 315076 299309 315077
rect 299243 315012 299244 315076
rect 299308 315012 299309 315076
rect 299243 315011 299309 315012
rect 298875 314260 298941 314261
rect 298875 314196 298876 314260
rect 298940 314196 298941 314260
rect 298875 314195 298941 314196
rect 299430 313853 299490 317459
rect 299427 313852 299493 313853
rect 299427 313788 299428 313852
rect 299492 313788 299493 313852
rect 299427 313787 299493 313788
rect 299614 313581 299674 317867
rect 299611 313580 299677 313581
rect 299611 313516 299612 313580
rect 299676 313516 299677 313580
rect 299611 313515 299677 313516
rect 299798 312629 299858 320043
rect 299795 312628 299861 312629
rect 299795 312564 299796 312628
rect 299860 312564 299861 312628
rect 299795 312563 299861 312564
rect 298691 310452 298757 310453
rect 298691 310388 298692 310452
rect 298756 310388 298757 310452
rect 298691 310387 298757 310388
rect 299979 308412 300045 308413
rect 299979 308348 299980 308412
rect 300044 308348 300045 308412
rect 299979 308347 300045 308348
rect 298139 300116 298205 300117
rect 298139 300052 298140 300116
rect 298204 300052 298205 300116
rect 298139 300051 298205 300052
rect 299982 232797 300042 308347
rect 299979 232796 300045 232797
rect 299979 232732 299980 232796
rect 300044 232732 300045 232796
rect 299979 232731 300045 232732
rect 295931 231572 295997 231573
rect 295931 231508 295932 231572
rect 295996 231508 295997 231572
rect 295931 231507 295997 231508
rect 300902 223277 300962 320179
rect 301270 320109 301330 321510
rect 301451 321196 301517 321197
rect 301451 321132 301452 321196
rect 301516 321132 301517 321196
rect 301451 321131 301517 321132
rect 301267 320108 301333 320109
rect 301267 320044 301268 320108
rect 301332 320044 301333 320108
rect 301267 320043 301333 320044
rect 301083 317524 301149 317525
rect 301083 317460 301084 317524
rect 301148 317460 301149 317524
rect 301083 317459 301149 317460
rect 301086 303517 301146 317459
rect 301270 307053 301330 320043
rect 301454 313581 301514 321131
rect 302006 320245 302066 392939
rect 302190 379530 302250 393075
rect 310283 391916 310349 391917
rect 310283 391852 310284 391916
rect 310348 391852 310349 391916
rect 310283 391851 310349 391852
rect 307707 390692 307773 390693
rect 307707 390628 307708 390692
rect 307772 390628 307773 390692
rect 307707 390627 307773 390628
rect 304947 383212 305013 383213
rect 304947 383148 304948 383212
rect 305012 383148 305013 383212
rect 304947 383147 305013 383148
rect 302190 379470 302434 379530
rect 302374 360770 302434 379470
rect 302739 369476 302805 369477
rect 302739 369412 302740 369476
rect 302804 369412 302805 369476
rect 302739 369411 302805 369412
rect 302190 360710 302434 360770
rect 302190 321330 302250 360710
rect 302742 360210 302802 369411
rect 302374 360150 302802 360210
rect 302374 328470 302434 360150
rect 304950 345030 305010 383147
rect 306971 378996 307037 378997
rect 306971 378932 306972 378996
rect 307036 378932 307037 378996
rect 306971 378931 307037 378932
rect 306235 373556 306301 373557
rect 306235 373492 306236 373556
rect 306300 373492 306301 373556
rect 306235 373491 306301 373492
rect 304950 344970 305378 345030
rect 302374 328410 302618 328470
rect 302190 321270 302434 321330
rect 302187 320516 302253 320517
rect 302187 320452 302188 320516
rect 302252 320452 302253 320516
rect 302187 320451 302253 320452
rect 302190 320245 302250 320451
rect 302003 320244 302069 320245
rect 302003 320180 302004 320244
rect 302068 320180 302069 320244
rect 302003 320179 302069 320180
rect 302187 320244 302253 320245
rect 302187 320180 302188 320244
rect 302252 320180 302253 320244
rect 302187 320179 302253 320180
rect 302374 320109 302434 321270
rect 302558 320789 302618 328410
rect 305318 325710 305378 344970
rect 306238 325710 306298 373491
rect 305318 325650 305562 325710
rect 303291 321060 303357 321061
rect 303291 320996 303292 321060
rect 303356 320996 303357 321060
rect 303291 320995 303357 320996
rect 302555 320788 302621 320789
rect 302555 320724 302556 320788
rect 302620 320724 302621 320788
rect 302555 320723 302621 320724
rect 302371 320108 302437 320109
rect 302371 320044 302372 320108
rect 302436 320044 302437 320108
rect 302371 320043 302437 320044
rect 301635 319972 301701 319973
rect 301635 319908 301636 319972
rect 301700 319908 301701 319972
rect 301635 319907 301701 319908
rect 301638 315757 301698 319907
rect 302374 319429 302434 320043
rect 302371 319428 302437 319429
rect 302371 319364 302372 319428
rect 302436 319364 302437 319428
rect 302371 319363 302437 319364
rect 302371 318748 302437 318749
rect 302371 318684 302372 318748
rect 302436 318684 302437 318748
rect 302371 318683 302437 318684
rect 301635 315756 301701 315757
rect 301635 315692 301636 315756
rect 301700 315692 301701 315756
rect 301635 315691 301701 315692
rect 301451 313580 301517 313581
rect 301451 313516 301452 313580
rect 301516 313516 301517 313580
rect 301451 313515 301517 313516
rect 302374 311910 302434 318683
rect 302558 318613 302618 320723
rect 303294 319701 303354 320995
rect 305315 320516 305381 320517
rect 305315 320452 305316 320516
rect 305380 320452 305381 320516
rect 305315 320451 305381 320452
rect 303291 319700 303357 319701
rect 303291 319636 303292 319700
rect 303356 319636 303357 319700
rect 303291 319635 303357 319636
rect 304211 318884 304277 318885
rect 304211 318820 304212 318884
rect 304276 318820 304277 318884
rect 304211 318819 304277 318820
rect 302555 318612 302621 318613
rect 302555 318548 302556 318612
rect 302620 318548 302621 318612
rect 302555 318547 302621 318548
rect 303475 318068 303541 318069
rect 303475 318004 303476 318068
rect 303540 318004 303541 318068
rect 303475 318003 303541 318004
rect 302739 317932 302805 317933
rect 302739 317868 302740 317932
rect 302804 317868 302805 317932
rect 302739 317867 302805 317868
rect 302190 311850 302434 311910
rect 301267 307052 301333 307053
rect 301267 306988 301268 307052
rect 301332 306988 301333 307052
rect 301267 306987 301333 306988
rect 301083 303516 301149 303517
rect 301083 303452 301084 303516
rect 301148 303452 301149 303516
rect 301083 303451 301149 303452
rect 302190 300253 302250 311850
rect 302555 302292 302621 302293
rect 302555 302228 302556 302292
rect 302620 302228 302621 302292
rect 302555 302227 302621 302228
rect 302187 300252 302253 300253
rect 302187 300188 302188 300252
rect 302252 300188 302253 300252
rect 302187 300187 302253 300188
rect 302558 226133 302618 302227
rect 302742 297669 302802 317867
rect 302923 317524 302989 317525
rect 302923 317460 302924 317524
rect 302988 317460 302989 317524
rect 302923 317459 302989 317460
rect 302926 303517 302986 317459
rect 303478 308685 303538 318003
rect 303475 308684 303541 308685
rect 303475 308620 303476 308684
rect 303540 308620 303541 308684
rect 303475 308619 303541 308620
rect 302923 303516 302989 303517
rect 302923 303452 302924 303516
rect 302988 303452 302989 303516
rect 302923 303451 302989 303452
rect 302926 302293 302986 303451
rect 302923 302292 302989 302293
rect 302923 302228 302924 302292
rect 302988 302228 302989 302292
rect 302923 302227 302989 302228
rect 302739 297668 302805 297669
rect 302739 297604 302740 297668
rect 302804 297604 302805 297668
rect 302739 297603 302805 297604
rect 302742 293589 302802 297603
rect 302739 293588 302805 293589
rect 302739 293524 302740 293588
rect 302804 293524 302805 293588
rect 302739 293523 302805 293524
rect 302555 226132 302621 226133
rect 302555 226068 302556 226132
rect 302620 226068 302621 226132
rect 302555 226067 302621 226068
rect 304214 224637 304274 318819
rect 304579 317932 304645 317933
rect 304579 317868 304580 317932
rect 304644 317868 304645 317932
rect 304579 317867 304645 317868
rect 304395 317524 304461 317525
rect 304395 317460 304396 317524
rect 304460 317460 304461 317524
rect 304395 317459 304461 317460
rect 304398 298077 304458 317459
rect 304582 304741 304642 317867
rect 305318 314125 305378 320451
rect 305502 320109 305562 325650
rect 306054 325650 306298 325710
rect 306054 320517 306114 325650
rect 306974 321197 307034 378931
rect 307523 373284 307589 373285
rect 307523 373220 307524 373284
rect 307588 373220 307589 373284
rect 307523 373219 307589 373220
rect 306971 321196 307037 321197
rect 306971 321132 306972 321196
rect 307036 321132 307037 321196
rect 306971 321131 307037 321132
rect 306974 320789 307034 321131
rect 306971 320788 307037 320789
rect 306971 320724 306972 320788
rect 307036 320724 307037 320788
rect 306971 320723 307037 320724
rect 306051 320516 306117 320517
rect 306051 320452 306052 320516
rect 306116 320452 306117 320516
rect 306051 320451 306117 320452
rect 307526 320109 307586 373219
rect 307710 325710 307770 390627
rect 308995 377500 309061 377501
rect 308995 377436 308996 377500
rect 309060 377436 309061 377500
rect 308995 377435 309061 377436
rect 307710 325650 307954 325710
rect 307894 321570 307954 325650
rect 308811 321876 308877 321877
rect 308811 321812 308812 321876
rect 308876 321812 308877 321876
rect 308811 321811 308877 321812
rect 307710 321510 307954 321570
rect 307710 320517 307770 321510
rect 308814 320789 308874 321811
rect 308811 320788 308877 320789
rect 308811 320724 308812 320788
rect 308876 320724 308877 320788
rect 308811 320723 308877 320724
rect 307707 320516 307773 320517
rect 307707 320452 307708 320516
rect 307772 320452 307773 320516
rect 307707 320451 307773 320452
rect 307710 320245 307770 320451
rect 307707 320244 307773 320245
rect 307707 320180 307708 320244
rect 307772 320180 307773 320244
rect 307707 320179 307773 320180
rect 308998 320109 309058 377435
rect 310099 369340 310165 369341
rect 310099 369276 310100 369340
rect 310164 369276 310165 369340
rect 310099 369275 310165 369276
rect 310102 368389 310162 369275
rect 310099 368388 310165 368389
rect 310099 368324 310100 368388
rect 310164 368324 310165 368388
rect 310099 368323 310165 368324
rect 310286 321570 310346 391851
rect 311019 369612 311085 369613
rect 311019 369548 311020 369612
rect 311084 369548 311085 369612
rect 311019 369547 311085 369548
rect 310102 321510 310346 321570
rect 309547 320380 309613 320381
rect 309547 320316 309548 320380
rect 309612 320316 309613 320380
rect 309547 320315 309613 320316
rect 309915 320380 309981 320381
rect 309915 320316 309916 320380
rect 309980 320316 309981 320380
rect 309915 320315 309981 320316
rect 305499 320108 305565 320109
rect 305499 320044 305500 320108
rect 305564 320044 305565 320108
rect 305499 320043 305565 320044
rect 307523 320108 307589 320109
rect 307523 320044 307524 320108
rect 307588 320044 307589 320108
rect 307523 320043 307589 320044
rect 307707 320108 307773 320109
rect 307707 320044 307708 320108
rect 307772 320044 307773 320108
rect 307707 320043 307773 320044
rect 308995 320108 309061 320109
rect 308995 320044 308996 320108
rect 309060 320044 309061 320108
rect 308995 320043 309061 320044
rect 305502 318885 305562 320043
rect 305683 319972 305749 319973
rect 305683 319908 305684 319972
rect 305748 319908 305749 319972
rect 305683 319907 305749 319908
rect 305499 318884 305565 318885
rect 305499 318820 305500 318884
rect 305564 318820 305565 318884
rect 305499 318819 305565 318820
rect 305315 314124 305381 314125
rect 305315 314060 305316 314124
rect 305380 314060 305381 314124
rect 305315 314059 305381 314060
rect 305686 311910 305746 319907
rect 306419 318340 306485 318341
rect 306419 318276 306420 318340
rect 306484 318276 306485 318340
rect 306419 318275 306485 318276
rect 305502 311850 305746 311910
rect 304579 304740 304645 304741
rect 304579 304676 304580 304740
rect 304644 304676 304645 304740
rect 304579 304675 304645 304676
rect 305502 302021 305562 311850
rect 304947 302020 305013 302021
rect 304947 301956 304948 302020
rect 305012 301956 305013 302020
rect 304947 301955 305013 301956
rect 305499 302020 305565 302021
rect 305499 301956 305500 302020
rect 305564 301956 305565 302020
rect 305499 301955 305565 301956
rect 304950 301613 305010 301955
rect 304947 301612 305013 301613
rect 304947 301548 304948 301612
rect 305012 301548 305013 301612
rect 304947 301547 305013 301548
rect 304395 298076 304461 298077
rect 304395 298012 304396 298076
rect 304460 298012 304461 298076
rect 304395 298011 304461 298012
rect 306422 225997 306482 318275
rect 306971 317932 307037 317933
rect 306971 317868 306972 317932
rect 307036 317868 307037 317932
rect 306971 317867 307037 317868
rect 306974 316981 307034 317867
rect 307523 317524 307589 317525
rect 307523 317460 307524 317524
rect 307588 317460 307589 317524
rect 307523 317459 307589 317460
rect 306971 316980 307037 316981
rect 306971 316916 306972 316980
rect 307036 316916 307037 316980
rect 306971 316915 307037 316916
rect 306419 225996 306485 225997
rect 306419 225932 306420 225996
rect 306484 225932 306485 225996
rect 306419 225931 306485 225932
rect 304211 224636 304277 224637
rect 304211 224572 304212 224636
rect 304276 224572 304277 224636
rect 304211 224571 304277 224572
rect 300899 223276 300965 223277
rect 300899 223212 300900 223276
rect 300964 223212 300965 223276
rect 300899 223211 300965 223212
rect 293514 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 294134 223174
rect 293514 222854 294134 222938
rect 293514 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 294134 222854
rect 290595 220420 290661 220421
rect 290595 220356 290596 220420
rect 290660 220356 290661 220420
rect 290595 220355 290661 220356
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 281395 71908 281461 71909
rect 281395 71844 281396 71908
rect 281460 71844 281461 71908
rect 281395 71843 281461 71844
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -1306 258134 6618
rect 257514 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 258134 -1306
rect 257514 -1626 258134 -1542
rect 257514 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 258134 -1626
rect 257514 -1894 258134 -1862
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 187174 294134 222618
rect 306974 219061 307034 316915
rect 307526 314669 307586 317459
rect 307523 314668 307589 314669
rect 307523 314604 307524 314668
rect 307588 314604 307589 314668
rect 307523 314603 307589 314604
rect 307710 228581 307770 320043
rect 309550 319701 309610 320315
rect 309547 319700 309613 319701
rect 309547 319636 309548 319700
rect 309612 319636 309613 319700
rect 309547 319635 309613 319636
rect 309918 319565 309978 320315
rect 309915 319564 309981 319565
rect 309915 319500 309916 319564
rect 309980 319500 309981 319564
rect 309915 319499 309981 319500
rect 310102 318613 310162 321510
rect 310835 320516 310901 320517
rect 310835 320452 310836 320516
rect 310900 320452 310901 320516
rect 310835 320451 310901 320452
rect 310283 320380 310349 320381
rect 310283 320316 310284 320380
rect 310348 320316 310349 320380
rect 310283 320315 310349 320316
rect 310651 320380 310717 320381
rect 310651 320316 310652 320380
rect 310716 320316 310717 320380
rect 310651 320315 310717 320316
rect 309363 318612 309429 318613
rect 309363 318548 309364 318612
rect 309428 318548 309429 318612
rect 309363 318547 309429 318548
rect 310099 318612 310165 318613
rect 310099 318548 310100 318612
rect 310164 318548 310165 318612
rect 310099 318547 310165 318548
rect 309366 313037 309426 318547
rect 309363 313036 309429 313037
rect 309363 312972 309364 313036
rect 309428 312972 309429 313036
rect 309363 312971 309429 312972
rect 310286 312221 310346 320315
rect 310654 319565 310714 320315
rect 310651 319564 310717 319565
rect 310651 319500 310652 319564
rect 310716 319500 310717 319564
rect 310651 319499 310717 319500
rect 310838 319293 310898 320451
rect 311022 320381 311082 369547
rect 311203 369476 311269 369477
rect 311203 369412 311204 369476
rect 311268 369412 311269 369476
rect 311203 369411 311269 369412
rect 312491 369476 312557 369477
rect 312491 369412 312492 369476
rect 312556 369412 312557 369476
rect 312491 369411 312557 369412
rect 311019 320380 311085 320381
rect 311019 320316 311020 320380
rect 311084 320316 311085 320380
rect 311019 320315 311085 320316
rect 311206 320109 311266 369411
rect 312494 325710 312554 369411
rect 312494 325650 312738 325710
rect 312678 321570 312738 325650
rect 312126 321510 312738 321570
rect 311387 320380 311453 320381
rect 311387 320316 311388 320380
rect 311452 320316 311453 320380
rect 311387 320315 311453 320316
rect 311203 320108 311269 320109
rect 311203 320044 311204 320108
rect 311268 320044 311269 320108
rect 311203 320043 311269 320044
rect 310835 319292 310901 319293
rect 310835 319228 310836 319292
rect 310900 319228 310901 319292
rect 310835 319227 310901 319228
rect 310283 312220 310349 312221
rect 310283 312156 310284 312220
rect 310348 312156 310349 312220
rect 310283 312155 310349 312156
rect 308259 309908 308325 309909
rect 308259 309844 308260 309908
rect 308324 309844 308325 309908
rect 308259 309843 308325 309844
rect 307707 228580 307773 228581
rect 307707 228516 307708 228580
rect 307772 228516 307773 228580
rect 307707 228515 307773 228516
rect 308262 222053 308322 309843
rect 310467 299300 310533 299301
rect 310467 299236 310468 299300
rect 310532 299236 310533 299300
rect 310467 299235 310533 299236
rect 310470 230213 310530 299235
rect 311206 296730 311266 320043
rect 311390 312493 311450 320315
rect 311939 320108 312005 320109
rect 311939 320044 311940 320108
rect 312004 320044 312005 320108
rect 311939 320043 312005 320044
rect 311755 317932 311821 317933
rect 311755 317868 311756 317932
rect 311820 317868 311821 317932
rect 311755 317867 311821 317868
rect 311387 312492 311453 312493
rect 311387 312428 311388 312492
rect 311452 312428 311453 312492
rect 311387 312427 311453 312428
rect 311758 299301 311818 317867
rect 311942 312629 312002 320043
rect 311939 312628 312005 312629
rect 311939 312564 311940 312628
rect 312004 312564 312005 312628
rect 311939 312563 312005 312564
rect 311755 299300 311821 299301
rect 311755 299236 311756 299300
rect 311820 299236 311821 299300
rect 311755 299235 311821 299236
rect 310654 296670 311266 296730
rect 310654 293725 310714 296670
rect 310651 293724 310717 293725
rect 310651 293660 310652 293724
rect 310716 293660 310717 293724
rect 310651 293659 310717 293660
rect 312126 291005 312186 321510
rect 312678 320653 312738 321510
rect 312675 320652 312741 320653
rect 312675 320588 312676 320652
rect 312740 320588 312741 320652
rect 312675 320587 312741 320588
rect 313046 320109 313106 395931
rect 314331 377772 314397 377773
rect 314331 377708 314332 377772
rect 314396 377708 314397 377772
rect 314331 377707 314397 377708
rect 313779 369612 313845 369613
rect 313779 369548 313780 369612
rect 313844 369548 313845 369612
rect 313779 369547 313845 369548
rect 313595 369476 313661 369477
rect 313595 369412 313596 369476
rect 313660 369412 313661 369476
rect 313595 369411 313661 369412
rect 313598 320109 313658 369411
rect 312491 320108 312557 320109
rect 312491 320044 312492 320108
rect 312556 320044 312557 320108
rect 312491 320043 312557 320044
rect 313043 320108 313109 320109
rect 313043 320044 313044 320108
rect 313108 320044 313109 320108
rect 313043 320043 313109 320044
rect 313595 320108 313661 320109
rect 313595 320044 313596 320108
rect 313660 320044 313661 320108
rect 313595 320043 313661 320044
rect 312494 296730 312554 320043
rect 313782 317933 313842 369547
rect 314334 320245 314394 377707
rect 315619 370564 315685 370565
rect 315619 370500 315620 370564
rect 315684 370500 315685 370564
rect 315619 370499 315685 370500
rect 315435 369748 315501 369749
rect 315435 369684 315436 369748
rect 315500 369684 315501 369748
rect 315435 369683 315501 369684
rect 314883 320652 314949 320653
rect 314883 320588 314884 320652
rect 314948 320588 314949 320652
rect 314883 320587 314949 320588
rect 313963 320244 314029 320245
rect 313963 320180 313964 320244
rect 314028 320180 314029 320244
rect 313963 320179 314029 320180
rect 314331 320244 314397 320245
rect 314331 320180 314332 320244
rect 314396 320180 314397 320244
rect 314331 320179 314397 320180
rect 313966 319701 314026 320179
rect 314147 320108 314213 320109
rect 314147 320044 314148 320108
rect 314212 320044 314213 320108
rect 314147 320043 314213 320044
rect 313963 319700 314029 319701
rect 313963 319636 313964 319700
rect 314028 319636 314029 319700
rect 313963 319635 314029 319636
rect 313779 317932 313845 317933
rect 313779 317868 313780 317932
rect 313844 317868 313845 317932
rect 313779 317867 313845 317868
rect 312675 317524 312741 317525
rect 312675 317460 312676 317524
rect 312740 317460 312741 317524
rect 312675 317459 312741 317460
rect 312678 308821 312738 317459
rect 312675 308820 312741 308821
rect 312675 308756 312676 308820
rect 312740 308756 312741 308820
rect 312675 308755 312741 308756
rect 312310 296670 312554 296730
rect 312123 291004 312189 291005
rect 312123 290940 312124 291004
rect 312188 290940 312189 291004
rect 312123 290939 312189 290940
rect 310467 230212 310533 230213
rect 310467 230148 310468 230212
rect 310532 230148 310533 230212
rect 310467 230147 310533 230148
rect 308259 222052 308325 222053
rect 308259 221988 308260 222052
rect 308324 221988 308325 222052
rect 308259 221987 308325 221988
rect 306971 219060 307037 219061
rect 306971 218996 306972 219060
rect 307036 218996 307037 219060
rect 306971 218995 307037 218996
rect 312310 218925 312370 296670
rect 313782 290733 313842 317867
rect 314150 315621 314210 320043
rect 314147 315620 314213 315621
rect 314147 315556 314148 315620
rect 314212 315556 314213 315620
rect 314147 315555 314213 315556
rect 313779 290732 313845 290733
rect 313779 290668 313780 290732
rect 313844 290668 313845 290732
rect 313779 290667 313845 290668
rect 314334 223141 314394 320179
rect 314331 223140 314397 223141
rect 314331 223076 314332 223140
rect 314396 223076 314397 223140
rect 314331 223075 314397 223076
rect 314886 220285 314946 320587
rect 315067 320108 315133 320109
rect 315067 320044 315068 320108
rect 315132 320044 315133 320108
rect 315067 320043 315133 320044
rect 314883 220284 314949 220285
rect 314883 220220 314884 220284
rect 314948 220220 314949 220284
rect 314883 220219 314949 220220
rect 315070 219197 315130 320043
rect 315438 319701 315498 369683
rect 315622 320109 315682 370499
rect 315806 320653 315866 396883
rect 317275 390556 317341 390557
rect 317275 390492 317276 390556
rect 317340 390492 317341 390556
rect 317275 390491 317341 390492
rect 317091 390148 317157 390149
rect 317091 390084 317092 390148
rect 317156 390084 317157 390148
rect 317091 390083 317157 390084
rect 315803 320652 315869 320653
rect 315803 320588 315804 320652
rect 315868 320588 315869 320652
rect 315803 320587 315869 320588
rect 316907 320652 316973 320653
rect 316907 320588 316908 320652
rect 316972 320588 316973 320652
rect 316907 320587 316973 320588
rect 315619 320108 315685 320109
rect 315619 320044 315620 320108
rect 315684 320044 315685 320108
rect 315619 320043 315685 320044
rect 316723 320108 316789 320109
rect 316723 320044 316724 320108
rect 316788 320044 316789 320108
rect 316723 320043 316789 320044
rect 315435 319700 315501 319701
rect 315435 319636 315436 319700
rect 315500 319636 315501 319700
rect 315435 319635 315501 319636
rect 316355 318748 316421 318749
rect 316355 318684 316356 318748
rect 316420 318684 316421 318748
rect 316355 318683 316421 318684
rect 315619 317524 315685 317525
rect 315619 317460 315620 317524
rect 315684 317460 315685 317524
rect 315619 317459 315685 317460
rect 315622 309909 315682 317459
rect 315619 309908 315685 309909
rect 315619 309844 315620 309908
rect 315684 309844 315685 309908
rect 315619 309843 315685 309844
rect 316358 264485 316418 318683
rect 316539 317524 316605 317525
rect 316539 317460 316540 317524
rect 316604 317460 316605 317524
rect 316539 317459 316605 317460
rect 316542 305829 316602 317459
rect 316726 315349 316786 320043
rect 316910 318477 316970 320587
rect 317094 318749 317154 390083
rect 317278 320109 317338 390491
rect 318011 369476 318077 369477
rect 318011 369412 318012 369476
rect 318076 369412 318077 369476
rect 318011 369411 318077 369412
rect 318014 328470 318074 369411
rect 317646 328410 318074 328470
rect 317459 320652 317525 320653
rect 317459 320588 317460 320652
rect 317524 320588 317525 320652
rect 317459 320587 317525 320588
rect 317275 320108 317341 320109
rect 317275 320044 317276 320108
rect 317340 320044 317341 320108
rect 317275 320043 317341 320044
rect 317462 319565 317522 320587
rect 317646 320109 317706 328410
rect 318011 320652 318077 320653
rect 318011 320588 318012 320652
rect 318076 320588 318077 320652
rect 318011 320587 318077 320588
rect 318195 320652 318261 320653
rect 318195 320588 318196 320652
rect 318260 320588 318261 320652
rect 318195 320587 318261 320588
rect 317643 320108 317709 320109
rect 317643 320044 317644 320108
rect 317708 320044 317709 320108
rect 317643 320043 317709 320044
rect 317459 319564 317525 319565
rect 317459 319500 317460 319564
rect 317524 319500 317525 319564
rect 317459 319499 317525 319500
rect 317091 318748 317157 318749
rect 317091 318684 317092 318748
rect 317156 318684 317157 318748
rect 317091 318683 317157 318684
rect 316907 318476 316973 318477
rect 316907 318412 316908 318476
rect 316972 318412 316973 318476
rect 316907 318411 316973 318412
rect 317275 317660 317341 317661
rect 317275 317596 317276 317660
rect 317340 317596 317341 317660
rect 317275 317595 317341 317596
rect 316723 315348 316789 315349
rect 316723 315284 316724 315348
rect 316788 315284 316789 315348
rect 316723 315283 316789 315284
rect 316539 305828 316605 305829
rect 316539 305764 316540 305828
rect 316604 305764 316605 305828
rect 316539 305763 316605 305764
rect 317278 299301 317338 317595
rect 317275 299300 317341 299301
rect 317275 299236 317276 299300
rect 317340 299236 317341 299300
rect 317275 299235 317341 299236
rect 317646 268429 317706 320043
rect 318014 319021 318074 320587
rect 318198 319429 318258 320587
rect 318566 320245 318626 397019
rect 320035 390420 320101 390421
rect 320035 390356 320036 390420
rect 320100 390356 320101 390420
rect 320035 390355 320101 390356
rect 319299 369612 319365 369613
rect 319299 369548 319300 369612
rect 319364 369548 319365 369612
rect 319299 369547 319365 369548
rect 319302 325710 319362 369547
rect 319667 369476 319733 369477
rect 319667 369412 319668 369476
rect 319732 369412 319733 369476
rect 319667 369411 319733 369412
rect 319118 325650 319362 325710
rect 318931 321196 318997 321197
rect 318931 321132 318932 321196
rect 318996 321132 318997 321196
rect 318931 321131 318997 321132
rect 318934 320653 318994 321131
rect 318931 320652 318997 320653
rect 318931 320588 318932 320652
rect 318996 320588 318997 320652
rect 318931 320587 318997 320588
rect 318563 320244 318629 320245
rect 318563 320180 318564 320244
rect 318628 320180 318629 320244
rect 318563 320179 318629 320180
rect 318195 319428 318261 319429
rect 318195 319364 318196 319428
rect 318260 319364 318261 319428
rect 318195 319363 318261 319364
rect 318011 319020 318077 319021
rect 318011 318956 318012 319020
rect 318076 318956 318077 319020
rect 318011 318955 318077 318956
rect 318379 317524 318445 317525
rect 318379 317460 318380 317524
rect 318444 317460 318445 317524
rect 318379 317459 318445 317460
rect 318382 311677 318442 317459
rect 318379 311676 318445 311677
rect 318379 311612 318380 311676
rect 318444 311612 318445 311676
rect 318379 311611 318445 311612
rect 318566 296730 318626 320179
rect 319118 320109 319178 325650
rect 319299 320380 319365 320381
rect 319299 320316 319300 320380
rect 319364 320316 319365 320380
rect 319299 320315 319365 320316
rect 319115 320108 319181 320109
rect 319115 320044 319116 320108
rect 319180 320044 319181 320108
rect 319115 320043 319181 320044
rect 318747 318068 318813 318069
rect 318747 318004 318748 318068
rect 318812 318004 318813 318068
rect 318747 318003 318813 318004
rect 318750 314533 318810 318003
rect 319118 316709 319178 320043
rect 319302 319429 319362 320315
rect 319483 320108 319549 320109
rect 319483 320044 319484 320108
rect 319548 320044 319549 320108
rect 319483 320043 319549 320044
rect 319299 319428 319365 319429
rect 319299 319364 319300 319428
rect 319364 319364 319365 319428
rect 319299 319363 319365 319364
rect 319115 316708 319181 316709
rect 319115 316644 319116 316708
rect 319180 316644 319181 316708
rect 319115 316643 319181 316644
rect 318747 314532 318813 314533
rect 318747 314468 318748 314532
rect 318812 314468 318813 314532
rect 318747 314467 318813 314468
rect 319486 311910 319546 320043
rect 319670 318749 319730 369411
rect 320038 320109 320098 390355
rect 324267 372332 324333 372333
rect 324267 372268 324268 372332
rect 324332 372268 324333 372332
rect 324267 372267 324333 372268
rect 323163 371516 323229 371517
rect 323163 371452 323164 371516
rect 323228 371452 323229 371516
rect 323163 371451 323229 371452
rect 320955 369612 321021 369613
rect 320955 369548 320956 369612
rect 321020 369548 321021 369612
rect 320955 369547 321021 369548
rect 320771 322012 320837 322013
rect 320771 321948 320772 322012
rect 320836 321948 320837 322012
rect 320771 321947 320837 321948
rect 320587 321468 320653 321469
rect 320587 321404 320588 321468
rect 320652 321404 320653 321468
rect 320587 321403 320653 321404
rect 320590 320381 320650 321403
rect 320587 320380 320653 320381
rect 320587 320316 320588 320380
rect 320652 320316 320653 320380
rect 320587 320315 320653 320316
rect 320035 320108 320101 320109
rect 320035 320044 320036 320108
rect 320100 320044 320101 320108
rect 320035 320043 320101 320044
rect 320403 320108 320469 320109
rect 320403 320044 320404 320108
rect 320468 320044 320469 320108
rect 320403 320043 320469 320044
rect 320406 319429 320466 320043
rect 320403 319428 320469 319429
rect 320403 319364 320404 319428
rect 320468 319364 320469 319428
rect 320403 319363 320469 319364
rect 319667 318748 319733 318749
rect 319667 318684 319668 318748
rect 319732 318684 319733 318748
rect 319667 318683 319733 318684
rect 320774 317933 320834 321947
rect 320958 321333 321018 369547
rect 321139 369476 321205 369477
rect 321139 369412 321140 369476
rect 321204 369412 321205 369476
rect 321139 369411 321205 369412
rect 320955 321332 321021 321333
rect 320955 321268 320956 321332
rect 321020 321268 321021 321332
rect 320955 321267 321021 321268
rect 320771 317932 320837 317933
rect 320771 317868 320772 317932
rect 320836 317868 320837 317932
rect 320771 317867 320837 317868
rect 320219 317796 320285 317797
rect 320219 317732 320220 317796
rect 320284 317732 320285 317796
rect 320219 317731 320285 317732
rect 318934 311850 319546 311910
rect 318747 311676 318813 311677
rect 318747 311612 318748 311676
rect 318812 311612 318813 311676
rect 318747 311611 318813 311612
rect 318750 310861 318810 311611
rect 318747 310860 318813 310861
rect 318747 310796 318748 310860
rect 318812 310796 318813 310860
rect 318747 310795 318813 310796
rect 317830 296670 318626 296730
rect 317643 268428 317709 268429
rect 317643 268364 317644 268428
rect 317708 268364 317709 268428
rect 317643 268363 317709 268364
rect 316355 264484 316421 264485
rect 316355 264420 316356 264484
rect 316420 264420 316421 264484
rect 316355 264419 316421 264420
rect 317830 246533 317890 296670
rect 318934 272509 318994 311850
rect 318931 272508 318997 272509
rect 318931 272444 318932 272508
rect 318996 272444 318997 272508
rect 318931 272443 318997 272444
rect 317827 246532 317893 246533
rect 317827 246468 317828 246532
rect 317892 246468 317893 246532
rect 317827 246467 317893 246468
rect 320222 224773 320282 317731
rect 320958 311910 321018 321267
rect 321142 319021 321202 369411
rect 323166 364989 323226 371451
rect 324270 366349 324330 372267
rect 324267 366348 324333 366349
rect 324267 366284 324268 366348
rect 324332 366284 324333 366348
rect 324267 366283 324333 366284
rect 323163 364988 323229 364989
rect 323163 364924 323164 364988
rect 323228 364924 323229 364988
rect 323163 364923 323229 364924
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 323715 356692 323781 356693
rect 323715 356628 323716 356692
rect 323780 356628 323781 356692
rect 323715 356627 323781 356628
rect 323531 324460 323597 324461
rect 323531 324396 323532 324460
rect 323596 324396 323597 324460
rect 323531 324395 323597 324396
rect 321507 321332 321573 321333
rect 321507 321268 321508 321332
rect 321572 321268 321573 321332
rect 321507 321267 321573 321268
rect 322979 321332 323045 321333
rect 322979 321268 322980 321332
rect 323044 321268 323045 321332
rect 322979 321267 323045 321268
rect 321323 321060 321389 321061
rect 321323 320996 321324 321060
rect 321388 320996 321389 321060
rect 321323 320995 321389 320996
rect 321326 320653 321386 320995
rect 321323 320652 321389 320653
rect 321323 320588 321324 320652
rect 321388 320588 321389 320652
rect 321323 320587 321389 320588
rect 321323 320380 321389 320381
rect 321323 320316 321324 320380
rect 321388 320316 321389 320380
rect 321323 320315 321389 320316
rect 321326 319429 321386 320315
rect 321510 320109 321570 321267
rect 322982 320653 323042 321267
rect 323534 320789 323594 324395
rect 323531 320788 323597 320789
rect 323531 320724 323532 320788
rect 323596 320724 323597 320788
rect 323531 320723 323597 320724
rect 322979 320652 323045 320653
rect 322979 320588 322980 320652
rect 323044 320588 323045 320652
rect 323718 320650 323778 356627
rect 323899 342956 323965 342957
rect 323899 342892 323900 342956
rect 323964 342892 323965 342956
rect 323899 342891 323965 342892
rect 322979 320587 323045 320588
rect 323534 320590 323778 320650
rect 323534 320517 323594 320590
rect 322059 320516 322125 320517
rect 322059 320452 322060 320516
rect 322124 320452 322125 320516
rect 322059 320451 322125 320452
rect 322611 320516 322677 320517
rect 322611 320452 322612 320516
rect 322676 320452 322677 320516
rect 322611 320451 322677 320452
rect 323347 320516 323413 320517
rect 323347 320452 323348 320516
rect 323412 320452 323413 320516
rect 323347 320451 323413 320452
rect 323531 320516 323597 320517
rect 323531 320452 323532 320516
rect 323596 320452 323597 320516
rect 323531 320451 323597 320452
rect 321507 320108 321573 320109
rect 321507 320044 321508 320108
rect 321572 320044 321573 320108
rect 321507 320043 321573 320044
rect 322062 319565 322122 320451
rect 322427 320380 322493 320381
rect 322427 320316 322428 320380
rect 322492 320316 322493 320380
rect 322427 320315 322493 320316
rect 322430 319701 322490 320315
rect 322427 319700 322493 319701
rect 322427 319636 322428 319700
rect 322492 319636 322493 319700
rect 322427 319635 322493 319636
rect 322059 319564 322125 319565
rect 322059 319500 322060 319564
rect 322124 319500 322125 319564
rect 322059 319499 322125 319500
rect 321323 319428 321389 319429
rect 321323 319364 321324 319428
rect 321388 319364 321389 319428
rect 321323 319363 321389 319364
rect 322614 319021 322674 320451
rect 323350 319021 323410 320451
rect 321139 319020 321205 319021
rect 321139 318956 321140 319020
rect 321204 318956 321205 319020
rect 321139 318955 321205 318956
rect 322611 319020 322677 319021
rect 322611 318956 322612 319020
rect 322676 318956 322677 319020
rect 322611 318955 322677 318956
rect 323347 319020 323413 319021
rect 323347 318956 323348 319020
rect 323412 318956 323413 319020
rect 323347 318955 323413 318956
rect 323347 318476 323413 318477
rect 323347 318412 323348 318476
rect 323412 318412 323413 318476
rect 323347 318411 323413 318412
rect 323163 317932 323229 317933
rect 323163 317868 323164 317932
rect 323228 317868 323229 317932
rect 323163 317867 323229 317868
rect 321323 317524 321389 317525
rect 321323 317460 321324 317524
rect 321388 317460 321389 317524
rect 321323 317459 321389 317460
rect 321691 317524 321757 317525
rect 321691 317460 321692 317524
rect 321756 317460 321757 317524
rect 321691 317459 321757 317460
rect 320406 311850 321018 311910
rect 320406 261493 320466 311850
rect 321326 306390 321386 317459
rect 321694 311910 321754 317459
rect 320774 306330 321386 306390
rect 321510 311850 321754 311910
rect 320774 304877 320834 306330
rect 320771 304876 320837 304877
rect 320771 304812 320772 304876
rect 320836 304812 320837 304876
rect 320771 304811 320837 304812
rect 320403 261492 320469 261493
rect 320403 261428 320404 261492
rect 320468 261428 320469 261492
rect 320403 261427 320469 261428
rect 320219 224772 320285 224773
rect 320219 224708 320220 224772
rect 320284 224708 320285 224772
rect 320219 224707 320285 224708
rect 320774 223413 320834 304811
rect 321510 301477 321570 311850
rect 321507 301476 321573 301477
rect 321507 301412 321508 301476
rect 321572 301412 321573 301476
rect 321507 301411 321573 301412
rect 323166 245173 323226 317867
rect 323350 258909 323410 318411
rect 323347 258908 323413 258909
rect 323347 258844 323348 258908
rect 323412 258844 323413 258908
rect 323347 258843 323413 258844
rect 323163 245172 323229 245173
rect 323163 245108 323164 245172
rect 323228 245108 323229 245172
rect 323163 245107 323229 245108
rect 323534 226269 323594 320451
rect 323902 320381 323962 342891
rect 325371 341460 325437 341461
rect 325371 341396 325372 341460
rect 325436 341396 325437 341460
rect 325371 341395 325437 341396
rect 324635 340100 324701 340101
rect 324635 340036 324636 340100
rect 324700 340036 324701 340100
rect 324635 340035 324701 340036
rect 324083 323644 324149 323645
rect 324083 323580 324084 323644
rect 324148 323580 324149 323644
rect 324083 323579 324149 323580
rect 324086 320789 324146 323579
rect 324451 322148 324517 322149
rect 324451 322084 324452 322148
rect 324516 322084 324517 322148
rect 324451 322083 324517 322084
rect 324083 320788 324149 320789
rect 324083 320724 324084 320788
rect 324148 320724 324149 320788
rect 324083 320723 324149 320724
rect 323899 320380 323965 320381
rect 323899 320316 323900 320380
rect 323964 320316 323965 320380
rect 323899 320315 323965 320316
rect 323902 319701 323962 320315
rect 324086 319701 324146 320723
rect 324454 320381 324514 322083
rect 324267 320380 324333 320381
rect 324267 320316 324268 320380
rect 324332 320316 324333 320380
rect 324267 320315 324333 320316
rect 324451 320380 324517 320381
rect 324451 320316 324452 320380
rect 324516 320316 324517 320380
rect 324451 320315 324517 320316
rect 323899 319700 323965 319701
rect 323899 319636 323900 319700
rect 323964 319636 323965 319700
rect 323899 319635 323965 319636
rect 324083 319700 324149 319701
rect 324083 319636 324084 319700
rect 324148 319636 324149 319700
rect 324083 319635 324149 319636
rect 324270 319021 324330 320315
rect 324267 319020 324333 319021
rect 324267 318956 324268 319020
rect 324332 318956 324333 319020
rect 324267 318955 324333 318956
rect 324454 255917 324514 320315
rect 324638 320109 324698 340035
rect 325374 327181 325434 341395
rect 325794 327454 326414 362898
rect 329514 705798 330134 705830
rect 329514 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 330134 705798
rect 329514 705478 330134 705562
rect 329514 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 330134 705478
rect 329514 691174 330134 705242
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 439174 330134 474618
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 343587 452164 343653 452165
rect 343587 452100 343588 452164
rect 343652 452100 343653 452164
rect 343587 452099 343653 452100
rect 343590 446453 343650 452099
rect 357387 451620 357453 451621
rect 357387 451556 357388 451620
rect 357452 451556 357453 451620
rect 357387 451555 357453 451556
rect 346347 451484 346413 451485
rect 346347 451420 346348 451484
rect 346412 451420 346413 451484
rect 346347 451419 346413 451420
rect 343955 449444 344021 449445
rect 343955 449380 343956 449444
rect 344020 449380 344021 449444
rect 343955 449379 344021 449380
rect 345243 449444 345309 449445
rect 345243 449380 345244 449444
rect 345308 449380 345309 449444
rect 345243 449379 345309 449380
rect 343587 446452 343653 446453
rect 343587 446388 343588 446452
rect 343652 446388 343653 446452
rect 343587 446387 343653 446388
rect 343958 444957 344018 449379
rect 344875 449308 344941 449309
rect 344875 449244 344876 449308
rect 344940 449244 344941 449308
rect 344875 449243 344941 449244
rect 343955 444956 344021 444957
rect 343955 444892 343956 444956
rect 344020 444892 344021 444956
rect 343955 444891 344021 444892
rect 329514 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 330134 439174
rect 329514 438854 330134 438938
rect 329514 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 330134 438854
rect 329514 403174 330134 438618
rect 329514 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 330134 403174
rect 329514 402854 330134 402938
rect 329514 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 330134 402854
rect 329514 367174 330134 402618
rect 343219 400620 343285 400621
rect 343219 400556 343220 400620
rect 343284 400556 343285 400620
rect 343219 400555 343285 400556
rect 343222 399261 343282 400555
rect 344878 400077 344938 449243
rect 345246 401981 345306 449379
rect 346350 447813 346410 451419
rect 347635 451348 347701 451349
rect 347635 451284 347636 451348
rect 347700 451284 347701 451348
rect 347635 451283 347701 451284
rect 355179 451348 355245 451349
rect 355179 451284 355180 451348
rect 355244 451284 355245 451348
rect 355179 451283 355245 451284
rect 346347 447812 346413 447813
rect 346347 447748 346348 447812
rect 346412 447748 346413 447812
rect 346347 447747 346413 447748
rect 345243 401980 345309 401981
rect 345243 401916 345244 401980
rect 345308 401916 345309 401980
rect 345243 401915 345309 401916
rect 347638 400893 347698 451283
rect 349659 449444 349725 449445
rect 349659 449380 349660 449444
rect 349724 449380 349725 449444
rect 349659 449379 349725 449380
rect 353339 449444 353405 449445
rect 353339 449380 353340 449444
rect 353404 449380 353405 449444
rect 353339 449379 353405 449380
rect 347635 400892 347701 400893
rect 346534 400830 347330 400890
rect 344875 400076 344941 400077
rect 344875 400012 344876 400076
rect 344940 400012 344941 400076
rect 344875 400011 344941 400012
rect 346534 399941 346594 400830
rect 346531 399940 346597 399941
rect 346531 399876 346532 399940
rect 346596 399876 346597 399940
rect 346531 399875 346597 399876
rect 346899 399940 346965 399941
rect 346899 399876 346900 399940
rect 346964 399876 346965 399940
rect 346899 399875 346965 399876
rect 347083 399940 347149 399941
rect 347083 399876 347084 399940
rect 347148 399876 347149 399940
rect 347083 399875 347149 399876
rect 346347 399804 346413 399805
rect 346347 399740 346348 399804
rect 346412 399802 346413 399804
rect 346715 399804 346781 399805
rect 346412 399742 346594 399802
rect 346412 399740 346413 399742
rect 346347 399739 346413 399740
rect 346347 399532 346413 399533
rect 346347 399468 346348 399532
rect 346412 399468 346413 399532
rect 346347 399467 346413 399468
rect 343219 399260 343285 399261
rect 343219 399196 343220 399260
rect 343284 399196 343285 399260
rect 343219 399195 343285 399196
rect 346350 398853 346410 399467
rect 346347 398852 346413 398853
rect 346347 398788 346348 398852
rect 346412 398788 346413 398852
rect 346347 398787 346413 398788
rect 346534 398581 346594 399742
rect 346715 399740 346716 399804
rect 346780 399740 346781 399804
rect 346715 399739 346781 399740
rect 346531 398580 346597 398581
rect 346531 398516 346532 398580
rect 346596 398516 346597 398580
rect 346531 398515 346597 398516
rect 345243 398036 345309 398037
rect 345243 397972 345244 398036
rect 345308 397972 345309 398036
rect 345243 397971 345309 397972
rect 345059 396132 345125 396133
rect 345059 396068 345060 396132
rect 345124 396068 345125 396132
rect 345059 396067 345125 396068
rect 343587 395860 343653 395861
rect 343587 395796 343588 395860
rect 343652 395796 343653 395860
rect 343587 395795 343653 395796
rect 343035 386884 343101 386885
rect 343035 386820 343036 386884
rect 343100 386820 343101 386884
rect 343035 386819 343101 386820
rect 342851 386748 342917 386749
rect 342851 386684 342852 386748
rect 342916 386684 342917 386748
rect 342851 386683 342917 386684
rect 330523 385932 330589 385933
rect 330523 385868 330524 385932
rect 330588 385868 330589 385932
rect 330523 385867 330589 385868
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 331174 330134 366618
rect 329514 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 330134 331174
rect 329514 330854 330134 330938
rect 329514 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 330134 330854
rect 329235 330580 329301 330581
rect 329235 330516 329236 330580
rect 329300 330516 329301 330580
rect 329235 330515 329301 330516
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325371 327180 325437 327181
rect 325371 327116 325372 327180
rect 325436 327116 325437 327180
rect 325371 327115 325437 327116
rect 325794 327134 326414 327218
rect 325374 320789 325434 327115
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 324819 320788 324885 320789
rect 324819 320724 324820 320788
rect 324884 320724 324885 320788
rect 324819 320723 324885 320724
rect 325371 320788 325437 320789
rect 325371 320724 325372 320788
rect 325436 320724 325437 320788
rect 325371 320723 325437 320724
rect 324635 320108 324701 320109
rect 324635 320044 324636 320108
rect 324700 320044 324701 320108
rect 324635 320043 324701 320044
rect 324451 255916 324517 255917
rect 324451 255852 324452 255916
rect 324516 255852 324517 255916
rect 324451 255851 324517 255852
rect 324638 250613 324698 320043
rect 324822 319701 324882 320723
rect 325003 320516 325069 320517
rect 325003 320452 325004 320516
rect 325068 320452 325069 320516
rect 325003 320451 325069 320452
rect 324819 319700 324885 319701
rect 324819 319636 324820 319700
rect 324884 319636 324885 319700
rect 324819 319635 324885 319636
rect 325006 319021 325066 320451
rect 325003 319020 325069 319021
rect 325003 318956 325004 319020
rect 325068 318956 325069 319020
rect 325003 318955 325069 318956
rect 325794 291454 326414 326898
rect 329238 325710 329298 330515
rect 328502 325650 329298 325710
rect 327763 322964 327829 322965
rect 327763 322900 327764 322964
rect 327828 322900 327829 322964
rect 327763 322899 327829 322900
rect 326659 322284 326725 322285
rect 326659 322220 326660 322284
rect 326724 322220 326725 322284
rect 326659 322219 326725 322220
rect 326662 320789 326722 322219
rect 327395 321604 327461 321605
rect 327395 321540 327396 321604
rect 327460 321540 327461 321604
rect 327395 321539 327461 321540
rect 326659 320788 326725 320789
rect 326659 320724 326660 320788
rect 326724 320724 326725 320788
rect 326659 320723 326725 320724
rect 327398 320381 327458 321539
rect 327766 320381 327826 322899
rect 326659 320380 326725 320381
rect 326659 320316 326660 320380
rect 326724 320316 326725 320380
rect 326659 320315 326725 320316
rect 327395 320380 327461 320381
rect 327395 320316 327396 320380
rect 327460 320316 327461 320380
rect 327395 320315 327461 320316
rect 327763 320380 327829 320381
rect 327763 320316 327764 320380
rect 327828 320316 327829 320380
rect 327763 320315 327829 320316
rect 326662 319021 326722 320315
rect 326843 320108 326909 320109
rect 326843 320044 326844 320108
rect 326908 320044 326909 320108
rect 326843 320043 326909 320044
rect 326846 319565 326906 320043
rect 326843 319564 326909 319565
rect 326843 319500 326844 319564
rect 326908 319500 326909 319564
rect 326843 319499 326909 319500
rect 327398 319021 327458 320315
rect 326659 319020 326725 319021
rect 326659 318956 326660 319020
rect 326724 318956 326725 319020
rect 326659 318955 326725 318956
rect 327395 319020 327461 319021
rect 327395 318956 327396 319020
rect 327460 318956 327461 319020
rect 327395 318955 327461 318956
rect 328502 318613 328562 325650
rect 328499 318612 328565 318613
rect 328499 318548 328500 318612
rect 328564 318548 328565 318612
rect 328499 318547 328565 318548
rect 326659 317796 326725 317797
rect 326659 317732 326660 317796
rect 326724 317732 326725 317796
rect 326659 317731 326725 317732
rect 328315 317796 328381 317797
rect 328315 317732 328316 317796
rect 328380 317732 328381 317796
rect 328315 317731 328381 317732
rect 326662 316437 326722 317731
rect 327027 317660 327093 317661
rect 327027 317596 327028 317660
rect 327092 317596 327093 317660
rect 327027 317595 327093 317596
rect 326659 316436 326725 316437
rect 326659 316372 326660 316436
rect 326724 316372 326725 316436
rect 326659 316371 326725 316372
rect 327030 312629 327090 317595
rect 327027 312628 327093 312629
rect 327027 312564 327028 312628
rect 327092 312564 327093 312628
rect 327027 312563 327093 312564
rect 328318 306390 328378 317731
rect 327582 306330 328378 306390
rect 327582 305013 327642 306330
rect 327579 305012 327645 305013
rect 327579 304948 327580 305012
rect 327644 304948 327645 305012
rect 327579 304947 327645 304948
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 324635 250612 324701 250613
rect 324635 250548 324636 250612
rect 324700 250548 324701 250612
rect 324635 250547 324701 250548
rect 323531 226268 323597 226269
rect 323531 226204 323532 226268
rect 323596 226204 323597 226268
rect 323531 226203 323597 226204
rect 320771 223412 320837 223413
rect 320771 223348 320772 223412
rect 320836 223348 320837 223412
rect 320771 223347 320837 223348
rect 325794 219454 326414 254898
rect 327582 228717 327642 304947
rect 327579 228716 327645 228717
rect 327579 228652 327580 228716
rect 327644 228652 327645 228716
rect 327579 228651 327645 228652
rect 328502 227357 328562 318547
rect 329051 317932 329117 317933
rect 329051 317868 329052 317932
rect 329116 317868 329117 317932
rect 329051 317867 329117 317868
rect 328867 316300 328933 316301
rect 328867 316236 328868 316300
rect 328932 316236 328933 316300
rect 328867 316235 328933 316236
rect 328683 316164 328749 316165
rect 328683 316100 328684 316164
rect 328748 316100 328749 316164
rect 328683 316099 328749 316100
rect 328686 235925 328746 316099
rect 328683 235924 328749 235925
rect 328683 235860 328684 235924
rect 328748 235860 328749 235924
rect 328683 235859 328749 235860
rect 328870 235517 328930 316235
rect 329054 306917 329114 317867
rect 329051 306916 329117 306917
rect 329051 306852 329052 306916
rect 329116 306852 329117 306916
rect 329051 306851 329117 306852
rect 329514 295174 330134 330618
rect 330339 322284 330405 322285
rect 330339 322220 330340 322284
rect 330404 322220 330405 322284
rect 330339 322219 330405 322220
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 328867 235516 328933 235517
rect 328867 235452 328868 235516
rect 328932 235452 328933 235516
rect 328867 235451 328933 235452
rect 328499 227356 328565 227357
rect 328499 227292 328500 227356
rect 328564 227292 328565 227356
rect 328499 227291 328565 227292
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 315067 219196 315133 219197
rect 315067 219132 315068 219196
rect 315132 219132 315133 219196
rect 315067 219131 315133 219132
rect 325794 219134 326414 219218
rect 312307 218924 312373 218925
rect 312307 218860 312308 218924
rect 312372 218860 312373 218924
rect 312307 218859 312373 218860
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 293514 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 294134 187174
rect 293514 186854 294134 186938
rect 293514 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 294134 186854
rect 293514 151174 294134 186618
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 115174 294134 150618
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 293514 79174 294134 114618
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -1306 294134 6618
rect 293514 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 294134 -1306
rect 293514 -1626 294134 -1542
rect 293514 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 294134 -1626
rect 293514 -1894 294134 -1862
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 223174 330134 258618
rect 330342 232661 330402 322219
rect 330526 319701 330586 385867
rect 333099 370156 333165 370157
rect 333099 370092 333100 370156
rect 333164 370092 333165 370156
rect 333099 370091 333165 370092
rect 331811 370020 331877 370021
rect 331811 369956 331812 370020
rect 331876 369956 331877 370020
rect 331811 369955 331877 369956
rect 330523 319700 330589 319701
rect 330523 319636 330524 319700
rect 330588 319636 330589 319700
rect 330523 319635 330589 319636
rect 330339 232660 330405 232661
rect 330339 232596 330340 232660
rect 330404 232596 330405 232660
rect 330339 232595 330405 232596
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 331814 31789 331874 369955
rect 333102 59397 333162 370091
rect 338619 326364 338685 326365
rect 338619 326300 338620 326364
rect 338684 326300 338685 326364
rect 338619 326299 338685 326300
rect 338622 316573 338682 326299
rect 338619 316572 338685 316573
rect 338619 316508 338620 316572
rect 338684 316508 338685 316572
rect 338619 316507 338685 316508
rect 342854 308549 342914 386683
rect 343038 370701 343098 386819
rect 343590 377637 343650 395795
rect 344139 389060 344205 389061
rect 344139 388996 344140 389060
rect 344204 388996 344205 389060
rect 344139 388995 344205 388996
rect 343587 377636 343653 377637
rect 343587 377572 343588 377636
rect 343652 377572 343653 377636
rect 343587 377571 343653 377572
rect 344142 371925 344202 388995
rect 344139 371924 344205 371925
rect 344139 371860 344140 371924
rect 344204 371860 344205 371924
rect 344139 371859 344205 371860
rect 343035 370700 343101 370701
rect 343035 370636 343036 370700
rect 343100 370636 343101 370700
rect 343035 370635 343101 370636
rect 342851 308548 342917 308549
rect 342851 308484 342852 308548
rect 342916 308484 342917 308548
rect 342851 308483 342917 308484
rect 345062 295085 345122 396067
rect 345246 388517 345306 397971
rect 346718 395045 346778 399739
rect 346715 395044 346781 395045
rect 346715 394980 346716 395044
rect 346780 394980 346781 395044
rect 346715 394979 346781 394980
rect 346902 390570 346962 399875
rect 347086 395453 347146 399875
rect 347270 399805 347330 400830
rect 347635 400828 347636 400892
rect 347700 400828 347701 400892
rect 347635 400827 347701 400828
rect 348555 400620 348621 400621
rect 348555 400556 348556 400620
rect 348620 400556 348621 400620
rect 348555 400555 348621 400556
rect 348558 400077 348618 400555
rect 348555 400076 348621 400077
rect 348555 400012 348556 400076
rect 348620 400012 348621 400076
rect 348555 400011 348621 400012
rect 347819 399940 347885 399941
rect 347819 399876 347820 399940
rect 347884 399876 347885 399940
rect 347819 399875 347885 399876
rect 348187 399940 348253 399941
rect 348187 399876 348188 399940
rect 348252 399876 348253 399940
rect 348187 399875 348253 399876
rect 348739 399940 348805 399941
rect 348739 399876 348740 399940
rect 348804 399876 348805 399940
rect 348739 399875 348805 399876
rect 347267 399804 347333 399805
rect 347267 399740 347268 399804
rect 347332 399740 347333 399804
rect 347267 399739 347333 399740
rect 347822 395453 347882 399875
rect 348003 397628 348069 397629
rect 348003 397564 348004 397628
rect 348068 397564 348069 397628
rect 348003 397563 348069 397564
rect 347083 395452 347149 395453
rect 347083 395388 347084 395452
rect 347148 395388 347149 395452
rect 347083 395387 347149 395388
rect 347819 395452 347885 395453
rect 347819 395388 347820 395452
rect 347884 395388 347885 395452
rect 347819 395387 347885 395388
rect 346718 390510 346962 390570
rect 346718 389877 346778 390510
rect 346715 389876 346781 389877
rect 346715 389812 346716 389876
rect 346780 389812 346781 389876
rect 346715 389811 346781 389812
rect 345243 388516 345309 388517
rect 345243 388452 345244 388516
rect 345308 388452 345309 388516
rect 345243 388451 345309 388452
rect 348006 388381 348066 397563
rect 348190 389197 348250 399875
rect 348742 394909 348802 399875
rect 348923 399396 348989 399397
rect 348923 399332 348924 399396
rect 348988 399332 348989 399396
rect 348923 399331 348989 399332
rect 348926 398853 348986 399331
rect 348923 398852 348989 398853
rect 348923 398788 348924 398852
rect 348988 398788 348989 398852
rect 348923 398787 348989 398788
rect 349291 398444 349357 398445
rect 349291 398380 349292 398444
rect 349356 398380 349357 398444
rect 349291 398379 349357 398380
rect 349107 395044 349173 395045
rect 349107 394980 349108 395044
rect 349172 394980 349173 395044
rect 349107 394979 349173 394980
rect 348739 394908 348805 394909
rect 348739 394844 348740 394908
rect 348804 394844 348805 394908
rect 348739 394843 348805 394844
rect 348187 389196 348253 389197
rect 348187 389132 348188 389196
rect 348252 389132 348253 389196
rect 348187 389131 348253 389132
rect 348003 388380 348069 388381
rect 348003 388316 348004 388380
rect 348068 388316 348069 388380
rect 348003 388315 348069 388316
rect 349110 295221 349170 394979
rect 349294 391373 349354 398379
rect 349291 391372 349357 391373
rect 349291 391308 349292 391372
rect 349356 391308 349357 391372
rect 349291 391307 349357 391308
rect 349662 386885 349722 449379
rect 352787 401844 352853 401845
rect 352787 401780 352788 401844
rect 352852 401780 352853 401844
rect 352787 401779 352853 401780
rect 351315 400076 351381 400077
rect 351315 400012 351316 400076
rect 351380 400012 351381 400076
rect 351315 400011 351381 400012
rect 349843 399940 349909 399941
rect 349843 399876 349844 399940
rect 349908 399876 349909 399940
rect 349843 399875 349909 399876
rect 350211 399940 350277 399941
rect 350211 399876 350212 399940
rect 350276 399876 350277 399940
rect 350211 399875 350277 399876
rect 351131 399940 351197 399941
rect 351131 399876 351132 399940
rect 351196 399876 351197 399940
rect 351131 399875 351197 399876
rect 349846 395453 349906 399875
rect 350214 396813 350274 399875
rect 350763 398036 350829 398037
rect 350763 397972 350764 398036
rect 350828 397972 350829 398036
rect 350763 397971 350829 397972
rect 350579 397900 350645 397901
rect 350579 397836 350580 397900
rect 350644 397836 350645 397900
rect 350579 397835 350645 397836
rect 350211 396812 350277 396813
rect 350211 396748 350212 396812
rect 350276 396748 350277 396812
rect 350211 396747 350277 396748
rect 349843 395452 349909 395453
rect 349843 395388 349844 395452
rect 349908 395388 349909 395452
rect 349843 395387 349909 395388
rect 349659 386884 349725 386885
rect 349659 386820 349660 386884
rect 349724 386820 349725 386884
rect 349659 386819 349725 386820
rect 350582 301885 350642 397835
rect 350766 304197 350826 397971
rect 350947 396812 351013 396813
rect 350947 396748 350948 396812
rect 351012 396748 351013 396812
rect 350947 396747 351013 396748
rect 350950 358053 351010 396747
rect 351134 393549 351194 399875
rect 351318 398581 351378 400011
rect 352419 399940 352485 399941
rect 352419 399876 352420 399940
rect 352484 399876 352485 399940
rect 352419 399875 352485 399876
rect 351315 398580 351381 398581
rect 351315 398516 351316 398580
rect 351380 398516 351381 398580
rect 351315 398515 351381 398516
rect 352051 398444 352117 398445
rect 352051 398380 352052 398444
rect 352116 398380 352117 398444
rect 352051 398379 352117 398380
rect 351867 397492 351933 397493
rect 351867 397428 351868 397492
rect 351932 397428 351933 397492
rect 351867 397427 351933 397428
rect 351131 393548 351197 393549
rect 351131 393484 351132 393548
rect 351196 393484 351197 393548
rect 351131 393483 351197 393484
rect 351870 383077 351930 397427
rect 352054 394093 352114 398379
rect 352051 394092 352117 394093
rect 352051 394028 352052 394092
rect 352116 394028 352117 394092
rect 352051 394027 352117 394028
rect 351867 383076 351933 383077
rect 351867 383012 351868 383076
rect 351932 383012 351933 383076
rect 351867 383011 351933 383012
rect 350947 358052 351013 358053
rect 350947 357988 350948 358052
rect 351012 357988 351013 358052
rect 350947 357987 351013 357988
rect 352422 319837 352482 399875
rect 352790 399533 352850 401779
rect 353342 399533 353402 449379
rect 353523 400756 353589 400757
rect 353523 400692 353524 400756
rect 353588 400692 353589 400756
rect 353523 400691 353589 400692
rect 353526 399941 353586 400691
rect 354259 400620 354325 400621
rect 354259 400556 354260 400620
rect 354324 400556 354325 400620
rect 354259 400555 354325 400556
rect 354262 399941 354322 400555
rect 355182 400213 355242 451283
rect 355179 400212 355245 400213
rect 355179 400148 355180 400212
rect 355244 400148 355245 400212
rect 355179 400147 355245 400148
rect 357390 400077 357450 451555
rect 357571 449444 357637 449445
rect 357571 449380 357572 449444
rect 357636 449380 357637 449444
rect 357571 449379 357637 449380
rect 357574 401029 357634 449379
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 357571 401028 357637 401029
rect 357571 400964 357572 401028
rect 357636 400964 357637 401028
rect 357571 400963 357637 400964
rect 357387 400076 357453 400077
rect 357387 400012 357388 400076
rect 357452 400012 357453 400076
rect 357387 400011 357453 400012
rect 353523 399940 353589 399941
rect 353523 399876 353524 399940
rect 353588 399876 353589 399940
rect 354262 399940 354371 399941
rect 354262 399878 354306 399940
rect 353523 399875 353589 399876
rect 354305 399876 354306 399878
rect 354370 399876 354371 399940
rect 354305 399875 354371 399876
rect 354811 399940 354877 399941
rect 354811 399876 354812 399940
rect 354876 399876 354877 399940
rect 354811 399875 354877 399876
rect 354995 399940 355061 399941
rect 354995 399876 354996 399940
rect 355060 399876 355061 399940
rect 354995 399875 355061 399876
rect 356467 399940 356533 399941
rect 356467 399876 356468 399940
rect 356532 399876 356533 399940
rect 356467 399875 356533 399876
rect 356835 399940 356901 399941
rect 356835 399876 356836 399940
rect 356900 399876 356901 399940
rect 356835 399875 356901 399876
rect 357571 399940 357637 399941
rect 357571 399876 357572 399940
rect 357636 399876 357637 399940
rect 357571 399875 357637 399876
rect 358123 399940 358189 399941
rect 358123 399876 358124 399940
rect 358188 399876 358189 399940
rect 358123 399875 358189 399876
rect 358675 399940 358741 399941
rect 358675 399876 358676 399940
rect 358740 399876 358741 399940
rect 358675 399875 358741 399876
rect 359043 399940 359109 399941
rect 359043 399876 359044 399940
rect 359108 399876 359109 399940
rect 359043 399875 359109 399876
rect 359779 399940 359845 399941
rect 359779 399876 359780 399940
rect 359844 399876 359845 399940
rect 359779 399875 359845 399876
rect 360331 399940 360397 399941
rect 360331 399876 360332 399940
rect 360396 399876 360397 399940
rect 360331 399875 360397 399876
rect 361067 399940 361133 399941
rect 361067 399876 361068 399940
rect 361132 399876 361133 399940
rect 361067 399875 361133 399876
rect 352787 399532 352853 399533
rect 352787 399468 352788 399532
rect 352852 399468 352853 399532
rect 352787 399467 352853 399468
rect 353339 399532 353405 399533
rect 353339 399468 353340 399532
rect 353404 399468 353405 399532
rect 353339 399467 353405 399468
rect 354814 399261 354874 399875
rect 354811 399260 354877 399261
rect 354811 399196 354812 399260
rect 354876 399196 354877 399260
rect 354811 399195 354877 399196
rect 353891 398988 353957 398989
rect 353891 398924 353892 398988
rect 353956 398924 353957 398988
rect 353891 398923 353957 398924
rect 353339 397492 353405 397493
rect 353339 397428 353340 397492
rect 353404 397428 353405 397492
rect 353339 397427 353405 397428
rect 353342 385661 353402 397427
rect 353339 385660 353405 385661
rect 353339 385596 353340 385660
rect 353404 385596 353405 385660
rect 353339 385595 353405 385596
rect 352419 319836 352485 319837
rect 352419 319772 352420 319836
rect 352484 319772 352485 319836
rect 352419 319771 352485 319772
rect 350763 304196 350829 304197
rect 350763 304132 350764 304196
rect 350828 304132 350829 304196
rect 350763 304131 350829 304132
rect 350579 301884 350645 301885
rect 350579 301820 350580 301884
rect 350644 301820 350645 301884
rect 350579 301819 350645 301820
rect 349107 295220 349173 295221
rect 349107 295156 349108 295220
rect 349172 295156 349173 295220
rect 349107 295155 349173 295156
rect 345059 295084 345125 295085
rect 345059 295020 345060 295084
rect 345124 295020 345125 295084
rect 345059 295019 345125 295020
rect 353894 291821 353954 398923
rect 354998 396677 355058 399875
rect 355363 398036 355429 398037
rect 355363 397972 355364 398036
rect 355428 397972 355429 398036
rect 355363 397971 355429 397972
rect 354995 396676 355061 396677
rect 354995 396612 354996 396676
rect 355060 396612 355061 396676
rect 354995 396611 355061 396612
rect 355179 395588 355245 395589
rect 355179 395524 355180 395588
rect 355244 395524 355245 395588
rect 355179 395523 355245 395524
rect 355182 308685 355242 395523
rect 355366 383485 355426 397971
rect 356470 387565 356530 399875
rect 356838 398309 356898 399875
rect 356835 398308 356901 398309
rect 356835 398244 356836 398308
rect 356900 398244 356901 398308
rect 356835 398243 356901 398244
rect 356835 398172 356901 398173
rect 356835 398108 356836 398172
rect 356900 398108 356901 398172
rect 356835 398107 356901 398108
rect 356651 397220 356717 397221
rect 356651 397156 356652 397220
rect 356716 397156 356717 397220
rect 356651 397155 356717 397156
rect 356467 387564 356533 387565
rect 356467 387500 356468 387564
rect 356532 387500 356533 387564
rect 356467 387499 356533 387500
rect 355363 383484 355429 383485
rect 355363 383420 355364 383484
rect 355428 383420 355429 383484
rect 355363 383419 355429 383420
rect 355179 308684 355245 308685
rect 355179 308620 355180 308684
rect 355244 308620 355245 308684
rect 355179 308619 355245 308620
rect 356654 307325 356714 397155
rect 356838 382941 356898 398107
rect 357387 397492 357453 397493
rect 357387 397428 357388 397492
rect 357452 397428 357453 397492
rect 357387 397427 357453 397428
rect 357019 396132 357085 396133
rect 357019 396068 357020 396132
rect 357084 396068 357085 396132
rect 357019 396067 357085 396068
rect 357022 390285 357082 396067
rect 357019 390284 357085 390285
rect 357019 390220 357020 390284
rect 357084 390220 357085 390284
rect 357019 390219 357085 390220
rect 357390 383670 357450 397427
rect 357574 392869 357634 399875
rect 357939 396812 358005 396813
rect 357939 396748 357940 396812
rect 358004 396748 358005 396812
rect 357939 396747 358005 396748
rect 357571 392868 357637 392869
rect 357571 392804 357572 392868
rect 357636 392804 357637 392868
rect 357571 392803 357637 392804
rect 357390 383610 357634 383670
rect 356835 382940 356901 382941
rect 356835 382876 356836 382940
rect 356900 382876 356901 382940
rect 356835 382875 356901 382876
rect 356651 307324 356717 307325
rect 356651 307260 356652 307324
rect 356716 307260 356717 307324
rect 356651 307259 356717 307260
rect 357574 304333 357634 383610
rect 357942 307461 358002 396747
rect 358126 395317 358186 399875
rect 358123 395316 358189 395317
rect 358123 395252 358124 395316
rect 358188 395252 358189 395316
rect 358123 395251 358189 395252
rect 358678 393957 358738 399875
rect 359046 399533 359106 399875
rect 359411 399804 359477 399805
rect 359411 399740 359412 399804
rect 359476 399740 359477 399804
rect 359411 399739 359477 399740
rect 359043 399532 359109 399533
rect 359043 399468 359044 399532
rect 359108 399468 359109 399532
rect 359043 399467 359109 399468
rect 358859 399260 358925 399261
rect 358859 399196 358860 399260
rect 358924 399196 358925 399260
rect 358859 399195 358925 399196
rect 358675 393956 358741 393957
rect 358675 393892 358676 393956
rect 358740 393892 358741 393956
rect 358675 393891 358741 393892
rect 357939 307460 358005 307461
rect 357939 307396 357940 307460
rect 358004 307396 358005 307460
rect 357939 307395 358005 307396
rect 357571 304332 357637 304333
rect 357571 304268 357572 304332
rect 357636 304268 357637 304332
rect 357571 304267 357637 304268
rect 358862 302157 358922 399195
rect 359043 398988 359109 398989
rect 359043 398924 359044 398988
rect 359108 398924 359109 398988
rect 359043 398923 359109 398924
rect 359046 387157 359106 398923
rect 359414 396541 359474 399739
rect 359411 396540 359477 396541
rect 359411 396476 359412 396540
rect 359476 396476 359477 396540
rect 359411 396475 359477 396476
rect 359411 395452 359477 395453
rect 359411 395388 359412 395452
rect 359476 395388 359477 395452
rect 359411 395387 359477 395388
rect 359043 387156 359109 387157
rect 359043 387092 359044 387156
rect 359108 387092 359109 387156
rect 359043 387091 359109 387092
rect 358859 302156 358925 302157
rect 358859 302092 358860 302156
rect 358924 302092 358925 302156
rect 358859 302091 358925 302092
rect 359414 297941 359474 395387
rect 359782 395045 359842 399875
rect 360334 398989 360394 399875
rect 360515 399804 360581 399805
rect 360515 399740 360516 399804
rect 360580 399740 360581 399804
rect 360515 399739 360581 399740
rect 360331 398988 360397 398989
rect 360331 398924 360332 398988
rect 360396 398924 360397 398988
rect 360331 398923 360397 398924
rect 360331 398852 360397 398853
rect 360331 398788 360332 398852
rect 360396 398788 360397 398852
rect 360331 398787 360397 398788
rect 359779 395044 359845 395045
rect 359779 394980 359780 395044
rect 359844 394980 359845 395044
rect 359779 394979 359845 394980
rect 360334 389190 360394 398787
rect 360518 392597 360578 399739
rect 360699 399532 360765 399533
rect 360699 399468 360700 399532
rect 360764 399468 360765 399532
rect 360699 399467 360765 399468
rect 360515 392596 360581 392597
rect 360515 392532 360516 392596
rect 360580 392532 360581 392596
rect 360515 392531 360581 392532
rect 360150 389130 360394 389190
rect 360150 315893 360210 389130
rect 360147 315892 360213 315893
rect 360147 315828 360148 315892
rect 360212 315828 360213 315892
rect 360147 315827 360213 315828
rect 360702 303245 360762 399467
rect 361070 396813 361130 399875
rect 361251 399804 361317 399805
rect 361251 399740 361252 399804
rect 361316 399740 361317 399804
rect 361251 399739 361317 399740
rect 361067 396812 361133 396813
rect 361067 396748 361068 396812
rect 361132 396748 361133 396812
rect 361067 396747 361133 396748
rect 361254 393005 361314 399739
rect 361794 399454 362414 434898
rect 365514 705798 366134 705830
rect 365514 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 366134 705798
rect 365514 705478 366134 705562
rect 365514 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 366134 705478
rect 365514 691174 366134 705242
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 372659 452572 372725 452573
rect 372659 452508 372660 452572
rect 372724 452508 372725 452572
rect 372659 452507 372725 452508
rect 374131 452572 374197 452573
rect 374131 452508 374132 452572
rect 374196 452508 374197 452572
rect 374131 452507 374197 452508
rect 368979 451484 369045 451485
rect 368979 451420 368980 451484
rect 369044 451420 369045 451484
rect 368979 451419 369045 451420
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 363275 399940 363341 399941
rect 363275 399876 363276 399940
rect 363340 399876 363341 399940
rect 363275 399875 363341 399876
rect 363827 399940 363893 399941
rect 363827 399876 363828 399940
rect 363892 399876 363893 399940
rect 363827 399875 363893 399876
rect 364379 399940 364445 399941
rect 364379 399876 364380 399940
rect 364444 399876 364445 399940
rect 364931 399940 364997 399941
rect 364931 399938 364932 399940
rect 364379 399875 364445 399876
rect 364566 399878 364932 399938
rect 362907 399804 362973 399805
rect 362907 399740 362908 399804
rect 362972 399740 362973 399804
rect 362907 399739 362973 399740
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361251 393004 361317 393005
rect 361251 392940 361252 393004
rect 361316 392940 361317 393004
rect 361251 392939 361317 392940
rect 361794 363454 362414 398898
rect 362723 398036 362789 398037
rect 362723 397972 362724 398036
rect 362788 397972 362789 398036
rect 362723 397971 362789 397972
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 360699 303244 360765 303245
rect 360699 303180 360700 303244
rect 360764 303180 360765 303244
rect 360699 303179 360765 303180
rect 359411 297940 359477 297941
rect 359411 297876 359412 297940
rect 359476 297876 359477 297940
rect 359411 297875 359477 297876
rect 353891 291820 353957 291821
rect 353891 291756 353892 291820
rect 353956 291756 353957 291820
rect 353891 291755 353957 291756
rect 353894 277410 353954 291755
rect 353342 277350 353954 277410
rect 361794 291454 362414 326898
rect 362726 319701 362786 397971
rect 362723 319700 362789 319701
rect 362723 319636 362724 319700
rect 362788 319636 362789 319700
rect 362723 319635 362789 319636
rect 362910 304741 362970 399739
rect 363278 395725 363338 399875
rect 363459 398172 363525 398173
rect 363459 398108 363460 398172
rect 363524 398108 363525 398172
rect 363459 398107 363525 398108
rect 363275 395724 363341 395725
rect 363275 395660 363276 395724
rect 363340 395660 363341 395724
rect 363275 395659 363341 395660
rect 362907 304740 362973 304741
rect 362907 304676 362908 304740
rect 362972 304676 362973 304740
rect 362907 304675 362973 304676
rect 363462 304469 363522 398107
rect 363643 397356 363709 397357
rect 363643 397292 363644 397356
rect 363708 397292 363709 397356
rect 363643 397291 363709 397292
rect 363646 388245 363706 397291
rect 363830 394501 363890 399875
rect 364382 395453 364442 399875
rect 364379 395452 364445 395453
rect 364379 395388 364380 395452
rect 364444 395388 364445 395452
rect 364379 395387 364445 395388
rect 364379 395316 364445 395317
rect 364379 395252 364380 395316
rect 364444 395252 364445 395316
rect 364379 395251 364445 395252
rect 363827 394500 363893 394501
rect 363827 394436 363828 394500
rect 363892 394436 363893 394500
rect 363827 394435 363893 394436
rect 363643 388244 363709 388245
rect 363643 388180 363644 388244
rect 363708 388180 363709 388244
rect 363643 388179 363709 388180
rect 363459 304468 363525 304469
rect 363459 304404 363460 304468
rect 363524 304404 363525 304468
rect 363459 304403 363525 304404
rect 364382 298077 364442 395251
rect 364566 383349 364626 399878
rect 364931 399876 364932 399878
rect 364996 399876 364997 399940
rect 364931 399875 364997 399876
rect 364931 399804 364997 399805
rect 364931 399740 364932 399804
rect 364996 399740 364997 399804
rect 364931 399739 364997 399740
rect 365299 399804 365365 399805
rect 365299 399740 365300 399804
rect 365364 399740 365365 399804
rect 365299 399739 365365 399740
rect 364747 398580 364813 398581
rect 364747 398516 364748 398580
rect 364812 398516 364813 398580
rect 364747 398515 364813 398516
rect 364750 397221 364810 398515
rect 364747 397220 364813 397221
rect 364747 397156 364748 397220
rect 364812 397156 364813 397220
rect 364747 397155 364813 397156
rect 364934 395045 364994 399739
rect 365302 397901 365362 399739
rect 365299 397900 365365 397901
rect 365299 397836 365300 397900
rect 365364 397836 365365 397900
rect 365299 397835 365365 397836
rect 364931 395044 364997 395045
rect 364931 394980 364932 395044
rect 364996 394980 364997 395044
rect 364931 394979 364997 394980
rect 364563 383348 364629 383349
rect 364563 383284 364564 383348
rect 364628 383284 364629 383348
rect 364563 383283 364629 383284
rect 365514 367174 366134 402618
rect 368982 401301 369042 451419
rect 372662 449445 372722 452507
rect 374134 449445 374194 452507
rect 375971 451348 376037 451349
rect 375971 451284 375972 451348
rect 376036 451284 376037 451348
rect 375971 451283 376037 451284
rect 370451 449444 370517 449445
rect 370451 449380 370452 449444
rect 370516 449380 370517 449444
rect 370451 449379 370517 449380
rect 371555 449444 371621 449445
rect 371555 449380 371556 449444
rect 371620 449380 371621 449444
rect 371555 449379 371621 449380
rect 372659 449444 372725 449445
rect 372659 449380 372660 449444
rect 372724 449380 372725 449444
rect 372659 449379 372725 449380
rect 374131 449444 374197 449445
rect 374131 449380 374132 449444
rect 374196 449380 374197 449444
rect 374131 449379 374197 449380
rect 368979 401300 369045 401301
rect 368979 401236 368980 401300
rect 369044 401236 369045 401300
rect 368979 401235 369045 401236
rect 368427 400076 368493 400077
rect 368427 400012 368428 400076
rect 368492 400012 368493 400076
rect 368427 400011 368493 400012
rect 368059 399940 368125 399941
rect 368059 399876 368060 399940
rect 368124 399876 368125 399940
rect 368059 399875 368125 399876
rect 366403 399804 366469 399805
rect 366403 399740 366404 399804
rect 366468 399740 366469 399804
rect 366403 399739 366469 399740
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 364379 298076 364445 298077
rect 364379 298012 364380 298076
rect 364444 298012 364445 298076
rect 364379 298011 364445 298012
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 333099 59396 333165 59397
rect 333099 59332 333100 59396
rect 333164 59332 333165 59396
rect 333099 59331 333165 59332
rect 331811 31788 331877 31789
rect 331811 31724 331812 31788
rect 331876 31724 331877 31788
rect 331811 31723 331877 31724
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -1306 330134 6618
rect 353342 3773 353402 277350
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 353339 3772 353405 3773
rect 353339 3708 353340 3772
rect 353404 3708 353405 3772
rect 353339 3707 353405 3708
rect 329514 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 330134 -1306
rect 329514 -1626 330134 -1542
rect 329514 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 330134 -1626
rect 329514 -1894 330134 -1862
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 295174 366134 330618
rect 366406 316981 366466 399739
rect 366587 399532 366653 399533
rect 366587 399468 366588 399532
rect 366652 399468 366653 399532
rect 366587 399467 366653 399468
rect 366590 398717 366650 399467
rect 366587 398716 366653 398717
rect 366587 398652 366588 398716
rect 366652 398652 366653 398716
rect 366587 398651 366653 398652
rect 367323 398172 367389 398173
rect 367323 398108 367324 398172
rect 367388 398108 367389 398172
rect 367323 398107 367389 398108
rect 367691 398172 367757 398173
rect 367691 398108 367692 398172
rect 367756 398108 367757 398172
rect 367691 398107 367757 398108
rect 366587 397356 366653 397357
rect 366587 397292 366588 397356
rect 366652 397292 366653 397356
rect 366587 397291 366653 397292
rect 367139 397356 367205 397357
rect 367139 397292 367140 397356
rect 367204 397292 367205 397356
rect 367139 397291 367205 397292
rect 366590 378997 366650 397291
rect 366587 378996 366653 378997
rect 366587 378932 366588 378996
rect 366652 378932 366653 378996
rect 366587 378931 366653 378932
rect 367142 319565 367202 397291
rect 367326 373285 367386 398107
rect 367323 373284 367389 373285
rect 367323 373220 367324 373284
rect 367388 373220 367389 373284
rect 367323 373219 367389 373220
rect 367139 319564 367205 319565
rect 367139 319500 367140 319564
rect 367204 319500 367205 319564
rect 367139 319499 367205 319500
rect 366403 316980 366469 316981
rect 366403 316916 366404 316980
rect 366468 316916 366469 316980
rect 366403 316915 366469 316916
rect 367694 304605 367754 398107
rect 368062 396133 368122 399875
rect 368243 399804 368309 399805
rect 368243 399740 368244 399804
rect 368308 399740 368309 399804
rect 368243 399739 368309 399740
rect 368246 398037 368306 399739
rect 368243 398036 368309 398037
rect 368243 397972 368244 398036
rect 368308 397972 368309 398036
rect 368243 397971 368309 397972
rect 368059 396132 368125 396133
rect 368059 396068 368060 396132
rect 368124 396068 368125 396132
rect 368059 396067 368125 396068
rect 367691 304604 367757 304605
rect 367691 304540 367692 304604
rect 367756 304540 367757 304604
rect 367691 304539 367757 304540
rect 368430 299437 368490 400011
rect 369163 399940 369229 399941
rect 369163 399876 369164 399940
rect 369228 399876 369229 399940
rect 369163 399875 369229 399876
rect 369531 399940 369597 399941
rect 369531 399876 369532 399940
rect 369596 399876 369597 399940
rect 369531 399875 369597 399876
rect 370083 399940 370149 399941
rect 370083 399876 370084 399940
rect 370148 399876 370149 399940
rect 370083 399875 370149 399876
rect 368611 399804 368677 399805
rect 368611 399740 368612 399804
rect 368676 399740 368677 399804
rect 368611 399739 368677 399740
rect 368614 392733 368674 399739
rect 368979 398036 369045 398037
rect 368979 397972 368980 398036
rect 369044 397972 369045 398036
rect 368979 397971 369045 397972
rect 368611 392732 368677 392733
rect 368611 392668 368612 392732
rect 368676 392668 368677 392732
rect 368611 392667 368677 392668
rect 368982 386069 369042 397971
rect 369166 397629 369226 399875
rect 369534 397901 369594 399875
rect 370086 398717 370146 399875
rect 370454 399533 370514 449379
rect 370635 399940 370701 399941
rect 370635 399876 370636 399940
rect 370700 399876 370701 399940
rect 370635 399875 370701 399876
rect 370451 399532 370517 399533
rect 370451 399468 370452 399532
rect 370516 399468 370517 399532
rect 370451 399467 370517 399468
rect 370083 398716 370149 398717
rect 370083 398652 370084 398716
rect 370148 398652 370149 398716
rect 370083 398651 370149 398652
rect 370083 398580 370149 398581
rect 370083 398516 370084 398580
rect 370148 398516 370149 398580
rect 370083 398515 370149 398516
rect 369531 397900 369597 397901
rect 369531 397836 369532 397900
rect 369596 397836 369597 397900
rect 369531 397835 369597 397836
rect 369899 397900 369965 397901
rect 369899 397836 369900 397900
rect 369964 397836 369965 397900
rect 369899 397835 369965 397836
rect 369163 397628 369229 397629
rect 369163 397564 369164 397628
rect 369228 397564 369229 397628
rect 369163 397563 369229 397564
rect 368979 386068 369045 386069
rect 368979 386004 368980 386068
rect 369044 386004 369045 386068
rect 368979 386003 369045 386004
rect 369902 318069 369962 397835
rect 370086 325277 370146 398515
rect 370638 398445 370698 399875
rect 370635 398444 370701 398445
rect 370635 398380 370636 398444
rect 370700 398380 370701 398444
rect 370635 398379 370701 398380
rect 370267 397764 370333 397765
rect 370267 397700 370268 397764
rect 370332 397700 370333 397764
rect 370267 397699 370333 397700
rect 370270 384301 370330 397699
rect 371371 397492 371437 397493
rect 371371 397428 371372 397492
rect 371436 397428 371437 397492
rect 371371 397427 371437 397428
rect 371374 393957 371434 397427
rect 371371 393956 371437 393957
rect 371371 393892 371372 393956
rect 371436 393892 371437 393956
rect 371371 393891 371437 393892
rect 371558 387701 371618 449379
rect 372662 399125 372722 449379
rect 373947 449308 374013 449309
rect 373947 449306 373948 449308
rect 373766 449246 373948 449306
rect 373766 408510 373826 449246
rect 373947 449244 373948 449246
rect 374012 449244 374013 449308
rect 373947 449243 374013 449244
rect 373766 408450 374010 408510
rect 372843 399396 372909 399397
rect 372843 399332 372844 399396
rect 372908 399332 372909 399396
rect 372843 399331 372909 399332
rect 372659 399124 372725 399125
rect 372659 399060 372660 399124
rect 372724 399060 372725 399124
rect 372659 399059 372725 399060
rect 372659 398308 372725 398309
rect 372659 398244 372660 398308
rect 372724 398244 372725 398308
rect 372659 398243 372725 398244
rect 371555 387700 371621 387701
rect 371555 387636 371556 387700
rect 371620 387636 371621 387700
rect 371555 387635 371621 387636
rect 370267 384300 370333 384301
rect 370267 384236 370268 384300
rect 370332 384236 370333 384300
rect 370267 384235 370333 384236
rect 372662 377637 372722 398243
rect 372846 397901 372906 399331
rect 372843 397900 372909 397901
rect 372843 397836 372844 397900
rect 372908 397836 372909 397900
rect 372843 397835 372909 397836
rect 373211 397492 373277 397493
rect 373211 397428 373212 397492
rect 373276 397428 373277 397492
rect 373211 397427 373277 397428
rect 372659 377636 372725 377637
rect 372659 377572 372660 377636
rect 372724 377572 372725 377636
rect 372659 377571 372725 377572
rect 370083 325276 370149 325277
rect 370083 325212 370084 325276
rect 370148 325212 370149 325276
rect 370083 325211 370149 325212
rect 369899 318068 369965 318069
rect 369899 318004 369900 318068
rect 369964 318004 369965 318068
rect 369899 318003 369965 318004
rect 373214 303381 373274 397427
rect 373950 396677 374010 408450
rect 374134 400077 374194 449379
rect 375974 401165 376034 451283
rect 382227 449444 382293 449445
rect 382227 449380 382228 449444
rect 382292 449380 382293 449444
rect 382227 449379 382293 449380
rect 383883 449444 383949 449445
rect 383883 449380 383884 449444
rect 383948 449380 383949 449444
rect 383883 449379 383949 449380
rect 384251 449444 384317 449445
rect 384251 449380 384252 449444
rect 384316 449380 384317 449444
rect 384251 449379 384317 449380
rect 385355 449444 385421 449445
rect 385355 449380 385356 449444
rect 385420 449380 385421 449444
rect 385355 449379 385421 449380
rect 375971 401164 376037 401165
rect 375971 401100 375972 401164
rect 376036 401100 376037 401164
rect 375971 401099 376037 401100
rect 381307 400348 381373 400349
rect 381307 400284 381308 400348
rect 381372 400284 381373 400348
rect 381307 400283 381373 400284
rect 374131 400076 374197 400077
rect 374131 400012 374132 400076
rect 374196 400012 374197 400076
rect 374131 400011 374197 400012
rect 376523 400076 376589 400077
rect 376523 400012 376524 400076
rect 376588 400012 376589 400076
rect 376523 400011 376589 400012
rect 377259 400076 377325 400077
rect 377259 400012 377260 400076
rect 377324 400012 377325 400076
rect 377259 400011 377325 400012
rect 375051 399940 375117 399941
rect 375051 399876 375052 399940
rect 375116 399876 375117 399940
rect 375051 399875 375117 399876
rect 375787 399940 375853 399941
rect 375787 399876 375788 399940
rect 375852 399876 375853 399940
rect 375787 399875 375853 399876
rect 374499 398852 374565 398853
rect 374499 398788 374500 398852
rect 374564 398788 374565 398852
rect 374499 398787 374565 398788
rect 373947 396676 374013 396677
rect 373947 396612 373948 396676
rect 374012 396612 374013 396676
rect 373947 396611 374013 396612
rect 374502 392189 374562 398787
rect 375054 395317 375114 399875
rect 375790 396949 375850 399875
rect 375787 396948 375853 396949
rect 375787 396884 375788 396948
rect 375852 396884 375853 396948
rect 375787 396883 375853 396884
rect 375051 395316 375117 395317
rect 375051 395252 375052 395316
rect 375116 395252 375117 395316
rect 375051 395251 375117 395252
rect 374499 392188 374565 392189
rect 374499 392124 374500 392188
rect 374564 392124 374565 392188
rect 374499 392123 374565 392124
rect 375419 391372 375485 391373
rect 375419 391308 375420 391372
rect 375484 391308 375485 391372
rect 375419 391307 375485 391308
rect 373211 303380 373277 303381
rect 373211 303316 373212 303380
rect 373276 303316 373277 303380
rect 373211 303315 373277 303316
rect 368427 299436 368493 299437
rect 368427 299372 368428 299436
rect 368492 299372 368493 299436
rect 368427 299371 368493 299372
rect 375422 299165 375482 391307
rect 376526 338197 376586 400011
rect 376707 399940 376773 399941
rect 376707 399876 376708 399940
rect 376772 399876 376773 399940
rect 376707 399875 376773 399876
rect 376710 398445 376770 399875
rect 376891 399396 376957 399397
rect 376891 399332 376892 399396
rect 376956 399332 376957 399396
rect 376891 399331 376957 399332
rect 376707 398444 376773 398445
rect 376707 398380 376708 398444
rect 376772 398380 376773 398444
rect 376707 398379 376773 398380
rect 376523 338196 376589 338197
rect 376523 338132 376524 338196
rect 376588 338132 376589 338196
rect 376523 338131 376589 338132
rect 376526 335370 376586 338131
rect 375974 335310 376586 335370
rect 375974 309909 376034 335310
rect 375971 309908 376037 309909
rect 375971 309844 375972 309908
rect 376036 309844 376037 309908
rect 375971 309843 376037 309844
rect 376894 299301 376954 399331
rect 377262 305965 377322 400011
rect 378731 399940 378797 399941
rect 378731 399876 378732 399940
rect 378796 399876 378797 399940
rect 378731 399875 378797 399876
rect 380203 399940 380269 399941
rect 380203 399876 380204 399940
rect 380268 399876 380269 399940
rect 380203 399875 380269 399876
rect 381077 399940 381143 399941
rect 381077 399876 381078 399940
rect 381142 399938 381143 399940
rect 381142 399876 381186 399938
rect 381077 399875 381186 399876
rect 378179 399260 378245 399261
rect 378179 399196 378180 399260
rect 378244 399196 378245 399260
rect 378179 399195 378245 399196
rect 378182 321061 378242 399195
rect 378363 397492 378429 397493
rect 378363 397428 378364 397492
rect 378428 397428 378429 397492
rect 378363 397427 378429 397428
rect 378366 325141 378426 397427
rect 378734 395317 378794 399875
rect 378915 399804 378981 399805
rect 378915 399740 378916 399804
rect 378980 399740 378981 399804
rect 378915 399739 378981 399740
rect 378918 395317 378978 399739
rect 379651 399260 379717 399261
rect 379651 399196 379652 399260
rect 379716 399196 379717 399260
rect 379651 399195 379717 399196
rect 378731 395316 378797 395317
rect 378731 395252 378732 395316
rect 378796 395252 378797 395316
rect 378731 395251 378797 395252
rect 378915 395316 378981 395317
rect 378915 395252 378916 395316
rect 378980 395252 378981 395316
rect 378915 395251 378981 395252
rect 379654 389190 379714 399195
rect 380206 396949 380266 399875
rect 380755 398716 380821 398717
rect 380755 398652 380756 398716
rect 380820 398652 380821 398716
rect 380755 398651 380821 398652
rect 380203 396948 380269 396949
rect 380203 396884 380204 396948
rect 380268 396884 380269 396948
rect 380203 396883 380269 396884
rect 379470 389130 379714 389190
rect 378363 325140 378429 325141
rect 378363 325076 378364 325140
rect 378428 325076 378429 325140
rect 378363 325075 378429 325076
rect 378179 321060 378245 321061
rect 378179 320996 378180 321060
rect 378244 320996 378245 321060
rect 378179 320995 378245 320996
rect 377259 305964 377325 305965
rect 377259 305900 377260 305964
rect 377324 305900 377325 305964
rect 377259 305899 377325 305900
rect 379470 304877 379530 389130
rect 380758 335477 380818 398651
rect 380939 397492 381005 397493
rect 380939 397428 380940 397492
rect 381004 397428 381005 397492
rect 380939 397427 381005 397428
rect 380755 335476 380821 335477
rect 380755 335412 380756 335476
rect 380820 335412 380821 335476
rect 380755 335411 380821 335412
rect 380758 334661 380818 335411
rect 380755 334660 380821 334661
rect 380755 334596 380756 334660
rect 380820 334596 380821 334660
rect 380755 334595 380821 334596
rect 380942 311405 381002 397427
rect 381126 393549 381186 399875
rect 381310 399669 381370 400283
rect 381491 399940 381557 399941
rect 381491 399876 381492 399940
rect 381556 399876 381557 399940
rect 381491 399875 381557 399876
rect 381307 399668 381373 399669
rect 381307 399604 381308 399668
rect 381372 399604 381373 399668
rect 381307 399603 381373 399604
rect 381494 398717 381554 399875
rect 382230 399805 382290 449379
rect 382963 449308 383029 449309
rect 382963 449244 382964 449308
rect 383028 449244 383029 449308
rect 382963 449243 383029 449244
rect 382227 399804 382293 399805
rect 382227 399740 382228 399804
rect 382292 399740 382293 399804
rect 382227 399739 382293 399740
rect 381675 399668 381741 399669
rect 381675 399604 381676 399668
rect 381740 399604 381741 399668
rect 381675 399603 381741 399604
rect 381491 398716 381557 398717
rect 381491 398652 381492 398716
rect 381556 398652 381557 398716
rect 381491 398651 381557 398652
rect 381678 394710 381738 399603
rect 382779 397900 382845 397901
rect 382779 397836 382780 397900
rect 382844 397836 382845 397900
rect 382779 397835 382845 397836
rect 382227 397628 382293 397629
rect 382227 397564 382228 397628
rect 382292 397564 382293 397628
rect 382227 397563 382293 397564
rect 381494 394650 381738 394710
rect 381123 393548 381189 393549
rect 381123 393484 381124 393548
rect 381188 393484 381189 393548
rect 381123 393483 381189 393484
rect 380939 311404 381005 311405
rect 380939 311340 380940 311404
rect 381004 311340 381005 311404
rect 380939 311339 381005 311340
rect 379467 304876 379533 304877
rect 379467 304812 379468 304876
rect 379532 304812 379533 304876
rect 379467 304811 379533 304812
rect 381494 300661 381554 394650
rect 382230 325005 382290 397563
rect 382227 325004 382293 325005
rect 382227 324940 382228 325004
rect 382292 324940 382293 325004
rect 382227 324939 382293 324940
rect 382782 315621 382842 397835
rect 382966 385797 383026 449243
rect 383699 398444 383765 398445
rect 383699 398380 383700 398444
rect 383764 398380 383765 398444
rect 383699 398379 383765 398380
rect 382963 385796 383029 385797
rect 382963 385732 382964 385796
rect 383028 385732 383029 385796
rect 382963 385731 383029 385732
rect 382779 315620 382845 315621
rect 382779 315556 382780 315620
rect 382844 315556 382845 315620
rect 382779 315555 382845 315556
rect 383702 302021 383762 398379
rect 383886 389061 383946 449379
rect 384254 408510 384314 449379
rect 384254 408450 384498 408510
rect 384438 399261 384498 408450
rect 384987 400076 385053 400077
rect 384987 400012 384988 400076
rect 385052 400012 385053 400076
rect 384987 400011 385053 400012
rect 384435 399260 384501 399261
rect 384435 399196 384436 399260
rect 384500 399196 384501 399260
rect 384435 399195 384501 399196
rect 383883 389060 383949 389061
rect 383883 388996 383884 389060
rect 383948 388996 383949 389060
rect 383883 388995 383949 388996
rect 384990 307597 385050 400011
rect 385171 396132 385237 396133
rect 385171 396068 385172 396132
rect 385236 396068 385237 396132
rect 385171 396067 385237 396068
rect 385174 322285 385234 396067
rect 385358 388517 385418 449379
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 385723 400484 385789 400485
rect 385723 400420 385724 400484
rect 385788 400420 385789 400484
rect 385723 400419 385789 400420
rect 385726 399669 385786 400419
rect 385723 399668 385789 399669
rect 385723 399604 385724 399668
rect 385788 399604 385789 399668
rect 385723 399603 385789 399604
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 385355 388516 385421 388517
rect 385355 388452 385356 388516
rect 385420 388452 385421 388516
rect 385355 388451 385421 388452
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 385171 322284 385237 322285
rect 385171 322220 385172 322284
rect 385236 322220 385237 322284
rect 385171 322219 385237 322220
rect 384987 307596 385053 307597
rect 384987 307532 384988 307596
rect 385052 307532 385053 307596
rect 384987 307531 385053 307532
rect 383699 302020 383765 302021
rect 383699 301956 383700 302020
rect 383764 301956 383765 302020
rect 383699 301955 383765 301956
rect 381491 300660 381557 300661
rect 381491 300596 381492 300660
rect 381556 300596 381557 300660
rect 381491 300595 381557 300596
rect 376891 299300 376957 299301
rect 376891 299236 376892 299300
rect 376956 299236 376957 299300
rect 376891 299235 376957 299236
rect 375419 299164 375485 299165
rect 375419 299100 375420 299164
rect 375484 299100 375485 299164
rect 375419 299099 375485 299100
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -1306 366134 6618
rect 365514 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 366134 -1306
rect 365514 -1626 366134 -1542
rect 365514 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 366134 -1626
rect 365514 -1894 366134 -1862
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 705798 402134 705830
rect 401514 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 402134 705798
rect 401514 705478 402134 705562
rect 401514 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 402134 705478
rect 401514 691174 402134 705242
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -1306 402134 6618
rect 401514 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 402134 -1306
rect 401514 -1626 402134 -1542
rect 401514 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 402134 -1626
rect 401514 -1894 402134 -1862
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 705798 438134 705830
rect 437514 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 438134 705798
rect 437514 705478 438134 705562
rect 437514 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 438134 705478
rect 437514 691174 438134 705242
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 151174 438134 186618
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 115174 438134 150618
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -1306 438134 6618
rect 437514 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 438134 -1306
rect 437514 -1626 438134 -1542
rect 437514 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 438134 -1626
rect 437514 -1894 438134 -1862
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 705798 474134 705830
rect 473514 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 474134 705798
rect 473514 705478 474134 705562
rect 473514 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 474134 705478
rect 473514 691174 474134 705242
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -1306 474134 6618
rect 473514 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 474134 -1306
rect 473514 -1626 474134 -1542
rect 473514 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 474134 -1626
rect 473514 -1894 474134 -1862
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 705798 510134 705830
rect 509514 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 510134 705798
rect 509514 705478 510134 705562
rect 509514 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 510134 705478
rect 509514 691174 510134 705242
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -1306 510134 6618
rect 509514 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 510134 -1306
rect 509514 -1626 510134 -1542
rect 509514 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 510134 -1626
rect 509514 -1894 510134 -1862
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 705798 546134 705830
rect 545514 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 546134 705798
rect 545514 705478 546134 705562
rect 545514 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 546134 705478
rect 545514 691174 546134 705242
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -1306 546134 6618
rect 545514 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 546134 -1306
rect 545514 -1626 546134 -1542
rect 545514 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 546134 -1626
rect 545514 -1894 546134 -1862
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 705798 582134 705830
rect 581514 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 582134 705798
rect 581514 705478 582134 705562
rect 581514 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 582134 705478
rect 581514 691174 582134 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -1306 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691174 586890 705242
rect 586270 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 586890 691174
rect 586270 690854 586890 690938
rect 586270 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 586890 690854
rect 586270 655174 586890 690618
rect 586270 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 586890 655174
rect 586270 654854 586890 654938
rect 586270 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 586890 654854
rect 586270 619174 586890 654618
rect 586270 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 586890 619174
rect 586270 618854 586890 618938
rect 586270 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 586890 618854
rect 586270 583174 586890 618618
rect 586270 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 586890 583174
rect 586270 582854 586890 582938
rect 586270 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 586890 582854
rect 586270 547174 586890 582618
rect 586270 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 586890 547174
rect 586270 546854 586890 546938
rect 586270 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 586890 546854
rect 586270 511174 586890 546618
rect 586270 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 586890 511174
rect 586270 510854 586890 510938
rect 586270 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 586890 510854
rect 586270 475174 586890 510618
rect 586270 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 586890 475174
rect 586270 474854 586890 474938
rect 586270 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 586890 474854
rect 586270 439174 586890 474618
rect 586270 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 586890 439174
rect 586270 438854 586890 438938
rect 586270 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 586890 438854
rect 586270 403174 586890 438618
rect 586270 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 586890 403174
rect 586270 402854 586890 402938
rect 586270 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 586890 402854
rect 586270 367174 586890 402618
rect 586270 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 586890 367174
rect 586270 366854 586890 366938
rect 586270 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 586890 366854
rect 586270 331174 586890 366618
rect 586270 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 586890 331174
rect 586270 330854 586890 330938
rect 586270 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 586890 330854
rect 586270 295174 586890 330618
rect 586270 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 586890 295174
rect 586270 294854 586890 294938
rect 586270 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 586890 294854
rect 586270 259174 586890 294618
rect 586270 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 586890 259174
rect 586270 258854 586890 258938
rect 586270 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 586890 258854
rect 586270 223174 586890 258618
rect 586270 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 586890 223174
rect 586270 222854 586890 222938
rect 586270 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 586890 222854
rect 586270 187174 586890 222618
rect 586270 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 586890 187174
rect 586270 186854 586890 186938
rect 586270 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 586890 186854
rect 586270 151174 586890 186618
rect 586270 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 586890 151174
rect 586270 150854 586890 150938
rect 586270 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 586890 150854
rect 586270 115174 586890 150618
rect 586270 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 586890 115174
rect 586270 114854 586890 114938
rect 586270 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 586890 114854
rect 586270 79174 586890 114618
rect 586270 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 586890 79174
rect 586270 78854 586890 78938
rect 586270 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 586890 78854
rect 586270 43174 586890 78618
rect 586270 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 586890 43174
rect 586270 42854 586890 42938
rect 586270 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 586890 42854
rect 586270 7174 586890 42618
rect 586270 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 586890 7174
rect 586270 6854 586890 6938
rect 586270 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 586890 6854
rect 581514 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 582134 -1306
rect 581514 -1626 582134 -1542
rect 581514 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 582134 -1626
rect 581514 -1894 582134 -1862
rect 586270 -1306 586890 6618
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
<< via4 >>
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 690938 -2698 691174
rect -2614 690938 -2378 691174
rect -2934 690618 -2698 690854
rect -2614 690618 -2378 690854
rect -2934 654938 -2698 655174
rect -2614 654938 -2378 655174
rect -2934 654618 -2698 654854
rect -2614 654618 -2378 654854
rect -2934 618938 -2698 619174
rect -2614 618938 -2378 619174
rect -2934 618618 -2698 618854
rect -2614 618618 -2378 618854
rect -2934 582938 -2698 583174
rect -2614 582938 -2378 583174
rect -2934 582618 -2698 582854
rect -2614 582618 -2378 582854
rect -2934 546938 -2698 547174
rect -2614 546938 -2378 547174
rect -2934 546618 -2698 546854
rect -2614 546618 -2378 546854
rect -2934 510938 -2698 511174
rect -2614 510938 -2378 511174
rect -2934 510618 -2698 510854
rect -2614 510618 -2378 510854
rect -2934 474938 -2698 475174
rect -2614 474938 -2378 475174
rect -2934 474618 -2698 474854
rect -2614 474618 -2378 474854
rect -2934 438938 -2698 439174
rect -2614 438938 -2378 439174
rect -2934 438618 -2698 438854
rect -2614 438618 -2378 438854
rect -2934 402938 -2698 403174
rect -2614 402938 -2378 403174
rect -2934 402618 -2698 402854
rect -2614 402618 -2378 402854
rect -2934 366938 -2698 367174
rect -2614 366938 -2378 367174
rect -2934 366618 -2698 366854
rect -2614 366618 -2378 366854
rect -2934 330938 -2698 331174
rect -2614 330938 -2378 331174
rect -2934 330618 -2698 330854
rect -2614 330618 -2378 330854
rect -2934 294938 -2698 295174
rect -2614 294938 -2378 295174
rect -2934 294618 -2698 294854
rect -2614 294618 -2378 294854
rect -2934 258938 -2698 259174
rect -2614 258938 -2378 259174
rect -2934 258618 -2698 258854
rect -2614 258618 -2378 258854
rect -2934 222938 -2698 223174
rect -2614 222938 -2378 223174
rect -2934 222618 -2698 222854
rect -2614 222618 -2378 222854
rect -2934 186938 -2698 187174
rect -2614 186938 -2378 187174
rect -2934 186618 -2698 186854
rect -2614 186618 -2378 186854
rect -2934 150938 -2698 151174
rect -2614 150938 -2378 151174
rect -2934 150618 -2698 150854
rect -2614 150618 -2378 150854
rect -2934 114938 -2698 115174
rect -2614 114938 -2378 115174
rect -2934 114618 -2698 114854
rect -2614 114618 -2378 114854
rect -2934 78938 -2698 79174
rect -2614 78938 -2378 79174
rect -2934 78618 -2698 78854
rect -2614 78618 -2378 78854
rect -2934 42938 -2698 43174
rect -2614 42938 -2378 43174
rect -2934 42618 -2698 42854
rect -2614 42618 -2378 42854
rect -2934 6938 -2698 7174
rect -2614 6938 -2378 7174
rect -2934 6618 -2698 6854
rect -2614 6618 -2378 6854
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 705562 5782 705798
rect 5866 705562 6102 705798
rect 5546 705242 5782 705478
rect 5866 705242 6102 705478
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect 5546 -1542 5782 -1306
rect 5866 -1542 6102 -1306
rect 5546 -1862 5782 -1626
rect 5866 -1862 6102 -1626
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 705562 41782 705798
rect 41866 705562 42102 705798
rect 41546 705242 41782 705478
rect 41866 705242 42102 705478
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -1542 41782 -1306
rect 41866 -1542 42102 -1306
rect 41546 -1862 41782 -1626
rect 41866 -1862 42102 -1626
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 705562 77782 705798
rect 77866 705562 78102 705798
rect 77546 705242 77782 705478
rect 77866 705242 78102 705478
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 77546 582938 77782 583174
rect 77866 582938 78102 583174
rect 77546 582618 77782 582854
rect 77866 582618 78102 582854
rect 77546 546938 77782 547174
rect 77866 546938 78102 547174
rect 77546 546618 77782 546854
rect 77866 546618 78102 546854
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 77546 438938 77782 439174
rect 77866 438938 78102 439174
rect 77546 438618 77782 438854
rect 77866 438618 78102 438854
rect 77546 402938 77782 403174
rect 77866 402938 78102 403174
rect 77546 402618 77782 402854
rect 77866 402618 78102 402854
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 77546 258938 77782 259174
rect 77866 258938 78102 259174
rect 77546 258618 77782 258854
rect 77866 258618 78102 258854
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 77546 150938 77782 151174
rect 77866 150938 78102 151174
rect 77546 150618 77782 150854
rect 77866 150618 78102 150854
rect 77546 114938 77782 115174
rect 77866 114938 78102 115174
rect 77546 114618 77782 114854
rect 77866 114618 78102 114854
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -1542 77782 -1306
rect 77866 -1542 78102 -1306
rect 77546 -1862 77782 -1626
rect 77866 -1862 78102 -1626
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 705562 113782 705798
rect 113866 705562 114102 705798
rect 113546 705242 113782 705478
rect 113866 705242 114102 705478
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 113546 402938 113782 403174
rect 113866 402938 114102 403174
rect 113546 402618 113782 402854
rect 113866 402618 114102 402854
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 113546 258938 113782 259174
rect 113866 258938 114102 259174
rect 113546 258618 113782 258854
rect 113866 258618 114102 258854
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 113546 150938 113782 151174
rect 113866 150938 114102 151174
rect 113546 150618 113782 150854
rect 113866 150618 114102 150854
rect 113546 114938 113782 115174
rect 113866 114938 114102 115174
rect 113546 114618 113782 114854
rect 113866 114618 114102 114854
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -1542 113782 -1306
rect 113866 -1542 114102 -1306
rect 113546 -1862 113782 -1626
rect 113866 -1862 114102 -1626
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 705562 149782 705798
rect 149866 705562 150102 705798
rect 149546 705242 149782 705478
rect 149866 705242 150102 705478
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 149546 150938 149782 151174
rect 149866 150938 150102 151174
rect 149546 150618 149782 150854
rect 149866 150618 150102 150854
rect 149546 114938 149782 115174
rect 149866 114938 150102 115174
rect 149546 114618 149782 114854
rect 149866 114618 150102 114854
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 164250 183218 164486 183454
rect 164250 182898 164486 183134
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 179610 186938 179846 187174
rect 179610 186618 179846 186854
rect 185546 705562 185782 705798
rect 185866 705562 186102 705798
rect 185546 705242 185782 705478
rect 185866 705242 186102 705478
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 221546 705562 221782 705798
rect 221866 705562 222102 705798
rect 221546 705242 221782 705478
rect 221866 705242 222102 705478
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 221546 438938 221782 439174
rect 221866 438938 222102 439174
rect 221546 438618 221782 438854
rect 221866 438618 222102 438854
rect 221546 402938 221782 403174
rect 221866 402938 222102 403174
rect 221546 402618 221782 402854
rect 221866 402618 222102 402854
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -1542 149782 -1306
rect 149866 -1542 150102 -1306
rect 149546 -1862 149782 -1626
rect 149866 -1862 150102 -1626
rect 185546 222938 185782 223174
rect 185866 222938 186102 223174
rect 185546 222618 185782 222854
rect 185866 222618 186102 222854
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 194970 183218 195206 183454
rect 194970 182898 195206 183134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 221546 330938 221782 331174
rect 221866 330938 222102 331174
rect 221546 330618 221782 330854
rect 221866 330618 222102 330854
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 221546 294938 221782 295174
rect 221866 294938 222102 295174
rect 221546 294618 221782 294854
rect 221866 294618 222102 294854
rect 221546 258938 221782 259174
rect 221866 258938 222102 259174
rect 221546 258618 221782 258854
rect 221866 258618 222102 258854
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 185546 -1542 185782 -1306
rect 185866 -1542 186102 -1306
rect 185546 -1862 185782 -1626
rect 185866 -1862 186102 -1626
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 222938 221782 223174
rect 221866 222938 222102 223174
rect 221546 222618 221782 222854
rect 221866 222618 222102 222854
rect 221546 186938 221782 187174
rect 221866 186938 222102 187174
rect 221546 186618 221782 186854
rect 221866 186618 222102 186854
rect 221546 150938 221782 151174
rect 221866 150938 222102 151174
rect 221546 150618 221782 150854
rect 221866 150618 222102 150854
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 257546 705562 257782 705798
rect 257866 705562 258102 705798
rect 257546 705242 257782 705478
rect 257866 705242 258102 705478
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 257546 438938 257782 439174
rect 257866 438938 258102 439174
rect 257546 438618 257782 438854
rect 257866 438618 258102 438854
rect 257546 402938 257782 403174
rect 257866 402938 258102 403174
rect 257546 402618 257782 402854
rect 257866 402618 258102 402854
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 257546 330938 257782 331174
rect 257866 330938 258102 331174
rect 257546 330618 257782 330854
rect 257866 330618 258102 330854
rect 257546 294938 257782 295174
rect 257866 294938 258102 295174
rect 257546 294618 257782 294854
rect 257866 294618 258102 294854
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 221546 114938 221782 115174
rect 221866 114938 222102 115174
rect 221546 114618 221782 114854
rect 221866 114618 222102 114854
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -1542 221782 -1306
rect 221866 -1542 222102 -1306
rect 221546 -1862 221782 -1626
rect 221866 -1862 222102 -1626
rect 257546 258938 257782 259174
rect 257866 258938 258102 259174
rect 257546 258618 257782 258854
rect 257866 258618 258102 258854
rect 257546 222938 257782 223174
rect 257866 222938 258102 223174
rect 257546 222618 257782 222854
rect 257866 222618 258102 222854
rect 257546 186938 257782 187174
rect 257866 186938 258102 187174
rect 257546 186618 257782 186854
rect 257866 186618 258102 186854
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 293546 705562 293782 705798
rect 293866 705562 294102 705798
rect 293546 705242 293782 705478
rect 293866 705242 294102 705478
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 293546 438938 293782 439174
rect 293866 438938 294102 439174
rect 293546 438618 293782 438854
rect 293866 438618 294102 438854
rect 293546 402938 293782 403174
rect 293866 402938 294102 403174
rect 293546 402618 293782 402854
rect 293866 402618 294102 402854
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 293546 330938 293782 331174
rect 293866 330938 294102 331174
rect 293546 330618 293782 330854
rect 293866 330618 294102 330854
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 293546 294938 293782 295174
rect 293866 294938 294102 295174
rect 293546 294618 293782 294854
rect 293866 294618 294102 294854
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 293546 222938 293782 223174
rect 293866 222938 294102 223174
rect 293546 222618 293782 222854
rect 293866 222618 294102 222854
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -1542 257782 -1306
rect 257866 -1542 258102 -1306
rect 257546 -1862 257782 -1626
rect 257866 -1862 258102 -1626
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 329546 705562 329782 705798
rect 329866 705562 330102 705798
rect 329546 705242 329782 705478
rect 329866 705242 330102 705478
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 329546 438938 329782 439174
rect 329866 438938 330102 439174
rect 329546 438618 329782 438854
rect 329866 438618 330102 438854
rect 329546 402938 329782 403174
rect 329866 402938 330102 403174
rect 329546 402618 329782 402854
rect 329866 402618 330102 402854
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 329546 330938 329782 331174
rect 329866 330938 330102 331174
rect 329546 330618 329782 330854
rect 329866 330618 330102 330854
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 293546 186938 293782 187174
rect 293866 186938 294102 187174
rect 293546 186618 293782 186854
rect 293866 186618 294102 186854
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -1542 293782 -1306
rect 293866 -1542 294102 -1306
rect 293546 -1862 293782 -1626
rect 293866 -1862 294102 -1626
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 365546 705562 365782 705798
rect 365866 705562 366102 705798
rect 365546 705242 365782 705478
rect 365866 705242 366102 705478
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 329546 -1542 329782 -1306
rect 329866 -1542 330102 -1306
rect 329546 -1862 329782 -1626
rect 329866 -1862 330102 -1626
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -1542 365782 -1306
rect 365866 -1542 366102 -1306
rect 365546 -1862 365782 -1626
rect 365866 -1862 366102 -1626
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 705562 401782 705798
rect 401866 705562 402102 705798
rect 401546 705242 401782 705478
rect 401866 705242 402102 705478
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -1542 401782 -1306
rect 401866 -1542 402102 -1306
rect 401546 -1862 401782 -1626
rect 401866 -1862 402102 -1626
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 705562 437782 705798
rect 437866 705562 438102 705798
rect 437546 705242 437782 705478
rect 437866 705242 438102 705478
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -1542 437782 -1306
rect 437866 -1542 438102 -1306
rect 437546 -1862 437782 -1626
rect 437866 -1862 438102 -1626
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 705562 473782 705798
rect 473866 705562 474102 705798
rect 473546 705242 473782 705478
rect 473866 705242 474102 705478
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -1542 473782 -1306
rect 473866 -1542 474102 -1306
rect 473546 -1862 473782 -1626
rect 473866 -1862 474102 -1626
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 705562 509782 705798
rect 509866 705562 510102 705798
rect 509546 705242 509782 705478
rect 509866 705242 510102 705478
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -1542 509782 -1306
rect 509866 -1542 510102 -1306
rect 509546 -1862 509782 -1626
rect 509866 -1862 510102 -1626
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 705562 545782 705798
rect 545866 705562 546102 705798
rect 545546 705242 545782 705478
rect 545866 705242 546102 705478
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -1542 545782 -1306
rect 545866 -1542 546102 -1306
rect 545546 -1862 545782 -1626
rect 545866 -1862 546102 -1626
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 581546 705562 581782 705798
rect 581866 705562 582102 705798
rect 581546 705242 581782 705478
rect 581866 705242 582102 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 690938 586538 691174
rect 586622 690938 586858 691174
rect 586302 690618 586538 690854
rect 586622 690618 586858 690854
rect 586302 654938 586538 655174
rect 586622 654938 586858 655174
rect 586302 654618 586538 654854
rect 586622 654618 586858 654854
rect 586302 618938 586538 619174
rect 586622 618938 586858 619174
rect 586302 618618 586538 618854
rect 586622 618618 586858 618854
rect 586302 582938 586538 583174
rect 586622 582938 586858 583174
rect 586302 582618 586538 582854
rect 586622 582618 586858 582854
rect 586302 546938 586538 547174
rect 586622 546938 586858 547174
rect 586302 546618 586538 546854
rect 586622 546618 586858 546854
rect 586302 510938 586538 511174
rect 586622 510938 586858 511174
rect 586302 510618 586538 510854
rect 586622 510618 586858 510854
rect 586302 474938 586538 475174
rect 586622 474938 586858 475174
rect 586302 474618 586538 474854
rect 586622 474618 586858 474854
rect 586302 438938 586538 439174
rect 586622 438938 586858 439174
rect 586302 438618 586538 438854
rect 586622 438618 586858 438854
rect 586302 402938 586538 403174
rect 586622 402938 586858 403174
rect 586302 402618 586538 402854
rect 586622 402618 586858 402854
rect 586302 366938 586538 367174
rect 586622 366938 586858 367174
rect 586302 366618 586538 366854
rect 586622 366618 586858 366854
rect 586302 330938 586538 331174
rect 586622 330938 586858 331174
rect 586302 330618 586538 330854
rect 586622 330618 586858 330854
rect 586302 294938 586538 295174
rect 586622 294938 586858 295174
rect 586302 294618 586538 294854
rect 586622 294618 586858 294854
rect 586302 258938 586538 259174
rect 586622 258938 586858 259174
rect 586302 258618 586538 258854
rect 586622 258618 586858 258854
rect 586302 222938 586538 223174
rect 586622 222938 586858 223174
rect 586302 222618 586538 222854
rect 586622 222618 586858 222854
rect 586302 186938 586538 187174
rect 586622 186938 586858 187174
rect 586302 186618 586538 186854
rect 586622 186618 586858 186854
rect 586302 150938 586538 151174
rect 586622 150938 586858 151174
rect 586302 150618 586538 150854
rect 586622 150618 586858 150854
rect 586302 114938 586538 115174
rect 586622 114938 586858 115174
rect 586302 114618 586538 114854
rect 586622 114618 586858 114854
rect 586302 78938 586538 79174
rect 586622 78938 586858 79174
rect 586302 78618 586538 78854
rect 586622 78618 586858 78854
rect 586302 42938 586538 43174
rect 586622 42938 586858 43174
rect 586302 42618 586538 42854
rect 586622 42618 586858 42854
rect 586302 6938 586538 7174
rect 586622 6938 586858 7174
rect 586302 6618 586538 6854
rect 586622 6618 586858 6854
rect 581546 -1542 581782 -1306
rect 581866 -1542 582102 -1306
rect 581546 -1862 581782 -1626
rect 581866 -1862 582102 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
<< metal5 >>
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -2966 691174 586890 691206
rect -2966 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 586890 691174
rect -2966 690854 586890 690938
rect -2966 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 586890 690854
rect -2966 690586 586890 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -2966 655174 586890 655206
rect -2966 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 586890 655174
rect -2966 654854 586890 654938
rect -2966 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 586890 654854
rect -2966 654586 586890 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -2966 619174 586890 619206
rect -2966 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 586890 619174
rect -2966 618854 586890 618938
rect -2966 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 586890 618854
rect -2966 618586 586890 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -2966 583174 586890 583206
rect -2966 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 586890 583174
rect -2966 582854 586890 582938
rect -2966 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 586890 582854
rect -2966 582586 586890 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -2966 547174 586890 547206
rect -2966 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 586890 547174
rect -2966 546854 586890 546938
rect -2966 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 586890 546854
rect -2966 546586 586890 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -2966 511174 586890 511206
rect -2966 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 586890 511174
rect -2966 510854 586890 510938
rect -2966 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 586890 510854
rect -2966 510586 586890 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -2966 475174 586890 475206
rect -2966 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 586890 475174
rect -2966 474854 586890 474938
rect -2966 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 586890 474854
rect -2966 474586 586890 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -2966 439174 586890 439206
rect -2966 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 586890 439174
rect -2966 438854 586890 438938
rect -2966 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 586890 438854
rect -2966 438586 586890 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -2966 403174 586890 403206
rect -2966 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 586890 403174
rect -2966 402854 586890 402938
rect -2966 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 586890 402854
rect -2966 402586 586890 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -2966 367174 586890 367206
rect -2966 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 586890 367174
rect -2966 366854 586890 366938
rect -2966 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 586890 366854
rect -2966 366586 586890 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -2966 331174 586890 331206
rect -2966 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 586890 331174
rect -2966 330854 586890 330938
rect -2966 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 586890 330854
rect -2966 330586 586890 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -2966 295174 586890 295206
rect -2966 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 586890 295174
rect -2966 294854 586890 294938
rect -2966 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 586890 294854
rect -2966 294586 586890 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -2966 259174 586890 259206
rect -2966 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 586890 259174
rect -2966 258854 586890 258938
rect -2966 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 586890 258854
rect -2966 258586 586890 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -2966 223174 586890 223206
rect -2966 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 586890 223174
rect -2966 222854 586890 222938
rect -2966 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 586890 222854
rect -2966 222586 586890 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -2966 187174 586890 187206
rect -2966 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 179610 187174
rect 179846 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 586890 187174
rect -2966 186854 586890 186938
rect -2966 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 179610 186854
rect 179846 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 586890 186854
rect -2966 186586 586890 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 164250 183454
rect 164486 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 194970 183454
rect 195206 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 164250 183134
rect 164486 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 194970 183134
rect 195206 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -2966 151174 586890 151206
rect -2966 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 586890 151174
rect -2966 150854 586890 150938
rect -2966 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 586890 150854
rect -2966 150586 586890 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -2966 115174 586890 115206
rect -2966 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 586890 115174
rect -2966 114854 586890 114938
rect -2966 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 586890 114854
rect -2966 114586 586890 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -2966 79174 586890 79206
rect -2966 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 586890 79174
rect -2966 78854 586890 78938
rect -2966 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 586890 78854
rect -2966 78586 586890 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -2966 43174 586890 43206
rect -2966 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 586890 43174
rect -2966 42854 586890 42938
rect -2966 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 586890 42854
rect -2966 42586 586890 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -2966 7174 586890 7206
rect -2966 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 586890 7174
rect -2966 6854 586890 6938
rect -2966 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 586890 6854
rect -2966 6586 586890 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
use macro_2to3  u_macro_2to3
timestamp 0
transform 1 0 280000 0 1 320000
box 1066 0 48890 50000
use macro_2xdrive  u_macro_2xdrive
timestamp 0
transform 1 0 220000 0 1 240000
box 1066 0 48890 50000
use macro_and_inv  u_macro_and_inv
timestamp 0
transform 1 0 340000 0 1 400000
box 1066 0 48890 50000
use macro_golden  u_macro_golden
timestamp 0
transform 1 0 160000 0 1 160000
box 1066 0 48890 50000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -1894 2414 705830 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -1894 38414 705830 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -1894 74414 705830 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -1894 110414 705830 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -1894 146414 705830 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -1894 182414 705830 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -1894 218414 705830 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -1894 254414 705830 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -1894 290414 705830 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -1894 326414 705830 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -1894 362414 705830 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -1894 398414 705830 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -1894 434414 705830 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -1894 470414 705830 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -1894 506414 705830 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -1894 542414 705830 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -1894 578414 705830 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2966 2866 586890 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2966 38866 586890 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2966 74866 586890 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2966 110866 586890 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2966 146866 586890 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2966 182866 586890 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2966 218866 586890 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2966 254866 586890 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2966 290866 586890 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2966 326866 586890 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2966 362866 586890 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2966 398866 586890 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2966 434866 586890 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2966 470866 586890 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2966 506866 586890 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2966 542866 586890 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2966 578866 586890 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2966 614866 586890 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2966 650866 586890 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2966 686866 586890 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 5514 -1894 6134 705830 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 41514 -1894 42134 705830 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 77514 -1894 78134 705830 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 113514 -1894 114134 705830 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 149514 -1894 150134 705830 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 185514 -1894 186134 705830 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 221514 -1894 222134 705830 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 257514 -1894 258134 705830 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 293514 -1894 294134 705830 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 329514 -1894 330134 705830 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 365514 -1894 366134 705830 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 401514 -1894 402134 705830 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 437514 -1894 438134 705830 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 473514 -1894 474134 705830 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 509514 -1894 510134 705830 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 545514 -1894 546134 705830 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 581514 -1894 582134 705830 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -2966 6586 586890 7206 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -2966 42586 586890 43206 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -2966 78586 586890 79206 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -2966 114586 586890 115206 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -2966 150586 586890 151206 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -2966 186586 586890 187206 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -2966 222586 586890 223206 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -2966 258586 586890 259206 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -2966 294586 586890 295206 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -2966 330586 586890 331206 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -2966 366586 586890 367206 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -2966 402586 586890 403206 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -2966 438586 586890 439206 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -2966 474586 586890 475206 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -2966 510586 586890 511206 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -2966 546586 586890 547206 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -2966 582586 586890 583206 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -2966 618586 586890 619206 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -2966 654586 586890 655206 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -2966 690586 586890 691206 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 533 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 534 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 535 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 536 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 537 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 538 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 539 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 540 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 541 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 542 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 543 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 544 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 545 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 546 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 547 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 548 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 549 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 550 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 551 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 552 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 553 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 554 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 555 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 556 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 557 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 558 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 559 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 560 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 561 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 562 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 563 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 564 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 565 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 566 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 567 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 568 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 569 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 570 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 571 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 572 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 573 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 574 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 575 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 576 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 577 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 578 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 579 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 580 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 581 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 582 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 583 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 584 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 585 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 586 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 587 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 588 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 589 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 590 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 591 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 592 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 593 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 594 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 595 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 596 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 597 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 598 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 599 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 600 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 601 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 602 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 603 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 604 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 605 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 606 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 607 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 608 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 609 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 610 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 611 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 612 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 613 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 614 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 615 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 616 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 617 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 618 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 619 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 620 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 621 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 622 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 623 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 624 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 625 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 626 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 627 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 628 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 629 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 630 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 631 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 632 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 633 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 634 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 635 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 636 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 637 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 638 nsew signal input
rlabel via4 195088 183336 195088 183336 0 vccd1
rlabel via4 185984 187056 185984 187056 0 vssd1
rlabel metal3 581954 6596 581954 6596 0 io_in[0]
rlabel metal2 175398 211028 175398 211028 0 io_in[10]
rlabel metal2 176357 209916 176357 209916 0 io_in[11]
rlabel metal2 237406 293148 237406 293148 0 io_in[12]
rlabel metal2 237498 293896 237498 293896 0 io_in[13]
rlabel via2 580198 670701 580198 670701 0 io_in[14]
rlabel metal2 558946 580625 558946 580625 0 io_in[15]
rlabel metal2 272458 333778 272458 333778 0 io_in[16]
rlabel metal2 213210 253198 213210 253198 0 io_in[17]
rlabel metal2 273102 333200 273102 333200 0 io_in[18]
rlabel via1 365102 449429 365102 449429 0 io_in[19]
rlabel metal3 581908 46308 581908 46308 0 io_in[1]
rlabel metal2 366314 449956 366314 449956 0 io_in[20]
rlabel metal2 273286 464032 273286 464032 0 io_in[21]
rlabel metal1 248906 295766 248906 295766 0 io_in[22]
rlabel metal2 369626 449956 369626 449956 0 io_in[23]
rlabel metal2 190801 209916 190801 209916 0 io_in[24]
rlabel metal2 191905 209916 191905 209916 0 io_in[25]
rlabel metal3 1832 579972 1832 579972 0 io_in[26]
rlabel metal3 1648 527884 1648 527884 0 io_in[27]
rlabel metal2 195125 209916 195125 209916 0 io_in[28]
rlabel metal3 1924 423572 1924 423572 0 io_in[29]
rlabel metal2 229770 332928 229770 332928 0 io_in[2]
rlabel metal3 1878 371348 1878 371348 0 io_in[30]
rlabel metal3 1878 319260 1878 319260 0 io_in[31]
rlabel metal3 1694 267172 1694 267172 0 io_in[32]
rlabel metal3 1878 214948 1878 214948 0 io_in[33]
rlabel metal3 1832 162860 1832 162860 0 io_in[34]
rlabel metal3 1740 110636 1740 110636 0 io_in[35]
rlabel metal2 383978 449956 383978 449956 0 io_in[36]
rlabel metal2 385128 449956 385128 449956 0 io_in[37]
rlabel metal3 582046 126004 582046 126004 0 io_in[3]
rlabel metal2 219282 289442 219282 289442 0 io_in[4]
rlabel metal2 173558 211752 173558 211752 0 io_in[5]
rlabel metal1 232760 295358 232760 295358 0 io_in[6]
rlabel metal2 172086 210926 172086 210926 0 io_in[7]
rlabel metal2 173045 209916 173045 209916 0 io_in[8]
rlabel metal2 174195 209916 174195 209916 0 io_in[9]
rlabel metal3 583556 32368 583556 32368 0 io_oeb[0]
rlabel metal2 175766 211198 175766 211198 0 io_oeb[10]
rlabel metal2 236854 295902 236854 295902 0 io_oeb[11]
rlabel metal2 237958 293299 237958 293299 0 io_oeb[12]
rlabel metal2 580198 643569 580198 643569 0 io_oeb[13]
rlabel metal2 580198 697085 580198 697085 0 io_oeb[14]
rlabel metal2 527206 586714 527206 586714 0 io_oeb[15]
rlabel metal2 210726 253028 210726 253028 0 io_oeb[16]
rlabel metal2 334650 413474 334650 413474 0 io_oeb[17]
rlabel metal2 364520 449956 364520 449956 0 io_oeb[18]
rlabel metal2 271354 370668 271354 370668 0 io_oeb[19]
rlabel metal3 583556 72352 583556 72352 0 io_oeb[1]
rlabel metal2 366682 449956 366682 449956 0 io_oeb[20]
rlabel metal2 367786 449956 367786 449956 0 io_oeb[21]
rlabel metal2 308154 411570 308154 411570 0 io_oeb[22]
rlabel metal2 370116 450099 370116 450099 0 io_oeb[23]
rlabel metal3 1556 658172 1556 658172 0 io_oeb[24]
rlabel metal2 192181 209916 192181 209916 0 io_oeb[25]
rlabel metal2 373428 450031 373428 450031 0 io_oeb[26]
rlabel metal3 1694 501772 1694 501772 0 io_oeb[27]
rlabel metal3 1694 449548 1694 449548 0 io_oeb[28]
rlabel metal2 256825 289884 256825 289884 0 io_oeb[29]
rlabel metal2 580198 112965 580198 112965 0 io_oeb[2]
rlabel metal3 1832 345372 1832 345372 0 io_oeb[30]
rlabel metal3 1878 293148 1878 293148 0 io_oeb[31]
rlabel metal3 1832 241060 1832 241060 0 io_oeb[32]
rlabel metal3 1740 188836 1740 188836 0 io_oeb[33]
rlabel metal3 1970 136748 1970 136748 0 io_oeb[34]
rlabel metal3 1924 84660 1924 84660 0 io_oeb[35]
rlabel metal3 1924 45492 1924 45492 0 io_oeb[36]
rlabel metal3 1878 6460 1878 6460 0 io_oeb[37]
rlabel metal2 579922 152915 579922 152915 0 io_oeb[3]
rlabel metal2 229126 292322 229126 292322 0 io_oeb[4]
rlabel metal2 230230 292118 230230 292118 0 io_oeb[5]
rlabel metal2 171297 209916 171297 209916 0 io_oeb[6]
rlabel metal2 172309 209916 172309 209916 0 io_oeb[7]
rlabel metal2 173413 209916 173413 209916 0 io_oeb[8]
rlabel metal2 174517 209916 174517 209916 0 io_oeb[9]
rlabel metal2 580106 20213 580106 20213 0 io_out[0]
rlabel metal2 176134 212320 176134 212320 0 io_out[10]
rlabel metal2 237123 289884 237123 289884 0 io_out[11]
rlabel metal2 237406 291992 237406 291992 0 io_out[12]
rlabel metal2 237498 292264 237498 292264 0 io_out[13]
rlabel metal3 581908 683876 581908 683876 0 io_out[14]
rlabel metal2 542386 583379 542386 583379 0 io_out[15]
rlabel metal2 242742 292084 242742 292084 0 io_out[16]
rlabel metal2 243747 289884 243747 289884 0 io_out[17]
rlabel metal2 364842 449956 364842 449956 0 io_out[18]
rlabel metal2 365946 449956 365946 449956 0 io_out[19]
rlabel metal3 193545 275196 193545 275196 0 io_out[1]
rlabel metal2 367202 449956 367202 449956 0 io_out[20]
rlabel metal2 368154 449956 368154 449956 0 io_out[21]
rlabel metal2 369258 449956 369258 449956 0 io_out[22]
rlabel metal2 190585 209780 190585 209780 0 io_out[23]
rlabel metal2 191445 209916 191445 209916 0 io_out[24]
rlabel metal3 1878 619140 1878 619140 0 io_out[25]
rlabel metal3 1786 566916 1786 566916 0 io_out[26]
rlabel metal2 254886 290928 254886 290928 0 io_out[27]
rlabel metal3 1924 462604 1924 462604 0 io_out[28]
rlabel metal3 1878 410516 1878 410516 0 io_out[29]
rlabel metal2 580198 100079 580198 100079 0 io_out[2]
rlabel metal3 1740 358428 1740 358428 0 io_out[30]
rlabel metal3 2200 306204 2200 306204 0 io_out[31]
rlabel metal3 1878 254116 1878 254116 0 io_out[32]
rlabel metal1 272320 291550 272320 291550 0 io_out[33]
rlabel metal3 2016 149804 2016 149804 0 io_out[34]
rlabel metal3 1924 97580 1924 97580 0 io_out[35]
rlabel metal3 1694 58548 1694 58548 0 io_out[36]
rlabel metal3 1878 19380 1878 19380 0 io_out[37]
rlabel metal3 581908 139332 581908 139332 0 io_out[3]
rlabel metal2 229494 290792 229494 290792 0 io_out[4]
rlabel metal2 230545 289884 230545 289884 0 io_out[5]
rlabel metal2 171573 209916 171573 209916 0 io_out[6]
rlabel metal2 172723 209916 172723 209916 0 io_out[7]
rlabel metal2 173926 211164 173926 211164 0 io_out[8]
rlabel metal2 174885 209916 174885 209916 0 io_out[9]
rlabel metal2 125757 340 125757 340 0 la_data_in[0]
rlabel metal2 199686 135891 199686 135891 0 la_data_in[100]
rlabel metal1 269652 154122 269652 154122 0 la_data_in[101]
rlabel metal2 487409 340 487409 340 0 la_data_in[102]
rlabel metal2 274114 127942 274114 127942 0 la_data_in[103]
rlabel metal1 274252 256734 274252 256734 0 la_data_in[104]
rlabel metal1 351210 307530 351210 307530 0 la_data_in[105]
rlabel metal2 501577 340 501577 340 0 la_data_in[106]
rlabel metal2 505402 8116 505402 8116 0 la_data_in[107]
rlabel metal2 295366 236317 295366 236317 0 la_data_in[108]
rlabel metal4 287684 274176 287684 274176 0 la_data_in[109]
rlabel metal2 161322 1928 161322 1928 0 la_data_in[10]
rlabel metal2 293986 145894 293986 145894 0 la_data_in[110]
rlabel metal1 289570 235994 289570 235994 0 la_data_in[111]
rlabel metal2 523066 1928 523066 1928 0 la_data_in[112]
rlabel metal2 526417 340 526417 340 0 la_data_in[113]
rlabel metal2 299046 237065 299046 237065 0 la_data_in[114]
rlabel metal2 268962 144432 268962 144432 0 la_data_in[115]
rlabel metal3 330556 310080 330556 310080 0 la_data_in[116]
rlabel metal1 270848 232458 270848 232458 0 la_data_in[117]
rlabel metal2 275218 148648 275218 148648 0 la_data_in[118]
rlabel metal2 390770 355997 390770 355997 0 la_data_in[119]
rlabel metal2 294998 272544 294998 272544 0 la_data_in[11]
rlabel metal2 288374 152796 288374 152796 0 la_data_in[120]
rlabel metal2 269054 138958 269054 138958 0 la_data_in[121]
rlabel metal2 558072 16560 558072 16560 0 la_data_in[122]
rlabel metal2 561890 16560 561890 16560 0 la_data_in[123]
rlabel metal2 272274 137258 272274 137258 0 la_data_in[124]
rlabel metal2 267950 141593 267950 141593 0 la_data_in[125]
rlabel metal2 271814 136204 271814 136204 0 la_data_in[126]
rlabel metal2 328992 325680 328992 325680 0 la_data_in[127]
rlabel metal1 175950 155890 175950 155890 0 la_data_in[12]
rlabel metal1 173466 155686 173466 155686 0 la_data_in[13]
rlabel metal1 175674 152966 175674 152966 0 la_data_in[14]
rlabel metal2 178841 340 178841 340 0 la_data_in[15]
rlabel metal2 237038 231075 237038 231075 0 la_data_in[16]
rlabel metal2 186162 1690 186162 1690 0 la_data_in[17]
rlabel metal2 189750 2098 189750 2098 0 la_data_in[18]
rlabel metal2 193246 1894 193246 1894 0 la_data_in[19]
rlabel metal1 232254 231438 232254 231438 0 la_data_in[1]
rlabel metal2 196834 1860 196834 1860 0 la_data_in[20]
rlabel metal1 178434 141474 178434 141474 0 la_data_in[21]
rlabel metal2 203918 2064 203918 2064 0 la_data_in[22]
rlabel metal2 207223 340 207223 340 0 la_data_in[23]
rlabel metal2 211002 2234 211002 2234 0 la_data_in[24]
rlabel metal2 214222 16560 214222 16560 0 la_data_in[25]
rlabel metal2 218086 1724 218086 1724 0 la_data_in[26]
rlabel metal2 221582 2166 221582 2166 0 la_data_in[27]
rlabel metal2 273010 320161 273010 320161 0 la_data_in[28]
rlabel metal2 228758 1690 228758 1690 0 la_data_in[29]
rlabel metal2 132756 16560 132756 16560 0 la_data_in[2]
rlabel metal2 232254 2098 232254 2098 0 la_data_in[30]
rlabel metal2 235842 2132 235842 2132 0 la_data_in[31]
rlabel metal1 217580 153170 217580 153170 0 la_data_in[32]
rlabel metal2 215970 77044 215970 77044 0 la_data_in[33]
rlabel metal2 232530 76908 232530 76908 0 la_data_in[34]
rlabel metal2 250010 2166 250010 2166 0 la_data_in[35]
rlabel metal2 253506 1860 253506 1860 0 la_data_in[36]
rlabel metal2 257094 1826 257094 1826 0 la_data_in[37]
rlabel metal2 253138 3570 253138 3570 0 la_data_in[38]
rlabel metal2 233128 229080 233128 229080 0 la_data_in[39]
rlabel metal2 136482 2030 136482 2030 0 la_data_in[3]
rlabel metal2 267766 2183 267766 2183 0 la_data_in[40]
rlabel metal2 271262 1860 271262 1860 0 la_data_in[41]
rlabel metal2 274850 1826 274850 1826 0 la_data_in[42]
rlabel metal1 274988 230418 274988 230418 0 la_data_in[43]
rlabel metal2 244168 231268 244168 231268 0 la_data_in[44]
rlabel metal2 285430 1690 285430 1690 0 la_data_in[45]
rlabel metal2 289018 2166 289018 2166 0 la_data_in[46]
rlabel metal1 273102 229874 273102 229874 0 la_data_in[47]
rlabel metal2 271814 156978 271814 156978 0 la_data_in[48]
rlabel metal2 296010 77350 296010 77350 0 la_data_in[49]
rlabel metal2 139833 340 139833 340 0 la_data_in[4]
rlabel metal2 303186 2200 303186 2200 0 la_data_in[50]
rlabel metal2 306774 2234 306774 2234 0 la_data_in[51]
rlabel metal2 269330 229772 269330 229772 0 la_data_in[52]
rlabel metal2 313858 1792 313858 1792 0 la_data_in[53]
rlabel metal2 275402 139094 275402 139094 0 la_data_in[54]
rlabel metal2 307510 308040 307510 308040 0 la_data_in[55]
rlabel metal2 307510 309060 307510 309060 0 la_data_in[56]
rlabel metal2 270066 232288 270066 232288 0 la_data_in[57]
rlabel metal1 276552 231778 276552 231778 0 la_data_in[58]
rlabel metal2 335110 1860 335110 1860 0 la_data_in[59]
rlabel metal1 278346 372062 278346 372062 0 la_data_in[5]
rlabel metal2 308292 306360 308292 306360 0 la_data_in[60]
rlabel metal2 308982 307581 308982 307581 0 la_data_in[61]
rlabel metal2 345545 340 345545 340 0 la_data_in[62]
rlabel metal2 349278 1163 349278 1163 0 la_data_in[63]
rlabel metal2 249642 136238 249642 136238 0 la_data_in[64]
rlabel metal2 309810 308703 309810 308703 0 la_data_in[65]
rlabel metal2 251114 125222 251114 125222 0 la_data_in[66]
rlabel metal1 270480 233206 270480 233206 0 la_data_in[67]
rlabel metal2 367034 2234 367034 2234 0 la_data_in[68]
rlabel metal2 251022 134912 251022 134912 0 la_data_in[69]
rlabel metal1 173558 152354 173558 152354 0 la_data_in[6]
rlabel metal1 252264 3162 252264 3162 0 la_data_in[70]
rlabel metal3 311190 303620 311190 303620 0 la_data_in[71]
rlabel metal1 270710 232356 270710 232356 0 la_data_in[72]
rlabel metal2 384790 2132 384790 2132 0 la_data_in[73]
rlabel metal2 388049 340 388049 340 0 la_data_in[74]
rlabel metal2 391874 1860 391874 1860 0 la_data_in[75]
rlabel metal2 252494 123828 252494 123828 0 la_data_in[76]
rlabel metal2 276046 232628 276046 232628 0 la_data_in[77]
rlabel metal1 272274 222802 272274 222802 0 la_data_in[78]
rlabel metal2 313306 311440 313306 311440 0 la_data_in[79]
rlabel metal2 150558 16560 150558 16560 0 la_data_in[7]
rlabel metal2 409393 340 409393 340 0 la_data_in[80]
rlabel metal2 412889 340 412889 340 0 la_data_in[81]
rlabel metal2 289754 231098 289754 231098 0 la_data_in[82]
rlabel metal2 285798 137598 285798 137598 0 la_data_in[83]
rlabel metal2 423798 1690 423798 1690 0 la_data_in[84]
rlabel metal2 427057 340 427057 340 0 la_data_in[85]
rlabel metal1 288788 237422 288788 237422 0 la_data_in[86]
rlabel metal2 434233 340 434233 340 0 la_data_in[87]
rlabel metal2 290950 144194 290950 144194 0 la_data_in[88]
rlabel metal2 262154 136272 262154 136272 0 la_data_in[89]
rlabel metal2 154001 340 154001 340 0 la_data_in[8]
rlabel metal2 256082 127942 256082 127942 0 la_data_in[90]
rlabel metal2 448638 59167 448638 59167 0 la_data_in[91]
rlabel metal2 291778 227086 291778 227086 0 la_data_in[92]
rlabel metal2 291962 133484 291962 133484 0 la_data_in[93]
rlabel metal2 289754 126548 289754 126548 0 la_data_in[94]
rlabel metal2 462569 340 462569 340 0 la_data_in[95]
rlabel metal2 466065 340 466065 340 0 la_data_in[96]
rlabel metal2 469890 1928 469890 1928 0 la_data_in[97]
rlabel metal2 473478 1928 473478 1928 0 la_data_in[98]
rlabel metal2 275402 125222 275402 125222 0 la_data_in[99]
rlabel metal1 214774 236198 214774 236198 0 la_data_in[9]
rlabel metal3 172017 153068 172017 153068 0 la_data_out[0]
rlabel metal4 329268 328114 329268 328114 0 la_data_out[100]
rlabel metal2 485017 340 485017 340 0 la_data_out[101]
rlabel metal2 488704 16560 488704 16560 0 la_data_out[102]
rlabel metal2 346058 348398 346058 348398 0 la_data_out[103]
rlabel metal2 380926 326723 380926 326723 0 la_data_out[104]
rlabel metal2 392242 355436 392242 355436 0 la_data_out[105]
rlabel metal2 502688 16560 502688 16560 0 la_data_out[106]
rlabel metal2 506506 161660 506506 161660 0 la_data_out[107]
rlabel metal3 322092 309060 322092 309060 0 la_data_out[108]
rlabel metal2 208242 160820 208242 160820 0 la_data_out[109]
rlabel metal2 174754 137659 174754 137659 0 la_data_out[10]
rlabel metal2 237038 191148 237038 191148 0 la_data_out[110]
rlabel metal2 520766 2064 520766 2064 0 la_data_out[111]
rlabel metal2 524025 340 524025 340 0 la_data_out[112]
rlabel metal1 273976 232186 273976 232186 0 la_data_out[113]
rlabel metal2 322966 273887 322966 273887 0 la_data_out[114]
rlabel metal1 384146 349078 384146 349078 0 la_data_out[115]
rlabel metal2 538331 340 538331 340 0 la_data_out[116]
rlabel metal2 392334 357068 392334 357068 0 la_data_out[117]
rlabel metal2 545514 1758 545514 1758 0 la_data_out[118]
rlabel metal2 330326 323340 330326 323340 0 la_data_out[119]
rlabel metal3 174593 149124 174593 149124 0 la_data_out[11]
rlabel metal1 385480 333982 385480 333982 0 la_data_out[120]
rlabel metal2 205666 159929 205666 159929 0 la_data_out[121]
rlabel metal2 559537 340 559537 340 0 la_data_out[122]
rlabel metal2 563171 340 563171 340 0 la_data_out[123]
rlabel metal2 326922 303144 326922 303144 0 la_data_out[124]
rlabel metal1 326646 291142 326646 291142 0 la_data_out[125]
rlabel metal2 387090 162605 387090 162605 0 la_data_out[126]
rlabel metal2 577438 1860 577438 1860 0 la_data_out[127]
rlabel metal2 174616 151800 174616 151800 0 la_data_out[12]
rlabel metal2 172953 340 172953 340 0 la_data_out[13]
rlabel metal1 176364 28934 176364 28934 0 la_data_out[14]
rlabel metal2 180274 1911 180274 1911 0 la_data_out[15]
rlabel metal1 293434 305898 293434 305898 0 la_data_out[16]
rlabel metal2 187121 340 187121 340 0 la_data_out[17]
rlabel metal2 190854 1724 190854 1724 0 la_data_out[18]
rlabel metal2 194442 2132 194442 2132 0 la_data_out[19]
rlabel metal1 291778 305286 291778 305286 0 la_data_out[1]
rlabel metal2 197662 16560 197662 16560 0 la_data_out[20]
rlabel metal1 294906 305728 294906 305728 0 la_data_out[21]
rlabel metal2 296194 263330 296194 263330 0 la_data_out[22]
rlabel metal1 298816 307734 298816 307734 0 la_data_out[23]
rlabel metal2 211961 340 211961 340 0 la_data_out[24]
rlabel metal2 215503 340 215503 340 0 la_data_out[25]
rlabel metal2 218730 16560 218730 16560 0 la_data_out[26]
rlabel metal2 222502 16560 222502 16560 0 la_data_out[27]
rlabel metal2 294722 268056 294722 268056 0 la_data_out[28]
rlabel metal2 229625 340 229625 340 0 la_data_out[29]
rlabel metal2 134037 340 134037 340 0 la_data_out[2]
rlabel metal2 233358 16560 233358 16560 0 la_data_out[30]
rlabel metal2 236801 340 236801 340 0 la_data_out[31]
rlabel metal2 351394 351220 351394 351220 0 la_data_out[32]
rlabel metal2 347438 349350 347438 349350 0 la_data_out[33]
rlabel metal2 288098 263874 288098 263874 0 la_data_out[34]
rlabel metal2 251206 1792 251206 1792 0 la_data_out[35]
rlabel metal2 254702 1996 254702 1996 0 la_data_out[36]
rlabel metal2 253414 3876 253414 3876 0 la_data_out[37]
rlabel metal2 289294 268464 289294 268464 0 la_data_out[38]
rlabel metal1 275356 231778 275356 231778 0 la_data_out[39]
rlabel metal2 137441 340 137441 340 0 la_data_out[3]
rlabel metal1 253230 3978 253230 3978 0 la_data_out[40]
rlabel metal2 272458 2098 272458 2098 0 la_data_out[41]
rlabel metal2 276046 71247 276046 71247 0 la_data_out[42]
rlabel metal2 279305 340 279305 340 0 la_data_out[43]
rlabel metal3 283222 236028 283222 236028 0 la_data_out[44]
rlabel metal2 286626 2064 286626 2064 0 la_data_out[45]
rlabel metal2 290214 1724 290214 1724 0 la_data_out[46]
rlabel metal2 293710 1622 293710 1622 0 la_data_out[47]
rlabel metal1 301668 295426 301668 295426 0 la_data_out[48]
rlabel metal2 300794 1962 300794 1962 0 la_data_out[49]
rlabel metal2 270434 308788 270434 308788 0 la_data_out[4]
rlabel metal2 304145 340 304145 340 0 la_data_out[50]
rlabel metal2 307970 1911 307970 1911 0 la_data_out[51]
rlabel metal2 311466 2030 311466 2030 0 la_data_out[52]
rlabel metal2 315054 1860 315054 1860 0 la_data_out[53]
rlabel metal1 307418 300526 307418 300526 0 la_data_out[54]
rlabel metal2 307050 115056 307050 115056 0 la_data_out[55]
rlabel metal1 306820 223006 306820 223006 0 la_data_out[56]
rlabel metal2 329222 2098 329222 2098 0 la_data_out[57]
rlabel metal2 332672 16560 332672 16560 0 la_data_out[58]
rlabel metal1 249412 218042 249412 218042 0 la_data_out[59]
rlabel metal1 269698 318410 269698 318410 0 la_data_out[5]
rlabel metal1 248998 222122 248998 222122 0 la_data_out[60]
rlabel metal2 343153 340 343153 340 0 la_data_out[61]
rlabel metal2 346978 2132 346978 2132 0 la_data_out[62]
rlabel metal2 350474 1860 350474 1860 0 la_data_out[63]
rlabel metal2 354062 2047 354062 2047 0 la_data_out[64]
rlabel metal2 211830 198220 211830 198220 0 la_data_out[65]
rlabel metal1 271078 230452 271078 230452 0 la_data_out[66]
rlabel metal1 311006 310930 311006 310930 0 la_data_out[67]
rlabel metal1 328578 4046 328578 4046 0 la_data_out[68]
rlabel metal2 371489 340 371489 340 0 la_data_out[69]
rlabel metal4 174800 151800 174800 151800 0 la_data_out[6]
rlabel metal1 311558 262174 311558 262174 0 la_data_out[70]
rlabel metal1 309396 292094 309396 292094 0 la_data_out[71]
rlabel metal1 312938 301886 312938 301886 0 la_data_out[72]
rlabel metal2 252126 188811 252126 188811 0 la_data_out[73]
rlabel metal1 313030 256734 313030 256734 0 la_data_out[74]
rlabel metal1 312846 311814 312846 311814 0 la_data_out[75]
rlabel metal1 253092 222054 253092 222054 0 la_data_out[76]
rlabel metal1 328578 309502 328578 309502 0 la_data_out[77]
rlabel metal1 253092 214574 253092 214574 0 la_data_out[78]
rlabel metal2 407238 1775 407238 1775 0 la_data_out[79]
rlabel metal2 151846 74722 151846 74722 0 la_data_out[7]
rlabel metal2 254886 192134 254886 192134 0 la_data_out[80]
rlabel metal2 254610 183235 254610 183235 0 la_data_out[81]
rlabel metal3 250815 222156 250815 222156 0 la_data_out[82]
rlabel metal1 254426 221374 254426 221374 0 la_data_out[83]
rlabel metal2 424994 1860 424994 1860 0 la_data_out[84]
rlabel metal3 256243 222020 256243 222020 0 la_data_out[85]
rlabel metal2 429870 160412 429870 160412 0 la_data_out[86]
rlabel metal2 255990 184280 255990 184280 0 la_data_out[87]
rlabel metal2 256174 192134 256174 192134 0 la_data_out[88]
rlabel metal2 442152 16560 442152 16560 0 la_data_out[89]
rlabel metal2 155020 16560 155020 16560 0 la_data_out[8]
rlabel metal2 446009 340 446009 340 0 la_data_out[90]
rlabel metal2 449834 1418 449834 1418 0 la_data_out[91]
rlabel metal2 257370 184586 257370 184586 0 la_data_out[92]
rlabel metal2 257462 192287 257462 192287 0 la_data_out[93]
rlabel metal1 294124 257346 294124 257346 0 la_data_out[94]
rlabel metal2 463864 16560 463864 16560 0 la_data_out[95]
rlabel metal2 466992 16560 466992 16560 0 la_data_out[96]
rlabel metal1 319976 251158 319976 251158 0 la_data_out[97]
rlabel metal1 319884 253062 319884 253062 0 la_data_out[98]
rlabel metal3 393300 313888 393300 313888 0 la_data_out[99]
rlabel metal2 270434 315622 270434 315622 0 la_data_out[9]
rlabel metal2 268686 354909 268686 354909 0 la_oenb[0]
rlabel metal2 482862 1843 482862 1843 0 la_oenb[100]
rlabel metal2 486128 16560 486128 16560 0 la_oenb[101]
rlabel metal2 489210 56916 489210 56916 0 la_oenb[102]
rlabel metal2 493297 340 493297 340 0 la_oenb[103]
rlabel metal3 231288 143820 231288 143820 0 la_oenb[104]
rlabel metal2 500112 16560 500112 16560 0 la_oenb[105]
rlabel metal2 503969 340 503969 340 0 la_oenb[106]
rlabel metal2 330418 310284 330418 310284 0 la_oenb[107]
rlabel metal2 329038 311236 329038 311236 0 la_oenb[108]
rlabel metal3 358777 102748 358777 102748 0 la_oenb[109]
rlabel metal2 293986 300339 293986 300339 0 la_oenb[10]
rlabel metal2 518137 340 518137 340 0 la_oenb[110]
rlabel metal2 521870 1928 521870 1928 0 la_oenb[111]
rlabel metal2 524952 16560 524952 16560 0 la_oenb[112]
rlabel metal2 528809 340 528809 340 0 la_oenb[113]
rlabel metal3 234255 179996 234255 179996 0 la_oenb[114]
rlabel metal1 369748 94486 369748 94486 0 la_oenb[115]
rlabel metal2 539626 60527 539626 60527 0 la_oenb[116]
rlabel metal2 542977 340 542977 340 0 la_oenb[117]
rlabel metal2 546710 3968 546710 3968 0 la_oenb[118]
rlabel metal3 235589 177276 235589 177276 0 la_oenb[119]
rlabel metal2 175490 153204 175490 153204 0 la_oenb[11]
rlabel metal3 295320 255884 295320 255884 0 la_oenb[120]
rlabel metal2 557145 340 557145 340 0 la_oenb[121]
rlabel metal2 560641 340 560641 340 0 la_oenb[122]
rlabel metal3 326232 307564 326232 307564 0 la_oenb[123]
rlabel via3 206563 159868 206563 159868 0 la_oenb[124]
rlabel via3 206885 159868 206885 159868 0 la_oenb[125]
rlabel metal2 207138 159113 207138 159113 0 la_oenb[126]
rlabel metal2 578450 16560 578450 16560 0 la_oenb[127]
rlabel via3 176203 153068 176203 153068 0 la_oenb[12]
rlabel metal2 174103 340 174103 340 0 la_oenb[13]
rlabel metal2 177882 2948 177882 2948 0 la_oenb[14]
rlabel metal1 175996 153102 175996 153102 0 la_oenb[15]
rlabel metal2 348726 339830 348726 339830 0 la_oenb[16]
rlabel metal2 188140 16560 188140 16560 0 la_oenb[17]
rlabel metal2 192050 1928 192050 1928 0 la_oenb[18]
rlabel metal2 195638 1928 195638 1928 0 la_oenb[19]
rlabel metal2 172960 151800 172960 151800 0 la_oenb[1]
rlabel metal3 177560 140828 177560 140828 0 la_oenb[20]
rlabel metal1 178664 141542 178664 141542 0 la_oenb[21]
rlabel metal1 201158 141610 201158 141610 0 la_oenb[22]
rlabel metal2 209806 3627 209806 3627 0 la_oenb[23]
rlabel metal2 213394 1911 213394 1911 0 la_oenb[24]
rlabel metal2 238694 293420 238694 293420 0 la_oenb[25]
rlabel metal2 238096 229080 238096 229080 0 la_oenb[26]
rlabel metal2 223783 340 223783 340 0 la_oenb[27]
rlabel metal2 269698 350472 269698 350472 0 la_oenb[28]
rlabel metal2 230782 16560 230782 16560 0 la_oenb[29]
rlabel metal2 135286 1911 135286 1911 0 la_oenb[2]
rlabel metal2 234646 3627 234646 3627 0 la_oenb[30]
rlabel metal2 237905 340 237905 340 0 la_oenb[31]
rlabel metal1 211738 134606 211738 134606 0 la_oenb[32]
rlabel metal3 212727 122196 212727 122196 0 la_oenb[33]
rlabel metal2 248814 1622 248814 1622 0 la_oenb[34]
rlabel metal2 252402 1911 252402 1911 0 la_oenb[35]
rlabel metal2 268778 315520 268778 315520 0 la_oenb[36]
rlabel metal2 292422 262871 292422 262871 0 la_oenb[37]
rlabel metal2 262745 340 262745 340 0 la_oenb[38]
rlabel metal3 210956 141780 210956 141780 0 la_oenb[39]
rlabel metal1 233036 233750 233036 233750 0 la_oenb[3]
rlabel metal2 270066 1911 270066 1911 0 la_oenb[40]
rlabel metal2 273463 340 273463 340 0 la_oenb[41]
rlabel metal2 276913 340 276913 340 0 la_oenb[42]
rlabel metal2 208518 234073 208518 234073 0 la_oenb[43]
rlabel metal2 211646 265693 211646 265693 0 la_oenb[44]
rlabel metal2 287585 340 287585 340 0 la_oenb[45]
rlabel metal2 291410 2030 291410 2030 0 la_oenb[46]
rlabel metal2 294906 1962 294906 1962 0 la_oenb[47]
rlabel metal2 298303 340 298303 340 0 la_oenb[48]
rlabel metal2 301990 3203 301990 3203 0 la_oenb[49]
rlabel metal4 292652 268880 292652 268880 0 la_oenb[4]
rlabel metal2 289570 258400 289570 258400 0 la_oenb[50]
rlabel metal2 309074 1962 309074 1962 0 la_oenb[51]
rlabel metal1 212198 233886 212198 233886 0 la_oenb[52]
rlabel metal2 315330 52105 315330 52105 0 la_oenb[53]
rlabel metal2 236762 180948 236762 180948 0 la_oenb[54]
rlabel metal2 323143 340 323143 340 0 la_oenb[55]
rlabel metal2 326593 340 326593 340 0 la_oenb[56]
rlabel metal2 330418 3611 330418 3611 0 la_oenb[57]
rlabel metal2 214774 234328 214774 234328 0 la_oenb[58]
rlabel metal2 337502 3475 337502 3475 0 la_oenb[59]
rlabel metal2 145721 340 145721 340 0 la_oenb[5]
rlabel metal2 308522 275629 308522 275629 0 la_oenb[60]
rlabel metal1 309718 297942 309718 297942 0 la_oenb[61]
rlabel metal2 347944 16560 347944 16560 0 la_oenb[62]
rlabel metal2 351670 2047 351670 2047 0 la_oenb[63]
rlabel metal1 248216 219266 248216 219266 0 la_oenb[64]
rlabel metal3 209967 138788 209967 138788 0 la_oenb[65]
rlabel metal4 250332 219028 250332 219028 0 la_oenb[66]
rlabel metal3 191429 209508 191429 209508 0 la_oenb[67]
rlabel metal2 219282 248400 219282 248400 0 la_oenb[68]
rlabel metal2 372784 16560 372784 16560 0 la_oenb[69]
rlabel metal2 149546 1860 149546 1860 0 la_oenb[6]
rlabel metal4 310684 295196 310684 295196 0 la_oenb[70]
rlabel metal3 207897 138516 207897 138516 0 la_oenb[71]
rlabel metal2 383594 3322 383594 3322 0 la_oenb[72]
rlabel metal2 387182 3288 387182 3288 0 la_oenb[73]
rlabel metal3 253299 218076 253299 218076 0 la_oenb[74]
rlabel metal4 312616 325680 312616 325680 0 la_oenb[75]
rlabel metal3 311144 299268 311144 299268 0 la_oenb[76]
rlabel metal4 193752 171120 193752 171120 0 la_oenb[77]
rlabel metal2 253414 116926 253414 116926 0 la_oenb[78]
rlabel metal2 408434 1860 408434 1860 0 la_oenb[79]
rlabel metal2 152490 16560 152490 16560 0 la_oenb[7]
rlabel metal4 194120 171120 194120 171120 0 la_oenb[80]
rlabel metal2 313306 303501 313306 303501 0 la_oenb[81]
rlabel metal3 195707 209508 195707 209508 0 la_oenb[82]
rlabel metal2 422602 4716 422602 4716 0 la_oenb[83]
rlabel metal2 425953 340 425953 340 0 la_oenb[84]
rlabel metal2 429449 340 429449 340 0 la_oenb[85]
rlabel metal3 196673 144364 196673 144364 0 la_oenb[86]
rlabel metal2 436770 1639 436770 1639 0 la_oenb[87]
rlabel metal4 196880 171120 196880 171120 0 la_oenb[88]
rlabel metal2 196972 219420 196972 219420 0 la_oenb[89]
rlabel metal2 156393 340 156393 340 0 la_oenb[8]
rlabel metal2 257646 173655 257646 173655 0 la_oenb[90]
rlabel metal2 257554 168895 257554 168895 0 la_oenb[91]
rlabel metal3 198122 139332 198122 139332 0 la_oenb[92]
rlabel metal2 458114 1979 458114 1979 0 la_oenb[93]
rlabel metal2 461288 16560 461288 16560 0 la_oenb[94]
rlabel metal2 465198 1911 465198 1911 0 la_oenb[95]
rlabel metal2 468503 340 468503 340 0 la_oenb[96]
rlabel metal2 472282 1894 472282 1894 0 la_oenb[97]
rlabel metal2 475778 3254 475778 3254 0 la_oenb[98]
rlabel metal1 260544 175202 260544 175202 0 la_oenb[99]
rlabel metal2 160126 1792 160126 1792 0 la_oenb[9]
rlabel metal2 1702 1928 1702 1928 0 wb_rst_i
rlabel metal2 2898 1962 2898 1962 0 wbs_ack_o
rlabel metal2 7314 16560 7314 16560 0 wbs_adr_i[0]
rlabel metal2 155618 194582 155618 194582 0 wbs_adr_i[10]
rlabel metal2 156998 192525 156998 192525 0 wbs_adr_i[11]
rlabel metal2 155802 194684 155802 194684 0 wbs_adr_i[12]
rlabel metal2 58236 16560 58236 16560 0 wbs_adr_i[13]
rlabel metal2 61863 340 61863 340 0 wbs_adr_i[14]
rlabel metal2 271446 358292 271446 358292 0 wbs_adr_i[15]
rlabel metal2 69138 1962 69138 1962 0 wbs_adr_i[16]
rlabel metal3 156722 156604 156722 156604 0 wbs_adr_i[17]
rlabel metal2 76077 340 76077 340 0 wbs_adr_i[18]
rlabel metal2 79481 340 79481 340 0 wbs_adr_i[19]
rlabel metal2 272826 321232 272826 321232 0 wbs_adr_i[1]
rlabel metal2 83076 16560 83076 16560 0 wbs_adr_i[20]
rlabel metal1 289064 299438 289064 299438 0 wbs_adr_i[21]
rlabel metal3 152766 159596 152766 159596 0 wbs_adr_i[22]
rlabel metal2 93978 1826 93978 1826 0 wbs_adr_i[23]
rlabel metal2 97060 16560 97060 16560 0 wbs_adr_i[24]
rlabel metal2 100917 340 100917 340 0 wbs_adr_i[25]
rlabel metal2 153134 194157 153134 194157 0 wbs_adr_i[26]
rlabel metal2 287730 269960 287730 269960 0 wbs_adr_i[27]
rlabel metal2 111642 1860 111642 1860 0 wbs_adr_i[28]
rlabel metal2 115230 1792 115230 1792 0 wbs_adr_i[29]
rlabel metal2 17066 1928 17066 1928 0 wbs_adr_i[2]
rlabel metal2 118818 1996 118818 1996 0 wbs_adr_i[30]
rlabel metal2 122314 1911 122314 1911 0 wbs_adr_i[31]
rlabel metal2 21298 16560 21298 16560 0 wbs_adr_i[3]
rlabel metal2 26397 340 26397 340 0 wbs_adr_i[4]
rlabel metal2 155342 157604 155342 157604 0 wbs_adr_i[5]
rlabel metal2 154514 199376 154514 199376 0 wbs_adr_i[6]
rlabel metal2 37214 1996 37214 1996 0 wbs_adr_i[7]
rlabel metal2 40473 340 40473 340 0 wbs_adr_i[8]
rlabel metal2 44298 3627 44298 3627 0 wbs_adr_i[9]
rlabel metal2 4094 1826 4094 1826 0 wbs_cyc_i
rlabel metal2 268594 319804 268594 319804 0 wbs_dat_i[0]
rlabel metal2 156722 194463 156722 194463 0 wbs_dat_i[10]
rlabel metal2 210910 274312 210910 274312 0 wbs_dat_i[11]
rlabel metal2 55660 16560 55660 16560 0 wbs_dat_i[12]
rlabel metal2 59517 340 59517 340 0 wbs_dat_i[13]
rlabel metal2 62698 16560 62698 16560 0 wbs_dat_i[14]
rlabel metal1 287960 294338 287960 294338 0 wbs_dat_i[15]
rlabel metal2 70097 340 70097 340 0 wbs_dat_i[16]
rlabel metal1 167486 139434 167486 139434 0 wbs_dat_i[17]
rlabel metal2 77418 1996 77418 1996 0 wbs_dat_i[18]
rlabel metal2 80914 1911 80914 1911 0 wbs_dat_i[19]
rlabel metal2 17250 72046 17250 72046 0 wbs_dat_i[1]
rlabel metal2 199042 231506 199042 231506 0 wbs_dat_i[20]
rlabel metal1 289202 298078 289202 298078 0 wbs_dat_i[21]
rlabel metal1 129766 134606 129766 134606 0 wbs_dat_i[22]
rlabel metal2 94937 340 94937 340 0 wbs_dat_i[23]
rlabel metal2 98433 340 98433 340 0 wbs_dat_i[24]
rlabel metal2 102212 16560 102212 16560 0 wbs_dat_i[25]
rlabel metal4 290628 258544 290628 258544 0 wbs_dat_i[26]
rlabel metal2 109342 1996 109342 1996 0 wbs_dat_i[27]
rlabel metal1 171350 156638 171350 156638 0 wbs_dat_i[28]
rlabel metal2 116196 16560 116196 16560 0 wbs_dat_i[29]
rlabel metal2 18262 1622 18262 1622 0 wbs_dat_i[2]
rlabel metal2 119922 1860 119922 1860 0 wbs_dat_i[30]
rlabel metal2 133170 76092 133170 76092 0 wbs_dat_i[31]
rlabel metal2 23046 1928 23046 1928 0 wbs_dat_i[3]
rlabel metal2 27738 1792 27738 1792 0 wbs_dat_i[4]
rlabel metal2 36570 66793 36570 66793 0 wbs_dat_i[5]
rlabel metal2 34677 340 34677 340 0 wbs_dat_i[6]
rlabel metal2 38410 1928 38410 1928 0 wbs_dat_i[7]
rlabel metal2 41906 1928 41906 1928 0 wbs_dat_i[8]
rlabel metal2 45257 340 45257 340 0 wbs_dat_i[9]
rlabel metal2 153042 200481 153042 200481 0 wbs_dat_o[0]
rlabel metal3 255484 294644 255484 294644 0 wbs_dat_o[10]
rlabel metal2 53537 340 53537 340 0 wbs_dat_o[11]
rlabel metal2 57033 340 57033 340 0 wbs_dat_o[12]
rlabel metal2 60858 60544 60858 60544 0 wbs_dat_o[13]
rlabel metal2 64354 2574 64354 2574 0 wbs_dat_o[14]
rlabel metal2 288006 296463 288006 296463 0 wbs_dat_o[15]
rlabel metal2 288282 299183 288282 299183 0 wbs_dat_o[16]
rlabel metal2 74796 16560 74796 16560 0 wbs_dat_o[17]
rlabel metal2 78614 1860 78614 1860 0 wbs_dat_o[18]
rlabel metal2 81873 340 81873 340 0 wbs_dat_o[19]
rlabel metal2 14529 340 14529 340 0 wbs_dat_o[1]
rlabel metal1 289248 301614 289248 301614 0 wbs_dat_o[20]
rlabel metal2 212106 272884 212106 272884 0 wbs_dat_o[21]
rlabel metal2 230092 229080 230092 229080 0 wbs_dat_o[22]
rlabel metal2 96041 340 96041 340 0 wbs_dat_o[23]
rlabel metal2 99636 16560 99636 16560 0 wbs_dat_o[24]
rlabel metal2 103362 4648 103362 4648 0 wbs_dat_o[25]
rlabel metal2 106713 340 106713 340 0 wbs_dat_o[26]
rlabel metal3 268870 257380 268870 257380 0 wbs_dat_o[27]
rlabel metal2 114034 1860 114034 1860 0 wbs_dat_o[28]
rlabel metal2 117477 340 117477 340 0 wbs_dat_o[29]
rlabel metal2 19412 16560 19412 16560 0 wbs_dat_o[2]
rlabel metal2 121118 1996 121118 1996 0 wbs_dat_o[30]
rlabel metal2 124706 1996 124706 1996 0 wbs_dat_o[31]
rlabel metal2 24242 1826 24242 1826 0 wbs_dat_o[3]
rlabel metal2 153962 127806 153962 127806 0 wbs_dat_o[4]
rlabel metal2 32193 340 32193 340 0 wbs_dat_o[5]
rlabel metal2 35972 16560 35972 16560 0 wbs_dat_o[6]
rlabel metal2 39369 340 39369 340 0 wbs_dat_o[7]
rlabel metal2 42957 340 42957 340 0 wbs_dat_o[8]
rlabel metal1 158102 3468 158102 3468 0 wbs_dat_o[9]
rlabel metal1 252448 309978 252448 309978 0 wbs_sel_i[0]
rlabel metal2 15962 1911 15962 1911 0 wbs_sel_i[1]
rlabel metal2 20417 340 20417 340 0 wbs_sel_i[2]
rlabel metal2 25346 6722 25346 6722 0 wbs_sel_i[3]
rlabel metal2 5290 2574 5290 2574 0 wbs_stb_i
rlabel metal2 6486 1894 6486 1894 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
