magic
tech sky130A
magscale 1 2
timestamp 1666199351
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 1 21 911 203
rect 30 -17 64 21
<< locali >>
rect 467 333 533 425
rect 635 333 701 493
rect 835 333 903 493
rect 467 299 903 333
rect 18 211 248 265
rect 282 211 444 265
rect 478 211 641 265
rect 735 119 801 299
rect 835 151 903 265
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 18 333 89 493
rect 123 367 157 527
rect 191 333 257 493
rect 291 459 601 493
rect 291 367 325 459
rect 359 333 425 425
rect 18 299 425 333
rect 567 367 601 459
rect 735 367 801 527
rect 18 143 701 177
rect 18 51 89 143
rect 123 17 157 109
rect 191 51 257 143
rect 291 17 393 109
rect 435 51 501 143
rect 535 17 601 109
rect 635 85 701 143
rect 835 85 903 117
rect 635 51 903 85
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
rlabel locali s 18 211 248 265 6 A1
port 1 nsew signal input
rlabel locali s 282 211 444 265 6 A2
port 2 nsew signal input
rlabel locali s 478 211 641 265 6 A3
port 3 nsew signal input
rlabel locali s 835 151 903 265 6 B1
port 4 nsew signal input
rlabel metal1 s 0 -48 920 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 21 911 203 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 958 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 920 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 735 119 801 299 6 Y
port 9 nsew signal output
rlabel locali s 467 299 903 333 6 Y
port 9 nsew signal output
rlabel locali s 835 333 903 493 6 Y
port 9 nsew signal output
rlabel locali s 635 333 701 493 6 Y
port 9 nsew signal output
rlabel locali s 467 333 533 425 6 Y
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 920 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1439140
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1430212
<< end >>
