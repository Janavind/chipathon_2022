magic
tech sky130B
magscale 1 2
timestamp 1666199351
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 361 163 642 203
rect 1 27 642 163
rect 29 -17 63 27
rect 361 21 642 27
<< scnmos >>
rect 79 53 109 137
rect 258 53 288 137
rect 342 53 372 137
rect 440 47 470 177
rect 524 47 554 177
<< scpmoshvt >>
rect 79 297 109 381
rect 270 297 300 381
rect 342 297 372 381
rect 440 297 470 497
rect 524 297 554 497
<< ndiff >>
rect 387 137 440 177
rect 27 106 79 137
rect 27 72 35 106
rect 69 72 79 106
rect 27 53 79 72
rect 109 97 258 137
rect 109 63 119 97
rect 153 63 214 97
rect 248 63 258 97
rect 109 53 258 63
rect 288 111 342 137
rect 288 77 298 111
rect 332 77 342 111
rect 288 53 342 77
rect 372 97 440 137
rect 372 63 392 97
rect 426 63 440 97
rect 372 53 440 63
rect 387 47 440 53
rect 470 135 524 177
rect 470 101 480 135
rect 514 101 524 135
rect 470 47 524 101
rect 554 162 616 177
rect 554 128 564 162
rect 598 128 616 162
rect 554 94 616 128
rect 554 60 564 94
rect 598 60 616 94
rect 554 47 616 60
<< pdiff >>
rect 387 485 440 497
rect 387 451 395 485
rect 429 451 440 485
rect 387 417 440 451
rect 387 383 395 417
rect 429 383 440 417
rect 387 381 440 383
rect 27 349 79 381
rect 27 315 35 349
rect 69 315 79 349
rect 27 297 79 315
rect 109 343 161 381
rect 109 309 119 343
rect 153 309 161 343
rect 109 297 161 309
rect 218 354 270 381
rect 218 320 226 354
rect 260 320 270 354
rect 218 297 270 320
rect 300 297 342 381
rect 372 297 440 381
rect 470 454 524 497
rect 470 420 480 454
rect 514 420 524 454
rect 470 386 524 420
rect 470 352 480 386
rect 514 352 524 386
rect 470 297 524 352
rect 554 483 616 497
rect 554 449 564 483
rect 598 449 616 483
rect 554 415 616 449
rect 554 381 564 415
rect 598 381 616 415
rect 554 347 616 381
rect 554 313 564 347
rect 598 313 616 347
rect 554 297 616 313
<< ndiffc >>
rect 35 72 69 106
rect 119 63 153 97
rect 214 63 248 97
rect 298 77 332 111
rect 392 63 426 97
rect 480 101 514 135
rect 564 128 598 162
rect 564 60 598 94
<< pdiffc >>
rect 395 451 429 485
rect 395 383 429 417
rect 35 315 69 349
rect 119 309 153 343
rect 226 320 260 354
rect 480 420 514 454
rect 480 352 514 386
rect 564 449 598 483
rect 564 381 598 415
rect 564 313 598 347
<< poly >>
rect 440 497 470 523
rect 524 497 554 523
rect 168 473 372 483
rect 168 439 184 473
rect 218 453 372 473
rect 218 439 234 453
rect 168 429 234 439
rect 79 381 109 407
rect 270 381 300 407
rect 342 381 372 453
rect 79 265 109 297
rect 270 265 300 297
rect 21 249 109 265
rect 21 215 35 249
rect 69 215 109 249
rect 21 199 109 215
rect 216 249 300 265
rect 216 215 226 249
rect 260 215 300 249
rect 216 199 300 215
rect 79 137 109 199
rect 258 137 288 199
rect 342 137 372 297
rect 440 265 470 297
rect 524 265 554 297
rect 414 249 554 265
rect 414 215 424 249
rect 458 215 554 249
rect 414 199 554 215
rect 440 177 470 199
rect 524 177 554 199
rect 79 27 109 53
rect 258 27 288 53
rect 342 27 372 53
rect 440 21 470 47
rect 524 21 554 47
<< polycont >>
rect 184 439 218 473
rect 35 215 69 249
rect 226 215 260 249
rect 424 215 458 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 17 349 69 527
rect 382 485 438 527
rect 108 473 346 483
rect 108 439 184 473
rect 218 439 346 473
rect 108 417 346 439
rect 382 451 395 485
rect 429 451 438 485
rect 382 417 438 451
rect 382 383 395 417
rect 429 383 438 417
rect 17 315 35 349
rect 17 299 69 315
rect 119 343 153 377
rect 119 265 153 309
rect 197 354 281 383
rect 382 367 438 383
rect 480 454 526 493
rect 514 420 526 454
rect 480 386 526 420
rect 197 320 226 354
rect 260 333 281 354
rect 514 352 526 386
rect 260 320 446 333
rect 197 299 446 320
rect 480 299 526 352
rect 412 265 446 299
rect 17 249 85 265
rect 17 215 35 249
rect 69 215 85 249
rect 119 249 266 265
rect 119 215 226 249
rect 260 215 266 249
rect 119 199 266 215
rect 412 249 458 265
rect 412 215 424 249
rect 412 199 458 215
rect 119 181 168 199
rect 21 147 168 181
rect 412 165 446 199
rect 21 106 84 147
rect 298 131 446 165
rect 492 152 526 299
rect 560 483 611 527
rect 560 449 564 483
rect 598 449 611 483
rect 560 415 611 449
rect 560 381 564 415
rect 598 381 611 415
rect 560 347 611 381
rect 560 313 564 347
rect 598 313 611 347
rect 560 292 611 313
rect 480 135 526 152
rect 21 72 35 106
rect 69 72 84 106
rect 21 53 84 72
rect 118 97 264 113
rect 118 63 119 97
rect 153 63 214 97
rect 248 63 264 97
rect 118 17 264 63
rect 298 111 332 131
rect 514 101 526 135
rect 298 61 332 77
rect 366 63 392 97
rect 426 63 442 97
rect 480 83 526 101
rect 560 162 611 185
rect 560 128 564 162
rect 598 128 611 162
rect 560 94 611 128
rect 366 17 442 63
rect 560 60 564 94
rect 598 60 611 94
rect 560 17 611 60
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
flabel locali s 213 425 247 459 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 400 0 0 0 B_N
port 2 nsew signal input
flabel locali s 489 357 523 391 0 FreeSans 400 0 0 0 X
port 7 nsew signal output
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 or2b_2
rlabel metal1 s 0 -48 644 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 644 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 644 544
string GDS_END 1004888
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 999424
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 3.220 0.000 
<< end >>
