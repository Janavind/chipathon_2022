magic
tech sky130A
magscale 1 2
timestamp 1666199351
<< pwell >>
rect 256 567 277 616
<< obsli1 >>
rect 13 0 47 2220
rect 493 0 527 2220
<< obsm1 >>
rect 14 2154 526 2220
rect 14 126 46 2154
rect 74 66 106 2094
rect 134 126 166 2154
rect 194 66 226 2094
rect 254 126 286 2154
rect 314 66 346 2094
rect 374 126 406 2154
rect 434 66 466 2094
rect 494 126 526 2154
rect 60 0 480 66
<< obsm2 >>
rect 14 2154 166 2220
rect 14 126 46 2154
rect 74 66 106 2094
rect 134 126 166 2154
rect 194 66 226 2220
rect 254 2154 526 2220
rect 254 126 286 2154
rect 314 66 346 2094
rect 374 126 406 2154
rect 434 66 466 2094
rect 494 126 526 2154
rect 60 0 480 66
<< obsm3 >>
rect 0 2154 540 2220
rect 0 126 60 2154
rect 120 66 180 2094
rect 240 126 300 2154
rect 360 66 420 2094
rect 480 126 540 2154
rect 60 0 480 66
<< metal4 >>
rect 0 2154 540 2220
rect 0 126 60 2154
rect 120 66 180 2094
rect 240 126 300 2154
rect 360 66 420 2094
rect 480 126 540 2154
rect 60 0 480 66
<< labels >>
rlabel metal4 s 480 126 540 2154 6 C0
port 1 nsew
rlabel metal4 s 240 126 300 2154 6 C0
port 1 nsew
rlabel metal4 s 0 2154 540 2220 6 C0
port 1 nsew
rlabel metal4 s 0 126 60 2154 6 C0
port 1 nsew
rlabel metal4 s 360 66 420 2094 6 C1
port 2 nsew
rlabel metal4 s 120 66 180 2094 6 C1
port 2 nsew
rlabel metal4 s 60 0 480 66 6 C1
port 2 nsew
rlabel pwell s 256 567 277 616 6 SUB
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 540 2220
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 18284
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 10556
string device primitive
<< end >>
