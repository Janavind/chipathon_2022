magic
tech sky130B
magscale 1 2
timestamp 1666199351
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 1 67 919 203
rect 1 21 727 67
rect 30 -17 64 21
<< scnmos >>
rect 83 47 113 177
rect 167 47 197 177
rect 251 47 281 177
rect 335 47 365 177
rect 531 47 561 177
rect 615 47 645 177
rect 811 93 841 177
<< scpmoshvt >>
rect 83 297 113 497
rect 167 297 197 497
rect 251 297 281 497
rect 335 297 365 497
rect 531 297 561 497
rect 615 297 645 497
rect 811 297 841 381
<< ndiff >>
rect 27 163 83 177
rect 27 129 39 163
rect 73 129 83 163
rect 27 95 83 129
rect 27 61 39 95
rect 73 61 83 95
rect 27 47 83 61
rect 113 163 167 177
rect 113 129 123 163
rect 157 129 167 163
rect 113 95 167 129
rect 113 61 123 95
rect 157 61 167 95
rect 113 47 167 61
rect 197 95 251 177
rect 197 61 207 95
rect 241 61 251 95
rect 197 47 251 61
rect 281 163 335 177
rect 281 129 291 163
rect 325 129 335 163
rect 281 95 335 129
rect 281 61 291 95
rect 325 61 335 95
rect 281 47 335 61
rect 365 95 417 177
rect 365 61 375 95
rect 409 61 417 95
rect 365 47 417 61
rect 479 95 531 177
rect 479 61 487 95
rect 521 61 531 95
rect 479 47 531 61
rect 561 163 615 177
rect 561 129 571 163
rect 605 129 615 163
rect 561 95 615 129
rect 561 61 571 95
rect 605 61 615 95
rect 561 47 615 61
rect 645 163 701 177
rect 645 129 655 163
rect 689 129 701 163
rect 645 95 701 129
rect 645 61 655 95
rect 689 61 701 95
rect 759 149 811 177
rect 759 115 767 149
rect 801 115 811 149
rect 759 93 811 115
rect 841 149 893 177
rect 841 115 851 149
rect 885 115 893 149
rect 841 93 893 115
rect 645 47 701 61
<< pdiff >>
rect 27 477 83 497
rect 27 443 39 477
rect 73 443 83 477
rect 27 409 83 443
rect 27 375 39 409
rect 73 375 83 409
rect 27 341 83 375
rect 27 307 39 341
rect 73 307 83 341
rect 27 297 83 307
rect 113 477 167 497
rect 113 443 123 477
rect 157 443 167 477
rect 113 409 167 443
rect 113 375 123 409
rect 157 375 167 409
rect 113 297 167 375
rect 197 477 251 497
rect 197 443 207 477
rect 241 443 251 477
rect 197 409 251 443
rect 197 375 207 409
rect 241 375 251 409
rect 197 341 251 375
rect 197 307 207 341
rect 241 307 251 341
rect 197 297 251 307
rect 281 477 335 497
rect 281 443 291 477
rect 325 443 335 477
rect 281 409 335 443
rect 281 375 291 409
rect 325 375 335 409
rect 281 297 335 375
rect 365 409 421 497
rect 365 375 375 409
rect 409 375 421 409
rect 365 341 421 375
rect 365 307 375 341
rect 409 307 421 341
rect 365 297 421 307
rect 475 477 531 497
rect 475 443 487 477
rect 521 443 531 477
rect 475 409 531 443
rect 475 375 487 409
rect 521 375 531 409
rect 475 341 531 375
rect 475 307 487 341
rect 521 307 531 341
rect 475 297 531 307
rect 561 409 615 497
rect 561 375 571 409
rect 605 375 615 409
rect 561 341 615 375
rect 561 307 571 341
rect 605 307 615 341
rect 561 297 615 307
rect 645 477 701 497
rect 645 443 655 477
rect 689 443 701 477
rect 645 409 701 443
rect 645 375 655 409
rect 689 375 701 409
rect 645 341 701 375
rect 645 307 655 341
rect 689 307 701 341
rect 645 297 701 307
rect 759 358 811 381
rect 759 324 767 358
rect 801 324 811 358
rect 759 297 811 324
rect 841 358 893 381
rect 841 324 851 358
rect 885 324 893 358
rect 841 297 893 324
<< ndiffc >>
rect 39 129 73 163
rect 39 61 73 95
rect 123 129 157 163
rect 123 61 157 95
rect 207 61 241 95
rect 291 129 325 163
rect 291 61 325 95
rect 375 61 409 95
rect 487 61 521 95
rect 571 129 605 163
rect 571 61 605 95
rect 655 129 689 163
rect 655 61 689 95
rect 767 115 801 149
rect 851 115 885 149
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 39 307 73 341
rect 123 443 157 477
rect 123 375 157 409
rect 207 443 241 477
rect 207 375 241 409
rect 207 307 241 341
rect 291 443 325 477
rect 291 375 325 409
rect 375 375 409 409
rect 375 307 409 341
rect 487 443 521 477
rect 487 375 521 409
rect 487 307 521 341
rect 571 375 605 409
rect 571 307 605 341
rect 655 443 689 477
rect 655 375 689 409
rect 655 307 689 341
rect 767 324 801 358
rect 851 324 885 358
<< poly >>
rect 83 497 113 523
rect 167 497 197 523
rect 251 497 281 523
rect 335 497 365 523
rect 531 497 561 523
rect 615 497 645 523
rect 811 381 841 407
rect 83 265 113 297
rect 167 265 197 297
rect 83 249 197 265
rect 83 215 112 249
rect 146 215 197 249
rect 83 199 197 215
rect 83 177 113 199
rect 167 177 197 199
rect 251 265 281 297
rect 335 265 365 297
rect 251 249 365 265
rect 251 215 288 249
rect 322 215 365 249
rect 251 199 365 215
rect 251 177 281 199
rect 335 177 365 199
rect 531 265 561 297
rect 615 265 645 297
rect 811 265 841 297
rect 531 249 707 265
rect 531 215 663 249
rect 697 215 707 249
rect 531 199 707 215
rect 811 249 866 265
rect 811 215 822 249
rect 856 215 866 249
rect 811 199 866 215
rect 531 177 561 199
rect 615 177 645 199
rect 811 177 841 199
rect 811 67 841 93
rect 83 21 113 47
rect 167 21 197 47
rect 251 21 281 47
rect 335 21 365 47
rect 531 21 561 47
rect 615 21 645 47
<< polycont >>
rect 112 215 146 249
rect 288 215 322 249
rect 663 215 697 249
rect 822 215 856 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 18 477 81 493
rect 18 443 39 477
rect 73 443 81 477
rect 18 409 81 443
rect 18 375 39 409
rect 73 375 81 409
rect 18 341 81 375
rect 115 477 165 527
rect 115 443 123 477
rect 157 443 165 477
rect 115 409 165 443
rect 115 375 123 409
rect 157 375 165 409
rect 115 359 165 375
rect 199 477 249 493
rect 199 443 207 477
rect 241 443 249 477
rect 199 409 249 443
rect 199 375 207 409
rect 241 375 249 409
rect 18 307 39 341
rect 73 325 81 341
rect 199 341 249 375
rect 283 477 696 493
rect 283 443 291 477
rect 325 459 487 477
rect 325 443 333 459
rect 283 409 333 443
rect 475 443 487 459
rect 521 459 655 477
rect 521 443 529 459
rect 283 375 291 409
rect 325 375 333 409
rect 283 359 333 375
rect 367 409 417 425
rect 367 375 375 409
rect 409 375 417 409
rect 199 325 207 341
rect 73 307 207 325
rect 241 325 249 341
rect 367 341 417 375
rect 367 325 375 341
rect 241 307 375 325
rect 409 307 417 341
rect 18 291 417 307
rect 475 409 529 443
rect 647 443 655 459
rect 689 443 696 477
rect 475 375 487 409
rect 521 375 529 409
rect 475 341 529 375
rect 475 307 487 341
rect 521 307 529 341
rect 475 291 529 307
rect 563 409 613 425
rect 563 375 571 409
rect 605 375 613 409
rect 563 341 613 375
rect 563 307 571 341
rect 605 307 613 341
rect 22 249 193 257
rect 22 215 112 249
rect 146 215 193 249
rect 227 249 528 257
rect 227 215 288 249
rect 322 215 528 249
rect 563 181 613 307
rect 647 409 696 443
rect 647 375 655 409
rect 689 375 696 409
rect 647 341 696 375
rect 647 307 655 341
rect 689 307 696 341
rect 647 291 696 307
rect 738 358 809 374
rect 738 324 767 358
rect 801 324 809 358
rect 738 291 809 324
rect 843 358 893 527
rect 843 324 851 358
rect 885 324 893 358
rect 843 308 893 324
rect 738 257 772 291
rect 647 249 772 257
rect 647 215 663 249
rect 697 215 772 249
rect 806 249 903 257
rect 806 215 822 249
rect 856 215 903 249
rect 738 181 772 215
rect 18 163 73 181
rect 18 129 39 163
rect 18 95 73 129
rect 18 61 39 95
rect 18 17 73 61
rect 107 163 621 181
rect 107 129 123 163
rect 157 145 291 163
rect 157 129 173 145
rect 107 95 173 129
rect 275 129 291 145
rect 325 145 571 163
rect 325 129 341 145
rect 107 61 123 95
rect 157 61 173 95
rect 107 51 173 61
rect 207 95 241 111
rect 207 17 241 61
rect 275 95 341 129
rect 555 129 571 145
rect 605 129 621 163
rect 275 61 291 95
rect 325 61 341 95
rect 275 51 341 61
rect 375 95 521 111
rect 409 61 487 95
rect 375 17 521 61
rect 555 95 621 129
rect 555 61 571 95
rect 605 61 621 95
rect 555 51 621 61
rect 655 163 696 179
rect 689 129 696 163
rect 655 95 696 129
rect 689 61 696 95
rect 738 149 809 181
rect 738 115 767 149
rect 801 115 809 149
rect 738 76 809 115
rect 843 149 901 165
rect 843 115 851 149
rect 885 115 901 149
rect 655 17 696 61
rect 843 17 901 115
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
flabel locali s 857 221 891 255 0 FreeSans 400 0 0 0 C_N
port 3 nsew signal input
flabel locali s 586 85 620 119 0 FreeSans 400 0 0 0 Y
port 8 nsew signal output
flabel locali s 122 221 156 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 306 221 340 255 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 nor3b_2
rlabel metal1 s 0 -48 920 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 920 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 920 544
string GDS_END 1117960
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1110144
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 4.600 0.000 
<< end >>
