magic
tech sky130A
magscale 1 2
timestamp 1666199351
<< poly >>
rect 721 3500 1121 3516
rect 721 3398 768 3500
rect 1074 3398 1121 3500
rect 721 2896 768 2998
rect 1074 2896 1121 2998
rect 721 2194 768 2296
rect 1074 2194 1121 2296
rect 721 1092 768 1194
rect 1074 1092 1121 1194
rect 721 1072 1121 1092
<< polycont >>
rect 768 3398 1074 3500
rect 768 2896 1074 2998
rect 768 2194 1074 2296
rect 768 1092 1074 1194
<< npolyres >>
rect 721 2998 1121 3398
rect 721 2296 1121 2896
rect 721 1194 1121 2194
<< locali >>
rect 2853 11344 2925 11378
rect 2127 11308 2187 11342
rect 2093 11261 2221 11308
rect 2127 11227 2187 11261
rect 2093 11180 2221 11227
rect 2127 11146 2187 11180
rect 2093 11099 2221 11146
rect 2127 11065 2187 11099
rect 2093 11019 2221 11065
rect 2127 10985 2187 11019
rect 2819 11305 2959 11344
rect 2853 11271 2925 11305
rect 2819 11233 2959 11271
rect 2853 11199 2925 11233
rect 2819 11161 2959 11199
rect 2853 11127 2925 11161
rect 2819 11089 2959 11127
rect 2853 11055 2925 11089
rect 2819 11017 2959 11055
rect 2853 10983 2925 11017
rect 752 3514 1090 3516
rect 752 3480 753 3514
rect 787 3500 828 3514
rect 862 3500 903 3514
rect 937 3500 979 3514
rect 1013 3500 1055 3514
rect 1089 3480 1090 3514
rect 752 3420 768 3480
rect 1074 3420 1090 3480
rect 752 3386 753 3420
rect 787 3386 828 3398
rect 862 3386 903 3398
rect 937 3386 979 3398
rect 1013 3386 1055 3398
rect 1089 3386 1090 3420
rect 752 3382 1090 3386
rect 752 2978 760 3012
rect 794 2998 863 3012
rect 897 2998 966 3012
rect 1000 2998 1090 3012
rect 752 2930 768 2978
rect 752 2896 760 2930
rect 1074 2896 1090 2998
rect 752 2294 768 2296
rect 752 2260 760 2294
rect 752 2212 768 2260
rect 752 2178 760 2212
rect 1074 2194 1090 2296
rect 794 2178 863 2194
rect 897 2178 966 2194
rect 1000 2178 1090 2194
rect 752 1197 1090 1210
rect 752 1091 753 1197
rect 1075 1091 1090 1197
rect 752 1076 1090 1091
<< viali >>
rect 2819 11344 2853 11378
rect 2925 11344 2959 11378
rect 2093 11308 2127 11342
rect 2187 11308 2221 11342
rect 2093 11227 2127 11261
rect 2187 11227 2221 11261
rect 2093 11146 2127 11180
rect 2187 11146 2221 11180
rect 2093 11065 2127 11099
rect 2187 11065 2221 11099
rect 2093 10985 2127 11019
rect 2187 10985 2221 11019
rect 2819 11271 2853 11305
rect 2925 11271 2959 11305
rect 2819 11199 2853 11233
rect 2925 11199 2959 11233
rect 2819 11127 2853 11161
rect 2925 11127 2959 11161
rect 2819 11055 2853 11089
rect 2925 11055 2959 11089
rect 2819 10983 2853 11017
rect 2925 10983 2959 11017
rect 753 3500 787 3514
rect 828 3500 862 3514
rect 903 3500 937 3514
rect 979 3500 1013 3514
rect 1055 3500 1089 3514
rect 753 3480 768 3500
rect 768 3480 787 3500
rect 828 3480 862 3500
rect 903 3480 937 3500
rect 979 3480 1013 3500
rect 1055 3480 1074 3500
rect 1074 3480 1089 3500
rect 753 3398 768 3420
rect 768 3398 787 3420
rect 828 3398 862 3420
rect 903 3398 937 3420
rect 979 3398 1013 3420
rect 1055 3398 1074 3420
rect 1074 3398 1089 3420
rect 753 3386 787 3398
rect 828 3386 862 3398
rect 903 3386 937 3398
rect 979 3386 1013 3398
rect 1055 3386 1089 3398
rect 760 2998 794 3012
rect 863 2998 897 3012
rect 966 2998 1000 3012
rect 760 2978 768 2998
rect 768 2978 794 2998
rect 863 2978 897 2998
rect 966 2978 1000 2998
rect 760 2896 768 2930
rect 768 2896 794 2930
rect 863 2896 897 2930
rect 966 2896 1000 2930
rect 760 2260 768 2294
rect 768 2260 794 2294
rect 863 2260 897 2294
rect 966 2260 1000 2294
rect 760 2194 768 2212
rect 768 2194 794 2212
rect 863 2194 897 2212
rect 966 2194 1000 2212
rect 760 2178 794 2194
rect 863 2178 897 2194
rect 966 2178 1000 2194
rect 753 1194 1075 1197
rect 753 1092 768 1194
rect 768 1092 1074 1194
rect 1074 1092 1075 1194
rect 753 1091 1075 1092
<< metal1 >>
rect 18589 20683 18620 20750
rect 4117 20425 4271 20431
rect 4169 20373 4271 20425
rect 4117 20361 4271 20373
rect 4169 20353 4271 20361
rect 4117 20303 4169 20309
tri 4169 20303 4219 20353 nw
rect 2648 16599 2694 16651
rect 3025 12926 3099 13014
rect 6438 11647 6540 11736
rect 2515 11386 2965 11390
rect 2087 11342 2227 11354
rect 2087 11308 2093 11342
rect 2127 11308 2187 11342
rect 2221 11308 2227 11342
rect 2087 11261 2227 11308
rect 2087 11227 2093 11261
rect 2127 11227 2187 11261
rect 2221 11238 2227 11261
rect 2515 11334 2521 11386
rect 2573 11334 2608 11386
rect 2660 11334 2694 11386
rect 2746 11378 2965 11386
rect 2746 11344 2819 11378
rect 2853 11344 2925 11378
rect 2959 11344 2965 11378
rect 2746 11334 2965 11344
rect 2515 11305 2965 11334
rect 2515 11294 2819 11305
rect 2515 11242 2521 11294
rect 2573 11242 2608 11294
rect 2660 11242 2694 11294
rect 2746 11271 2819 11294
rect 2853 11271 2925 11305
rect 2959 11271 2965 11305
rect 2746 11242 2965 11271
tri 2227 11238 2230 11241 sw
rect 2515 11238 2965 11242
rect 2221 11233 2230 11238
tri 2230 11233 2235 11238 sw
rect 2813 11233 2965 11238
rect 2221 11227 2235 11233
rect 2087 11199 2235 11227
tri 2235 11199 2269 11233 sw
rect 2813 11199 2819 11233
rect 2853 11199 2925 11233
rect 2959 11199 2965 11233
rect 2087 11180 2269 11199
rect 2087 11146 2093 11180
rect 2127 11146 2187 11180
rect 2221 11172 2269 11180
tri 2269 11172 2296 11199 sw
rect 2221 11146 2393 11172
rect 2087 11120 2393 11146
rect 2445 11120 2473 11172
rect 2525 11120 2552 11172
rect 2604 11120 2631 11172
rect 2683 11120 2710 11172
rect 2762 11120 2768 11172
rect 2087 11108 2768 11120
rect 2087 11099 2393 11108
rect 2087 11065 2093 11099
rect 2127 11065 2187 11099
rect 2221 11065 2393 11099
rect 2087 11056 2393 11065
rect 2445 11056 2473 11108
rect 2525 11056 2552 11108
rect 2604 11056 2631 11108
rect 2683 11056 2710 11108
rect 2762 11056 2768 11108
rect 2813 11161 2965 11199
rect 2813 11127 2819 11161
rect 2853 11127 2925 11161
rect 2959 11127 2965 11161
rect 2813 11089 2965 11127
rect 2087 11055 2295 11056
tri 2295 11055 2296 11056 nw
rect 2813 11055 2819 11089
rect 2853 11055 2925 11089
rect 2959 11055 2965 11089
rect 2087 11019 2257 11055
rect 2087 10985 2093 11019
rect 2127 10985 2187 11019
rect 2221 11017 2257 11019
tri 2257 11017 2295 11055 nw
rect 2813 11017 2965 11055
rect 2221 10985 2227 11017
tri 2227 10987 2257 11017 nw
rect 2087 10973 2227 10985
rect 2813 10983 2819 11017
rect 2853 10983 2925 11017
rect 2959 10983 2965 11017
rect 2813 10971 2965 10983
rect 7198 11048 8251 11062
rect 7198 10996 7204 11048
rect 7256 10996 7287 11048
rect 7339 10996 7370 11048
rect 7422 10996 7453 11048
rect 7505 10996 7536 11048
rect 7588 10996 7619 11048
rect 7671 10996 7701 11048
rect 7753 10996 7783 11048
rect 7835 10996 7865 11048
rect 7917 10996 7947 11048
rect 7999 10996 8029 11048
rect 8081 10996 8111 11048
rect 8163 10996 8193 11048
rect 8245 10996 8251 11048
rect 7198 10982 8251 10996
tri 2366 10593 2387 10614 se
rect 2387 10612 2768 10614
rect 2387 10593 2393 10612
tri 1077 10517 1153 10593 se
rect 1153 10560 2393 10593
rect 2445 10560 2473 10612
rect 2525 10560 2552 10612
rect 2604 10560 2631 10612
rect 2683 10560 2710 10612
rect 2762 10560 2768 10612
rect 1153 10542 2768 10560
rect 1153 10517 2393 10542
rect 554 10511 2393 10517
rect 606 10459 618 10511
rect 670 10459 682 10511
rect 734 10459 746 10511
rect 798 10490 2393 10511
rect 2445 10490 2473 10542
rect 2525 10490 2552 10542
rect 2604 10490 2631 10542
rect 2683 10490 2710 10542
rect 2762 10490 2768 10542
rect 798 10472 2768 10490
rect 798 10459 2393 10472
rect 554 10429 2393 10459
rect 606 10377 618 10429
rect 670 10377 682 10429
rect 734 10377 746 10429
rect 798 10420 2393 10429
rect 2445 10420 2473 10472
rect 2525 10420 2552 10472
rect 2604 10420 2631 10472
rect 2683 10420 2710 10472
rect 2762 10420 2768 10472
rect 798 10402 2768 10420
rect 798 10377 2393 10402
rect 554 10350 2393 10377
rect 2445 10350 2473 10402
rect 2525 10350 2552 10402
rect 2604 10350 2631 10402
rect 2683 10350 2710 10402
rect 2762 10350 2768 10402
rect 554 10346 2768 10350
rect 606 10294 618 10346
rect 670 10294 682 10346
rect 734 10294 746 10346
rect 798 10332 2768 10346
rect 798 10294 2393 10332
rect 554 10280 2393 10294
rect 2445 10280 2473 10332
rect 2525 10280 2552 10332
rect 2604 10280 2631 10332
rect 2683 10280 2710 10332
rect 2762 10280 2768 10332
rect 554 10277 2768 10280
rect 554 10263 2496 10277
rect 606 10211 618 10263
rect 670 10211 682 10263
rect 734 10211 746 10263
rect 798 10211 2496 10263
rect 554 10205 2496 10211
tri 2496 10205 2568 10277 nw
rect 25593 9506 25712 9623
rect 409 8610 415 8726
rect 531 8678 537 8726
rect 531 8610 541 8678
tri 2477 8229 2490 8242 se
rect 2490 8229 3338 8242
rect 2399 8223 3338 8229
rect 2515 8158 3338 8223
rect 2399 8101 2515 8107
rect 26411 8083 26446 8129
tri 26411 8054 26440 8083 ne
rect 26440 8013 26446 8083
rect 26562 8013 26568 8129
tri 26698 7972 26704 7978 se
rect 26704 7972 26821 7978
rect 26669 7886 26705 7972
tri 26669 7850 26705 7886 ne
rect 26705 7850 26821 7856
tri 26555 7306 26599 7350 se
rect 26599 7306 26605 7350
rect 24520 7190 24526 7306
rect 24642 7234 26605 7306
rect 26721 7234 26727 7350
rect 24642 7190 24648 7234
tri 24648 7190 24692 7234 nw
rect 3667 6447 3717 6497
rect 10742 5629 10937 5723
tri 343 5111 382 5150 se
rect 382 5144 498 5150
tri 330 5098 343 5111 se
rect 343 5098 382 5111
rect 330 4964 382 5098
tri 498 5077 532 5111 sw
rect 498 4964 532 5077
rect 330 4958 532 4964
rect 3629 4839 3739 4967
rect 24718 4674 24764 4720
rect 741 3632 747 3684
rect 799 3632 827 3684
rect 879 3632 906 3684
rect 958 3632 985 3684
rect 1037 3632 1064 3684
rect 1116 3632 1122 3684
rect 741 3600 1122 3632
rect 741 3548 747 3600
rect 799 3548 827 3600
rect 879 3548 906 3600
rect 958 3548 985 3600
rect 1037 3548 1064 3600
rect 1116 3548 1122 3600
rect 24021 3550 24066 3596
rect 741 3516 1122 3548
rect 741 3464 747 3516
rect 799 3464 827 3516
rect 879 3514 906 3516
rect 958 3514 985 3516
rect 1037 3514 1064 3516
rect 879 3480 903 3514
rect 958 3480 979 3514
rect 1037 3480 1055 3514
rect 879 3464 906 3480
rect 958 3464 985 3480
rect 1037 3464 1064 3480
rect 1116 3464 1122 3516
rect 741 3432 1122 3464
rect 741 3380 747 3432
rect 799 3380 827 3432
rect 879 3420 906 3432
rect 958 3420 985 3432
rect 1037 3420 1064 3432
rect 879 3386 903 3420
rect 958 3386 979 3420
rect 1037 3386 1055 3420
rect 879 3380 906 3386
rect 958 3380 985 3386
rect 1037 3380 1064 3386
rect 1116 3380 1122 3432
rect 748 3012 1012 3018
rect 748 2978 760 3012
rect 794 2978 863 3012
rect 897 2978 966 3012
rect 1000 2978 1012 3012
rect 748 2930 1012 2978
rect 748 2896 760 2930
rect 794 2896 863 2930
rect 897 2896 966 2930
rect 1000 2896 1012 2930
rect 748 2767 1012 2896
rect 749 2765 1011 2766
rect 748 2465 1012 2765
rect 749 2464 1011 2465
rect 748 2294 1012 2463
rect 748 2260 760 2294
rect 794 2260 863 2294
rect 897 2260 966 2294
rect 1000 2260 1012 2294
rect 2384 2271 2528 2439
rect 748 2212 1012 2260
rect 748 2178 760 2212
rect 794 2178 863 2212
rect 897 2178 966 2212
rect 1000 2178 1012 2212
rect 748 2172 1012 2178
rect 747 1744 753 1796
rect 805 1744 842 1796
rect 894 1744 932 1796
rect 984 1744 1022 1796
rect 1074 1744 1081 1796
rect 747 1728 1081 1744
rect 747 1676 753 1728
rect 805 1676 842 1728
rect 894 1676 932 1728
rect 984 1676 1022 1728
rect 1074 1676 1081 1728
rect 747 1197 1081 1676
rect 1991 1303 2116 1444
rect 747 1091 753 1197
rect 1075 1091 1081 1197
rect 747 1079 1081 1091
rect 1538 892 1717 1071
<< rmetal1 >>
rect 748 2766 1012 2767
rect 748 2765 749 2766
rect 1011 2765 1012 2766
rect 748 2464 749 2465
rect 1011 2464 1012 2465
rect 748 2463 1012 2464
<< via1 >>
rect 4117 20373 4169 20425
rect 4117 20309 4169 20361
rect 2521 11334 2573 11386
rect 2608 11334 2660 11386
rect 2694 11334 2746 11386
rect 2521 11242 2573 11294
rect 2608 11242 2660 11294
rect 2694 11242 2746 11294
rect 2393 11120 2445 11172
rect 2473 11120 2525 11172
rect 2552 11120 2604 11172
rect 2631 11120 2683 11172
rect 2710 11120 2762 11172
rect 2393 11056 2445 11108
rect 2473 11056 2525 11108
rect 2552 11056 2604 11108
rect 2631 11056 2683 11108
rect 2710 11056 2762 11108
rect 7204 10996 7256 11048
rect 7287 10996 7339 11048
rect 7370 10996 7422 11048
rect 7453 10996 7505 11048
rect 7536 10996 7588 11048
rect 7619 10996 7671 11048
rect 7701 10996 7753 11048
rect 7783 10996 7835 11048
rect 7865 10996 7917 11048
rect 7947 10996 7999 11048
rect 8029 10996 8081 11048
rect 8111 10996 8163 11048
rect 8193 10996 8245 11048
rect 2393 10560 2445 10612
rect 2473 10560 2525 10612
rect 2552 10560 2604 10612
rect 2631 10560 2683 10612
rect 2710 10560 2762 10612
rect 554 10459 606 10511
rect 618 10459 670 10511
rect 682 10459 734 10511
rect 746 10459 798 10511
rect 2393 10490 2445 10542
rect 2473 10490 2525 10542
rect 2552 10490 2604 10542
rect 2631 10490 2683 10542
rect 2710 10490 2762 10542
rect 554 10377 606 10429
rect 618 10377 670 10429
rect 682 10377 734 10429
rect 746 10377 798 10429
rect 2393 10420 2445 10472
rect 2473 10420 2525 10472
rect 2552 10420 2604 10472
rect 2631 10420 2683 10472
rect 2710 10420 2762 10472
rect 2393 10350 2445 10402
rect 2473 10350 2525 10402
rect 2552 10350 2604 10402
rect 2631 10350 2683 10402
rect 2710 10350 2762 10402
rect 554 10294 606 10346
rect 618 10294 670 10346
rect 682 10294 734 10346
rect 746 10294 798 10346
rect 2393 10280 2445 10332
rect 2473 10280 2525 10332
rect 2552 10280 2604 10332
rect 2631 10280 2683 10332
rect 2710 10280 2762 10332
rect 554 10211 606 10263
rect 618 10211 670 10263
rect 682 10211 734 10263
rect 746 10211 798 10263
rect 415 8610 531 8726
rect 2399 8107 2515 8223
rect 26446 8013 26562 8129
rect 26705 7856 26821 7972
rect 24526 7190 24642 7306
rect 26605 7234 26721 7350
rect 382 4964 498 5144
rect 747 3632 799 3684
rect 827 3632 879 3684
rect 906 3632 958 3684
rect 985 3632 1037 3684
rect 1064 3632 1116 3684
rect 747 3548 799 3600
rect 827 3548 879 3600
rect 906 3548 958 3600
rect 985 3548 1037 3600
rect 1064 3548 1116 3600
rect 747 3514 799 3516
rect 747 3480 753 3514
rect 753 3480 787 3514
rect 787 3480 799 3514
rect 747 3464 799 3480
rect 827 3514 879 3516
rect 906 3514 958 3516
rect 985 3514 1037 3516
rect 1064 3514 1116 3516
rect 827 3480 828 3514
rect 828 3480 862 3514
rect 862 3480 879 3514
rect 906 3480 937 3514
rect 937 3480 958 3514
rect 985 3480 1013 3514
rect 1013 3480 1037 3514
rect 1064 3480 1089 3514
rect 1089 3480 1116 3514
rect 827 3464 879 3480
rect 906 3464 958 3480
rect 985 3464 1037 3480
rect 1064 3464 1116 3480
rect 747 3420 799 3432
rect 747 3386 753 3420
rect 753 3386 787 3420
rect 787 3386 799 3420
rect 747 3380 799 3386
rect 827 3420 879 3432
rect 906 3420 958 3432
rect 985 3420 1037 3432
rect 1064 3420 1116 3432
rect 827 3386 828 3420
rect 828 3386 862 3420
rect 862 3386 879 3420
rect 906 3386 937 3420
rect 937 3386 958 3420
rect 985 3386 1013 3420
rect 1013 3386 1037 3420
rect 1064 3386 1089 3420
rect 1089 3386 1116 3420
rect 827 3380 879 3386
rect 906 3380 958 3386
rect 985 3380 1037 3386
rect 1064 3380 1116 3386
rect 753 1744 805 1796
rect 842 1744 894 1796
rect 932 1744 984 1796
rect 1022 1744 1074 1796
rect 753 1676 805 1728
rect 842 1676 894 1728
rect 932 1676 984 1728
rect 1022 1676 1074 1728
<< metal2 >>
rect 18324 21491 18391 21543
rect 18324 21411 18392 21451
rect 18322 21020 18391 21072
tri 2996 20991 3017 21012 se
rect 3017 20991 4051 21012
tri 4051 20991 4072 21012 sw
tri 2907 20902 2996 20991 se
rect 2996 20930 4072 20991
rect 2996 20902 3023 20930
tri 3023 20902 3051 20930 nw
tri 4017 20902 4045 20930 ne
rect 4045 20902 4072 20930
rect 2907 20875 2996 20902
tri 2996 20875 3023 20902 nw
tri 4045 20875 4072 20902 ne
tri 4072 20875 4188 20991 sw
rect 2907 20373 2989 20875
tri 2989 20868 2996 20875 nw
tri 4072 20868 4079 20875 ne
rect 4079 20868 4188 20875
tri 4079 20830 4117 20868 ne
rect 4117 20425 4188 20868
tri 2989 20373 2992 20376 sw
rect 4169 20373 4188 20425
rect 2907 20362 2992 20373
tri 2992 20362 3003 20373 sw
rect 2907 20361 3003 20362
tri 3003 20361 3004 20362 sw
rect 4117 20361 4188 20373
rect 2907 20342 3004 20361
tri 3004 20342 3023 20361 sw
tri 2907 20309 2940 20342 ne
rect 2940 20322 3023 20342
tri 3023 20322 3043 20342 sw
rect 2940 20309 3309 20322
tri 3309 20309 3322 20322 sw
rect 4169 20309 4188 20361
rect 18320 20353 18405 20431
tri 2940 20303 2946 20309 ne
rect 2946 20303 3322 20309
tri 3322 20303 3328 20309 sw
rect 4117 20303 4188 20309
tri 2946 20246 3003 20303 ne
rect 3003 20293 3328 20303
tri 3328 20293 3338 20303 sw
rect 3003 20246 3338 20293
tri 3338 20246 3385 20293 sw
tri 3279 20206 3319 20246 ne
rect 3319 20217 3385 20246
tri 3385 20217 3414 20246 sw
rect 3319 20206 3414 20217
rect 368 20197 506 20206
rect 368 20061 370 20197
tri 506 20176 536 20206 sw
tri 3319 20187 3338 20206 ne
rect 506 20061 794 20176
rect 368 20056 794 20061
rect 368 20052 506 20056
tri 506 20052 510 20056 nw
rect 144 20037 288 20046
rect 144 19901 152 20037
tri 288 20016 318 20046 sw
rect 288 19901 794 20016
rect 144 19896 794 19901
tri 144 19892 148 19896 ne
rect 148 19892 288 19896
tri 288 19892 292 19896 nw
tri 3245 18143 3338 18236 se
rect 3338 18206 3414 20206
rect 3338 18143 3351 18206
tri 3351 18143 3414 18206 nw
rect 2406 18092 3300 18143
tri 3300 18092 3351 18143 nw
rect 2406 18083 3275 18092
rect 2406 18067 2411 18083
rect 2467 18067 3275 18083
tri 3275 18067 3300 18092 nw
rect 2411 18003 2467 18027
rect 2411 17938 2467 17947
rect 2515 11946 2540 12002
rect 2596 11946 2661 12002
rect 2717 11946 2766 12002
rect 2515 11922 2766 11946
rect 2515 11866 2540 11922
rect 2596 11866 2661 11922
rect 2717 11866 2766 11922
rect 2515 11842 2766 11866
rect 2515 11786 2540 11842
rect 2596 11786 2661 11842
rect 2717 11786 2766 11842
rect 2515 11386 2766 11786
rect 2515 11334 2521 11386
rect 2573 11334 2608 11386
rect 2660 11334 2694 11386
rect 2746 11334 2766 11386
rect 2515 11294 2766 11334
rect 2515 11242 2521 11294
rect 2573 11242 2608 11294
rect 2660 11242 2694 11294
rect 2746 11242 2766 11294
rect 2370 11172 2768 11184
rect 2370 11120 2393 11172
rect 2445 11120 2473 11172
rect 2525 11120 2552 11172
rect 2604 11120 2631 11172
rect 2683 11120 2710 11172
rect 2762 11120 2768 11172
rect 2370 11108 2768 11120
rect 2370 11056 2393 11108
rect 2445 11056 2473 11108
rect 2525 11056 2552 11108
rect 2604 11056 2631 11108
rect 2683 11056 2710 11108
rect 2762 11056 2768 11108
rect 2370 10612 2768 11056
rect 7197 11051 8251 11062
rect 7197 11048 7206 11051
rect 7262 11048 7288 11051
rect 7197 10996 7204 11048
rect 7262 10996 7287 11048
rect 7197 10995 7206 10996
rect 7262 10995 7288 10996
rect 7344 10995 7370 11051
rect 7426 10995 7452 11051
rect 7508 10995 7534 11051
rect 7590 10995 7616 11051
rect 7672 10995 7698 11051
rect 7754 10995 7780 11051
rect 7836 10995 7862 11051
rect 7918 10995 7944 11051
rect 8000 10995 8025 11051
rect 8081 10995 8106 11051
rect 8162 11048 8187 11051
rect 8243 11048 8252 11051
rect 8163 10996 8187 11048
rect 8245 10996 8252 11048
rect 8162 10995 8187 10996
rect 8243 10995 8252 10996
rect 7197 10982 8251 10995
rect 2370 10560 2393 10612
rect 2445 10560 2473 10612
rect 2525 10560 2552 10612
rect 2604 10560 2631 10612
rect 2683 10560 2710 10612
rect 2762 10560 2768 10612
rect 2370 10542 2768 10560
rect 554 10511 798 10517
rect 606 10459 618 10511
rect 670 10459 682 10511
rect 734 10459 746 10511
rect 554 10429 798 10459
rect 606 10377 618 10429
rect 670 10377 682 10429
rect 734 10377 746 10429
rect 554 10346 798 10377
rect 606 10294 618 10346
rect 670 10294 682 10346
rect 734 10294 746 10346
rect 554 10263 798 10294
rect 606 10211 618 10263
rect 670 10211 682 10263
rect 734 10211 746 10263
tri 515 8726 554 8765 se
rect 554 8726 798 10211
rect 409 8610 415 8726
rect 531 8610 798 8726
tri 523 8579 554 8610 ne
rect 368 5182 504 5191
rect 368 4964 382 4966
rect 498 4964 504 4966
rect 368 4957 504 4964
rect 554 3684 798 8610
rect 2370 10490 2393 10542
rect 2445 10490 2473 10542
rect 2525 10490 2552 10542
rect 2604 10490 2631 10542
rect 2683 10490 2710 10542
rect 2762 10490 2768 10542
rect 2370 10472 2768 10490
rect 2370 10420 2393 10472
rect 2445 10420 2473 10472
rect 2525 10420 2552 10472
rect 2604 10420 2631 10472
rect 2683 10420 2710 10472
rect 2762 10420 2768 10472
rect 2370 10402 2768 10420
rect 2370 10350 2393 10402
rect 2445 10350 2473 10402
rect 2525 10350 2552 10402
rect 2604 10350 2631 10402
rect 2683 10350 2710 10402
rect 2762 10350 2768 10402
rect 2370 10332 2768 10350
rect 2370 10280 2393 10332
rect 2445 10280 2473 10332
rect 2525 10280 2552 10332
rect 2604 10280 2631 10332
rect 2683 10280 2710 10332
rect 2762 10280 2768 10332
rect 2370 10277 2768 10280
rect 2370 8260 2498 10277
tri 2498 10191 2584 10277 nw
rect 25972 10001 26779 10049
tri 26779 10001 26827 10049 sw
rect 25972 9921 26827 10001
tri 26658 9873 26706 9921 ne
rect 26023 9770 26536 9818
tri 26536 9770 26584 9818 sw
rect 26023 9690 26584 9770
tri 26400 9657 26433 9690 ne
tri 2498 8260 2515 8277 sw
rect 2370 8223 2515 8260
rect 2370 8107 2399 8223
rect 2370 8101 2515 8107
rect 26433 8129 26584 9690
rect 2905 7979 2957 8017
rect 26433 8013 26446 8129
rect 26562 8013 26584 8129
rect 2813 7932 2865 7966
rect 3674 7709 3753 7759
rect 26433 7350 26584 8013
tri 26674 7978 26706 8010 se
rect 26706 7978 26827 9921
rect 26652 7972 26827 7978
rect 26652 7856 26705 7972
rect 26821 7856 26827 7972
rect 26652 7850 26827 7856
tri 26584 7350 26658 7424 sw
rect 24520 7190 24526 7306
rect 24642 7190 24648 7306
rect 26433 7234 26605 7350
rect 26721 7234 26727 7350
rect 3092 7071 3139 7121
rect 2815 6972 2863 7022
rect 2537 6045 2589 6123
rect 3951 5695 4002 5740
tri 798 3684 945 3831 sw
rect 554 3632 747 3684
rect 799 3632 827 3684
rect 879 3632 906 3684
rect 958 3632 985 3684
rect 1037 3632 1064 3684
rect 1116 3632 1122 3684
rect 554 3600 1122 3632
rect 554 3548 747 3600
rect 799 3548 827 3600
rect 879 3548 906 3600
rect 958 3548 985 3600
rect 1037 3548 1064 3600
rect 1116 3548 1122 3600
rect 554 3516 1122 3548
rect 554 3464 747 3516
rect 799 3464 827 3516
rect 879 3464 906 3516
rect 958 3464 985 3516
rect 1037 3464 1064 3516
rect 1116 3464 1122 3516
rect 554 3432 1122 3464
rect 554 3380 747 3432
rect 799 3380 827 3432
rect 879 3380 906 3432
rect 958 3380 985 3432
rect 1037 3380 1064 3432
rect 1116 3380 1122 3432
rect 364 2799 513 2808
rect 420 2743 448 2799
rect 504 2758 513 2799
tri 513 2758 563 2808 sw
rect 504 2743 1258 2758
rect 364 2708 1258 2743
rect 420 2652 448 2708
rect 504 2652 1258 2708
rect 364 2616 1258 2652
rect 420 2560 448 2616
rect 504 2560 1258 2616
rect 364 2551 1258 2560
rect 148 2418 1244 2427
rect 148 2362 149 2418
rect 205 2362 233 2418
rect 289 2362 1244 2418
rect 148 2327 1244 2362
rect 148 2271 149 2327
rect 205 2271 233 2327
rect 289 2271 1244 2327
rect 148 2235 1244 2271
rect 148 2179 149 2235
rect 205 2179 233 2235
rect 289 2179 1244 2235
rect 148 2170 1244 2179
tri 686 2109 747 2170 ne
rect 747 1796 1080 2170
tri 1080 2109 1141 2170 nw
rect 747 1744 753 1796
rect 805 1744 842 1796
rect 894 1744 932 1796
rect 984 1744 1022 1796
rect 1074 1744 1080 1796
rect 747 1728 1080 1744
rect 747 1676 753 1728
rect 805 1676 842 1728
rect 894 1676 932 1728
rect 984 1676 1022 1728
rect 1074 1676 1080 1728
rect 2587 -2362 2643 -2353
rect 2587 -2442 2643 -2418
rect 2587 -2507 2643 -2498
<< via2 >>
rect 370 20061 506 20197
rect 152 19901 288 20037
rect 2411 18027 2467 18083
rect 2411 17947 2467 18003
rect 2540 11946 2596 12002
rect 2661 11946 2717 12002
rect 2540 11866 2596 11922
rect 2661 11866 2717 11922
rect 2540 11786 2596 11842
rect 2661 11786 2717 11842
rect 7206 11048 7262 11051
rect 7288 11048 7344 11051
rect 7206 10996 7256 11048
rect 7256 10996 7262 11048
rect 7288 10996 7339 11048
rect 7339 10996 7344 11048
rect 7206 10995 7262 10996
rect 7288 10995 7344 10996
rect 7370 11048 7426 11051
rect 7370 10996 7422 11048
rect 7422 10996 7426 11048
rect 7370 10995 7426 10996
rect 7452 11048 7508 11051
rect 7452 10996 7453 11048
rect 7453 10996 7505 11048
rect 7505 10996 7508 11048
rect 7452 10995 7508 10996
rect 7534 11048 7590 11051
rect 7534 10996 7536 11048
rect 7536 10996 7588 11048
rect 7588 10996 7590 11048
rect 7534 10995 7590 10996
rect 7616 11048 7672 11051
rect 7616 10996 7619 11048
rect 7619 10996 7671 11048
rect 7671 10996 7672 11048
rect 7616 10995 7672 10996
rect 7698 11048 7754 11051
rect 7698 10996 7701 11048
rect 7701 10996 7753 11048
rect 7753 10996 7754 11048
rect 7698 10995 7754 10996
rect 7780 11048 7836 11051
rect 7780 10996 7783 11048
rect 7783 10996 7835 11048
rect 7835 10996 7836 11048
rect 7780 10995 7836 10996
rect 7862 11048 7918 11051
rect 7862 10996 7865 11048
rect 7865 10996 7917 11048
rect 7917 10996 7918 11048
rect 7862 10995 7918 10996
rect 7944 11048 8000 11051
rect 7944 10996 7947 11048
rect 7947 10996 7999 11048
rect 7999 10996 8000 11048
rect 7944 10995 8000 10996
rect 8025 11048 8081 11051
rect 8025 10996 8029 11048
rect 8029 10996 8081 11048
rect 8025 10995 8081 10996
rect 8106 11048 8162 11051
rect 8187 11048 8243 11051
rect 8106 10996 8111 11048
rect 8111 10996 8162 11048
rect 8187 10996 8193 11048
rect 8193 10996 8243 11048
rect 8106 10995 8162 10996
rect 8187 10995 8243 10996
rect 368 5144 504 5182
rect 368 4966 382 5144
rect 382 4966 498 5144
rect 498 4966 504 5144
rect 364 2743 420 2799
rect 448 2743 504 2799
rect 364 2652 420 2708
rect 448 2652 504 2708
rect 364 2560 420 2616
rect 448 2560 504 2616
rect 149 2362 205 2418
rect 233 2362 289 2418
rect 149 2271 205 2327
rect 233 2271 289 2327
rect 149 2179 205 2235
rect 233 2179 289 2235
rect 2587 -2418 2643 -2362
rect 2587 -2498 2643 -2442
<< metal3 >>
rect 365 20197 511 20202
rect 365 20061 370 20197
rect 506 20061 511 20197
rect 365 20056 511 20061
tri 365 20053 368 20056 ne
rect 368 20055 511 20056
rect 144 20037 294 20042
rect 144 19901 152 20037
rect 288 19901 294 20037
rect 144 2418 294 19901
tri 363 5187 368 5192 se
rect 368 5187 509 20055
tri 509 20053 511 20055 nw
rect 2406 18083 2472 18092
rect 2406 18027 2411 18083
rect 2467 18027 2472 18083
rect 2406 18003 2472 18027
rect 2406 17947 2411 18003
rect 2467 17947 2472 18003
tri 2373 17838 2406 17871 se
rect 2406 17838 2472 17947
rect 2373 17826 2472 17838
rect 2373 8511 2439 17826
tri 2439 17793 2472 17826 nw
rect 2499 12002 2739 12007
rect 2499 11979 2540 12002
rect 2596 11979 2661 12002
rect 2717 11979 2739 12002
rect 2499 11915 2505 11979
rect 2651 11946 2661 11979
rect 2569 11922 2587 11946
rect 2651 11922 2669 11946
rect 2651 11915 2661 11922
rect 2733 11915 2739 11979
rect 2499 11869 2540 11915
rect 2596 11869 2661 11915
rect 2717 11869 2739 11915
rect 2499 11805 2505 11869
rect 2651 11866 2661 11869
rect 2569 11842 2587 11866
rect 2651 11842 2669 11866
rect 2651 11805 2661 11842
rect 2733 11805 2739 11869
rect 2499 11786 2540 11805
rect 2596 11786 2661 11805
rect 2717 11786 2739 11805
rect 2499 11781 2739 11786
rect 7196 11051 8252 11056
rect 7196 10995 7206 11051
rect 7262 10995 7288 11051
rect 7344 10995 7370 11051
rect 7426 10995 7452 11051
rect 7508 10995 7534 11051
rect 7590 10995 7616 11051
rect 7672 10995 7698 11051
rect 7754 10995 7780 11051
rect 7836 10995 7862 11051
rect 7918 10995 7944 11051
rect 8000 10995 8025 11051
rect 8081 10995 8106 11051
rect 8162 10995 8187 11051
rect 8243 10995 8252 11051
rect 7196 9226 8252 10995
tri 8252 9226 8566 9540 sw
tri 2373 8452 2432 8511 ne
rect 2432 8452 2439 8511
tri 2439 8452 2540 8553 sw
tri 2432 8445 2439 8452 ne
rect 2439 8445 2540 8452
tri 2439 8344 2540 8445 ne
tri 2540 8344 2648 8452 sw
tri 2540 8302 2582 8344 ne
rect 363 5182 509 5187
rect 363 4966 368 5182
rect 504 4966 509 5182
rect 363 4960 509 4966
tri 363 4955 368 4960 ne
tri 359 2808 368 2817 se
rect 368 2808 509 4960
rect 359 2799 509 2808
rect 359 2743 364 2799
rect 420 2743 448 2799
rect 504 2743 509 2799
rect 359 2708 509 2743
rect 359 2652 364 2708
rect 420 2652 448 2708
rect 504 2652 509 2708
rect 359 2616 509 2652
rect 359 2560 364 2616
rect 420 2560 448 2616
rect 504 2560 509 2616
rect 359 2551 509 2560
rect 144 2362 149 2418
rect 205 2362 233 2418
rect 289 2362 294 2418
rect 144 2327 294 2362
rect 144 2271 149 2327
rect 205 2271 233 2327
rect 289 2271 294 2327
rect 144 2235 294 2271
rect 144 2179 149 2235
rect 205 2179 233 2235
rect 289 2179 294 2235
rect 144 2170 294 2179
rect 2582 -2362 2648 8344
rect 2582 -2418 2587 -2362
rect 2643 -2418 2648 -2362
rect 2582 -2442 2648 -2418
rect 2582 -2498 2587 -2442
rect 2643 -2498 2648 -2442
rect 2582 -2507 2648 -2498
<< via3 >>
rect 2505 11946 2540 11979
rect 2540 11946 2569 11979
rect 2587 11946 2596 11979
rect 2596 11946 2651 11979
rect 2669 11946 2717 11979
rect 2717 11946 2733 11979
rect 2505 11922 2569 11946
rect 2587 11922 2651 11946
rect 2669 11922 2733 11946
rect 2505 11915 2540 11922
rect 2540 11915 2569 11922
rect 2587 11915 2596 11922
rect 2596 11915 2651 11922
rect 2669 11915 2717 11922
rect 2717 11915 2733 11922
rect 2505 11866 2540 11869
rect 2540 11866 2569 11869
rect 2587 11866 2596 11869
rect 2596 11866 2651 11869
rect 2669 11866 2717 11869
rect 2717 11866 2733 11869
rect 2505 11842 2569 11866
rect 2587 11842 2651 11866
rect 2669 11842 2733 11866
rect 2505 11805 2540 11842
rect 2540 11805 2569 11842
rect 2587 11805 2596 11842
rect 2596 11805 2651 11842
rect 2669 11805 2717 11842
rect 2717 11805 2733 11842
<< metal4 >>
tri 4007 25022 4385 25400 se
rect 2307 22622 4385 25022
rect 5267 20954 16876 21494
tri 3161 11980 3329 12148 se
rect 3329 11980 3866 12148
rect 2504 11979 3866 11980
rect 2504 11915 2505 11979
rect 2569 11915 2587 11979
rect 2651 11915 2669 11979
rect 2733 11915 3866 11979
rect 2504 11869 3866 11915
rect 2504 11805 2505 11869
rect 2569 11805 2587 11869
rect 2651 11805 2669 11869
rect 2733 11805 3866 11869
rect 2504 11804 3866 11805
tri 3185 11663 3326 11804 ne
rect 3326 9720 3866 11804
tri 3866 9720 4090 9944 sw
tri 17642 9720 17866 9944 se
rect 17866 9720 18406 9986
tri 3326 9718 3328 9720 ne
rect 3328 9718 4090 9720
tri 4090 9718 4092 9720 sw
tri 17640 9718 17642 9720 se
rect 17642 9718 18406 9720
tri 3328 9180 3866 9718 ne
rect 3866 9349 4092 9718
tri 4092 9349 4461 9718 sw
tri 17271 9349 17640 9718 se
rect 17640 9349 18406 9718
tri 18406 9349 18777 9720 sw
rect 3866 9180 4461 9349
tri 3866 8954 4092 9180 ne
rect 4092 8954 4461 9180
tri 4461 8954 4856 9349 sw
tri 16876 8954 17271 9349 se
rect 17271 8954 22978 9349
tri 4092 8414 4632 8954 ne
rect 4632 8414 22978 8954
use sky130_fd_io__gpio_ovtv2_pddrvr_sub  sky130_fd_io__gpio_ovtv2_pddrvr_sub_0
timestamp 1666199351
transform 1 0 414 0 1 -13002
box 380 12107 23743 39298
use sky130_fd_io__gpio_ovtv2_pudrvr_sub  sky130_fd_io__gpio_ovtv2_pudrvr_sub_0
timestamp 1666199351
transform 1 0 0 0 1 0
box 144 -1579 28211 25028
use sky130_fd_io__gpio_ovtv2_res_weak  sky130_fd_io__gpio_ovtv2_res_weak_0
timestamp 1666199351
transform 1 0 -126 0 1 -363
box 263 1014 681 10278
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_0
timestamp 1666199351
transform 1 0 2081 0 1 10971
box 0 0 882 404
use sky130_fd_io__tk_em1s_cdns_5595914180852  sky130_fd_io__tk_em1s_cdns_5595914180852_0
timestamp 1666199351
transform 0 1 748 -1 0 2819
box 0 0 1 1
use sky130_fd_pr__res_generic_po__example_5595914180853  sky130_fd_pr__res_generic_po__example_5595914180853_0
timestamp 1666199351
transform 0 -1 1121 -1 0 2896
box 15 31 585 32
use sky130_fd_pr__res_generic_po__example_5595914180855  sky130_fd_pr__res_generic_po__example_5595914180855_0
timestamp 1666199351
transform 0 -1 1121 -1 0 2194
box 15 31 985 32
use sky130_fd_pr__res_generic_po__example_5595914180856  sky130_fd_pr__res_generic_po__example_5595914180856_0
timestamp 1666199351
transform 0 -1 1121 -1 0 3398
box 15 31 385 32
use sky130_fd_pr__via_l1m1__example_5595914180832  sky130_fd_pr__via_l1m1__example_5595914180832_0
timestamp 1666199351
transform 0 -1 1075 1 0 1091
box 0 0 1 1
use sky130_fd_pr__via_pol1_centered__example_559591418080  sky130_fd_pr__via_pol1_centered__example_559591418080_0
timestamp 1666199351
transform -1 0 921 0 1 1143
box 0 0 1 1
use sky130_fd_pr__via_pol1_centered__example_559591418080  sky130_fd_pr__via_pol1_centered__example_559591418080_1
timestamp 1666199351
transform -1 0 921 0 -1 3449
box 0 0 1 1
<< labels >>
flabel metal2 s 3951 5695 4002 5740 3 FreeSans 200 0 0 0 PUG_H[2]
port 1 nsew
flabel metal2 s 3092 7071 3139 7121 3 FreeSans 200 0 0 0 PU_H_N[3]
port 2 nsew
flabel metal2 s 2815 6972 2863 7022 3 FreeSans 200 0 0 0 PU_H_N[2]
port 3 nsew
flabel metal2 s 2905 7979 2957 8017 3 FreeSans 200 0 0 0 PU_H_N[1]
port 4 nsew
flabel metal2 s 2813 7932 2865 7966 3 FreeSans 200 0 0 0 PU_H_N[0]
port 5 nsew
flabel metal2 s 2537 6045 2589 6123 3 FreeSans 200 0 0 0 PU_CSD_H
port 6 nsew
flabel metal2 s 3674 7709 3753 7759 3 FreeSans 200 0 0 0 PGHS_H
port 7 nsew
flabel metal2 s 18320 20353 18405 20431 3 FreeSans 200 0 0 0 PD_H[3]
port 8 nsew
flabel metal2 s 18322 21020 18391 21072 3 FreeSans 200 0 0 0 PD_H[2]
port 9 nsew
flabel metal2 s 18324 21411 18392 21451 3 FreeSans 200 0 0 0 PD_H[1]
port 10 nsew
flabel metal2 s 18324 21491 18391 21543 3 FreeSans 200 0 0 0 PD_H[0]
port 11 nsew
flabel metal2 s 4132 20500 4184 20578 3 FreeSans 200 0 0 0 PD_CSD_H
port 12 nsew
flabel comment s 26465 8104 26465 8104 0 FreeSans 200 0 0 0 VCC_IO_SOFT
flabel comment s 428 19861 428 19861 0 FreeSans 400 90 0 0 WEAK
flabel comment s 209 19861 209 19861 0 FreeSans 400 90 0 0 SLOW
flabel comment s 229 2527 229 2527 0 FreeSans 400 90 0 0 SLOW
flabel metal1 s 2384 2271 2528 2439 3 FreeSans 200 0 0 0 VPB_DRVR
port 13 nsew
flabel metal1 s 10742 5629 10937 5723 3 FreeSans 200 0 0 0 VDDIO_AMX
port 14 nsew
flabel metal1 s 18589 20683 18620 20750 3 FreeSans 200 90 0 0 TIE_LO_ESD
port 15 nsew
flabel metal1 s 25593 9506 25712 9623 3 FreeSans 200 0 0 0 TIE_HI_ESD
port 16 nsew
flabel metal1 s 3629 4839 3739 4967 3 FreeSans 200 0 0 0 PUG_H[4]
port 17 nsew
flabel metal1 s 3667 6447 3717 6497 3 FreeSans 200 0 0 0 PUG_H[3]
port 18 nsew
flabel metal1 s 24021 3550 24066 3596 3 FreeSans 200 0 0 0 PUG_H[1]
port 19 nsew
flabel metal1 s 24718 4674 24764 4720 3 FreeSans 200 0 0 0 PUG_H[0]
port 20 nsew
flabel metal1 s 6438 11647 6540 11736 3 FreeSans 200 0 0 0 VSSIO_AMX
port 21 nsew
flabel metal1 s 3025 12926 3099 13014 3 FreeSans 200 0 0 0 VSSIO
port 22 nsew
flabel metal1 s 1991 1303 2116 1444 3 FreeSans 200 0 0 0 VSSD
port 23 nsew
flabel metal1 s 1538 892 1717 1071 3 FreeSans 200 0 0 0 VDDIO
port 24 nsew
flabel metal1 s 2648 16599 2694 16651 3 FreeSans 200 0 0 0 NGHS_H
port 25 nsew
flabel metal1 s 1605 10206 1660 10593 3 FreeSans 520 180 0 0 PAD_ESD
port 26 nsew
flabel metal1 s 2862 11026 2917 11357 3 FreeSans 520 180 0 0 PAD
port 27 nsew
<< properties >>
string GDS_END 42045062
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 42017882
<< end >>
