magic
tech sky130A
magscale 1 2
timestamp 1666464484
<< pwell >>
rect 10 66 1950 1128
<< mvnmos >>
rect 228 92 328 1102
rect 384 92 484 1102
rect 540 92 640 1102
rect 696 92 796 1102
rect 852 92 952 1102
rect 1008 92 1108 1102
rect 1164 92 1264 1102
rect 1320 92 1420 1102
rect 1476 92 1576 1102
rect 1632 92 1732 1102
<< mvndiff >>
rect 172 1090 228 1102
rect 172 1056 183 1090
rect 217 1056 228 1090
rect 172 1022 228 1056
rect 172 988 183 1022
rect 217 988 228 1022
rect 172 954 228 988
rect 172 920 183 954
rect 217 920 228 954
rect 172 886 228 920
rect 172 852 183 886
rect 217 852 228 886
rect 172 818 228 852
rect 172 784 183 818
rect 217 784 228 818
rect 172 750 228 784
rect 172 716 183 750
rect 217 716 228 750
rect 172 682 228 716
rect 172 648 183 682
rect 217 648 228 682
rect 172 614 228 648
rect 172 580 183 614
rect 217 580 228 614
rect 172 546 228 580
rect 172 512 183 546
rect 217 512 228 546
rect 172 478 228 512
rect 172 444 183 478
rect 217 444 228 478
rect 172 410 228 444
rect 172 376 183 410
rect 217 376 228 410
rect 172 342 228 376
rect 172 308 183 342
rect 217 308 228 342
rect 172 274 228 308
rect 172 240 183 274
rect 217 240 228 274
rect 172 206 228 240
rect 172 172 183 206
rect 217 172 228 206
rect 172 138 228 172
rect 172 104 183 138
rect 217 104 228 138
rect 172 92 228 104
rect 328 1090 384 1102
rect 328 1056 339 1090
rect 373 1056 384 1090
rect 328 1022 384 1056
rect 328 988 339 1022
rect 373 988 384 1022
rect 328 954 384 988
rect 328 920 339 954
rect 373 920 384 954
rect 328 886 384 920
rect 328 852 339 886
rect 373 852 384 886
rect 328 818 384 852
rect 328 784 339 818
rect 373 784 384 818
rect 328 750 384 784
rect 328 716 339 750
rect 373 716 384 750
rect 328 682 384 716
rect 328 648 339 682
rect 373 648 384 682
rect 328 614 384 648
rect 328 580 339 614
rect 373 580 384 614
rect 328 546 384 580
rect 328 512 339 546
rect 373 512 384 546
rect 328 478 384 512
rect 328 444 339 478
rect 373 444 384 478
rect 328 410 384 444
rect 328 376 339 410
rect 373 376 384 410
rect 328 342 384 376
rect 328 308 339 342
rect 373 308 384 342
rect 328 274 384 308
rect 328 240 339 274
rect 373 240 384 274
rect 328 206 384 240
rect 328 172 339 206
rect 373 172 384 206
rect 328 138 384 172
rect 328 104 339 138
rect 373 104 384 138
rect 328 92 384 104
rect 484 1090 540 1102
rect 484 1056 495 1090
rect 529 1056 540 1090
rect 484 1022 540 1056
rect 484 988 495 1022
rect 529 988 540 1022
rect 484 954 540 988
rect 484 920 495 954
rect 529 920 540 954
rect 484 886 540 920
rect 484 852 495 886
rect 529 852 540 886
rect 484 818 540 852
rect 484 784 495 818
rect 529 784 540 818
rect 484 750 540 784
rect 484 716 495 750
rect 529 716 540 750
rect 484 682 540 716
rect 484 648 495 682
rect 529 648 540 682
rect 484 614 540 648
rect 484 580 495 614
rect 529 580 540 614
rect 484 546 540 580
rect 484 512 495 546
rect 529 512 540 546
rect 484 478 540 512
rect 484 444 495 478
rect 529 444 540 478
rect 484 410 540 444
rect 484 376 495 410
rect 529 376 540 410
rect 484 342 540 376
rect 484 308 495 342
rect 529 308 540 342
rect 484 274 540 308
rect 484 240 495 274
rect 529 240 540 274
rect 484 206 540 240
rect 484 172 495 206
rect 529 172 540 206
rect 484 138 540 172
rect 484 104 495 138
rect 529 104 540 138
rect 484 92 540 104
rect 640 1090 696 1102
rect 640 1056 651 1090
rect 685 1056 696 1090
rect 640 1022 696 1056
rect 640 988 651 1022
rect 685 988 696 1022
rect 640 954 696 988
rect 640 920 651 954
rect 685 920 696 954
rect 640 886 696 920
rect 640 852 651 886
rect 685 852 696 886
rect 640 818 696 852
rect 640 784 651 818
rect 685 784 696 818
rect 640 750 696 784
rect 640 716 651 750
rect 685 716 696 750
rect 640 682 696 716
rect 640 648 651 682
rect 685 648 696 682
rect 640 614 696 648
rect 640 580 651 614
rect 685 580 696 614
rect 640 546 696 580
rect 640 512 651 546
rect 685 512 696 546
rect 640 478 696 512
rect 640 444 651 478
rect 685 444 696 478
rect 640 410 696 444
rect 640 376 651 410
rect 685 376 696 410
rect 640 342 696 376
rect 640 308 651 342
rect 685 308 696 342
rect 640 274 696 308
rect 640 240 651 274
rect 685 240 696 274
rect 640 206 696 240
rect 640 172 651 206
rect 685 172 696 206
rect 640 138 696 172
rect 640 104 651 138
rect 685 104 696 138
rect 640 92 696 104
rect 796 1090 852 1102
rect 796 1056 807 1090
rect 841 1056 852 1090
rect 796 1022 852 1056
rect 796 988 807 1022
rect 841 988 852 1022
rect 796 954 852 988
rect 796 920 807 954
rect 841 920 852 954
rect 796 886 852 920
rect 796 852 807 886
rect 841 852 852 886
rect 796 818 852 852
rect 796 784 807 818
rect 841 784 852 818
rect 796 750 852 784
rect 796 716 807 750
rect 841 716 852 750
rect 796 682 852 716
rect 796 648 807 682
rect 841 648 852 682
rect 796 614 852 648
rect 796 580 807 614
rect 841 580 852 614
rect 796 546 852 580
rect 796 512 807 546
rect 841 512 852 546
rect 796 478 852 512
rect 796 444 807 478
rect 841 444 852 478
rect 796 410 852 444
rect 796 376 807 410
rect 841 376 852 410
rect 796 342 852 376
rect 796 308 807 342
rect 841 308 852 342
rect 796 274 852 308
rect 796 240 807 274
rect 841 240 852 274
rect 796 206 852 240
rect 796 172 807 206
rect 841 172 852 206
rect 796 138 852 172
rect 796 104 807 138
rect 841 104 852 138
rect 796 92 852 104
rect 952 1090 1008 1102
rect 952 1056 963 1090
rect 997 1056 1008 1090
rect 952 1022 1008 1056
rect 952 988 963 1022
rect 997 988 1008 1022
rect 952 954 1008 988
rect 952 920 963 954
rect 997 920 1008 954
rect 952 886 1008 920
rect 952 852 963 886
rect 997 852 1008 886
rect 952 818 1008 852
rect 952 784 963 818
rect 997 784 1008 818
rect 952 750 1008 784
rect 952 716 963 750
rect 997 716 1008 750
rect 952 682 1008 716
rect 952 648 963 682
rect 997 648 1008 682
rect 952 614 1008 648
rect 952 580 963 614
rect 997 580 1008 614
rect 952 546 1008 580
rect 952 512 963 546
rect 997 512 1008 546
rect 952 478 1008 512
rect 952 444 963 478
rect 997 444 1008 478
rect 952 410 1008 444
rect 952 376 963 410
rect 997 376 1008 410
rect 952 342 1008 376
rect 952 308 963 342
rect 997 308 1008 342
rect 952 274 1008 308
rect 952 240 963 274
rect 997 240 1008 274
rect 952 206 1008 240
rect 952 172 963 206
rect 997 172 1008 206
rect 952 138 1008 172
rect 952 104 963 138
rect 997 104 1008 138
rect 952 92 1008 104
rect 1108 1090 1164 1102
rect 1108 1056 1119 1090
rect 1153 1056 1164 1090
rect 1108 1022 1164 1056
rect 1108 988 1119 1022
rect 1153 988 1164 1022
rect 1108 954 1164 988
rect 1108 920 1119 954
rect 1153 920 1164 954
rect 1108 886 1164 920
rect 1108 852 1119 886
rect 1153 852 1164 886
rect 1108 818 1164 852
rect 1108 784 1119 818
rect 1153 784 1164 818
rect 1108 750 1164 784
rect 1108 716 1119 750
rect 1153 716 1164 750
rect 1108 682 1164 716
rect 1108 648 1119 682
rect 1153 648 1164 682
rect 1108 614 1164 648
rect 1108 580 1119 614
rect 1153 580 1164 614
rect 1108 546 1164 580
rect 1108 512 1119 546
rect 1153 512 1164 546
rect 1108 478 1164 512
rect 1108 444 1119 478
rect 1153 444 1164 478
rect 1108 410 1164 444
rect 1108 376 1119 410
rect 1153 376 1164 410
rect 1108 342 1164 376
rect 1108 308 1119 342
rect 1153 308 1164 342
rect 1108 274 1164 308
rect 1108 240 1119 274
rect 1153 240 1164 274
rect 1108 206 1164 240
rect 1108 172 1119 206
rect 1153 172 1164 206
rect 1108 138 1164 172
rect 1108 104 1119 138
rect 1153 104 1164 138
rect 1108 92 1164 104
rect 1264 1090 1320 1102
rect 1264 1056 1275 1090
rect 1309 1056 1320 1090
rect 1264 1022 1320 1056
rect 1264 988 1275 1022
rect 1309 988 1320 1022
rect 1264 954 1320 988
rect 1264 920 1275 954
rect 1309 920 1320 954
rect 1264 886 1320 920
rect 1264 852 1275 886
rect 1309 852 1320 886
rect 1264 818 1320 852
rect 1264 784 1275 818
rect 1309 784 1320 818
rect 1264 750 1320 784
rect 1264 716 1275 750
rect 1309 716 1320 750
rect 1264 682 1320 716
rect 1264 648 1275 682
rect 1309 648 1320 682
rect 1264 614 1320 648
rect 1264 580 1275 614
rect 1309 580 1320 614
rect 1264 546 1320 580
rect 1264 512 1275 546
rect 1309 512 1320 546
rect 1264 478 1320 512
rect 1264 444 1275 478
rect 1309 444 1320 478
rect 1264 410 1320 444
rect 1264 376 1275 410
rect 1309 376 1320 410
rect 1264 342 1320 376
rect 1264 308 1275 342
rect 1309 308 1320 342
rect 1264 274 1320 308
rect 1264 240 1275 274
rect 1309 240 1320 274
rect 1264 206 1320 240
rect 1264 172 1275 206
rect 1309 172 1320 206
rect 1264 138 1320 172
rect 1264 104 1275 138
rect 1309 104 1320 138
rect 1264 92 1320 104
rect 1420 1090 1476 1102
rect 1420 1056 1431 1090
rect 1465 1056 1476 1090
rect 1420 1022 1476 1056
rect 1420 988 1431 1022
rect 1465 988 1476 1022
rect 1420 954 1476 988
rect 1420 920 1431 954
rect 1465 920 1476 954
rect 1420 886 1476 920
rect 1420 852 1431 886
rect 1465 852 1476 886
rect 1420 818 1476 852
rect 1420 784 1431 818
rect 1465 784 1476 818
rect 1420 750 1476 784
rect 1420 716 1431 750
rect 1465 716 1476 750
rect 1420 682 1476 716
rect 1420 648 1431 682
rect 1465 648 1476 682
rect 1420 614 1476 648
rect 1420 580 1431 614
rect 1465 580 1476 614
rect 1420 546 1476 580
rect 1420 512 1431 546
rect 1465 512 1476 546
rect 1420 478 1476 512
rect 1420 444 1431 478
rect 1465 444 1476 478
rect 1420 410 1476 444
rect 1420 376 1431 410
rect 1465 376 1476 410
rect 1420 342 1476 376
rect 1420 308 1431 342
rect 1465 308 1476 342
rect 1420 274 1476 308
rect 1420 240 1431 274
rect 1465 240 1476 274
rect 1420 206 1476 240
rect 1420 172 1431 206
rect 1465 172 1476 206
rect 1420 138 1476 172
rect 1420 104 1431 138
rect 1465 104 1476 138
rect 1420 92 1476 104
rect 1576 1090 1632 1102
rect 1576 1056 1587 1090
rect 1621 1056 1632 1090
rect 1576 1022 1632 1056
rect 1576 988 1587 1022
rect 1621 988 1632 1022
rect 1576 954 1632 988
rect 1576 920 1587 954
rect 1621 920 1632 954
rect 1576 886 1632 920
rect 1576 852 1587 886
rect 1621 852 1632 886
rect 1576 818 1632 852
rect 1576 784 1587 818
rect 1621 784 1632 818
rect 1576 750 1632 784
rect 1576 716 1587 750
rect 1621 716 1632 750
rect 1576 682 1632 716
rect 1576 648 1587 682
rect 1621 648 1632 682
rect 1576 614 1632 648
rect 1576 580 1587 614
rect 1621 580 1632 614
rect 1576 546 1632 580
rect 1576 512 1587 546
rect 1621 512 1632 546
rect 1576 478 1632 512
rect 1576 444 1587 478
rect 1621 444 1632 478
rect 1576 410 1632 444
rect 1576 376 1587 410
rect 1621 376 1632 410
rect 1576 342 1632 376
rect 1576 308 1587 342
rect 1621 308 1632 342
rect 1576 274 1632 308
rect 1576 240 1587 274
rect 1621 240 1632 274
rect 1576 206 1632 240
rect 1576 172 1587 206
rect 1621 172 1632 206
rect 1576 138 1632 172
rect 1576 104 1587 138
rect 1621 104 1632 138
rect 1576 92 1632 104
rect 1732 1090 1788 1102
rect 1732 1056 1743 1090
rect 1777 1056 1788 1090
rect 1732 1022 1788 1056
rect 1732 988 1743 1022
rect 1777 988 1788 1022
rect 1732 954 1788 988
rect 1732 920 1743 954
rect 1777 920 1788 954
rect 1732 886 1788 920
rect 1732 852 1743 886
rect 1777 852 1788 886
rect 1732 818 1788 852
rect 1732 784 1743 818
rect 1777 784 1788 818
rect 1732 750 1788 784
rect 1732 716 1743 750
rect 1777 716 1788 750
rect 1732 682 1788 716
rect 1732 648 1743 682
rect 1777 648 1788 682
rect 1732 614 1788 648
rect 1732 580 1743 614
rect 1777 580 1788 614
rect 1732 546 1788 580
rect 1732 512 1743 546
rect 1777 512 1788 546
rect 1732 478 1788 512
rect 1732 444 1743 478
rect 1777 444 1788 478
rect 1732 410 1788 444
rect 1732 376 1743 410
rect 1777 376 1788 410
rect 1732 342 1788 376
rect 1732 308 1743 342
rect 1777 308 1788 342
rect 1732 274 1788 308
rect 1732 240 1743 274
rect 1777 240 1788 274
rect 1732 206 1788 240
rect 1732 172 1743 206
rect 1777 172 1788 206
rect 1732 138 1788 172
rect 1732 104 1743 138
rect 1777 104 1788 138
rect 1732 92 1788 104
<< mvndiffc >>
rect 183 1056 217 1090
rect 183 988 217 1022
rect 183 920 217 954
rect 183 852 217 886
rect 183 784 217 818
rect 183 716 217 750
rect 183 648 217 682
rect 183 580 217 614
rect 183 512 217 546
rect 183 444 217 478
rect 183 376 217 410
rect 183 308 217 342
rect 183 240 217 274
rect 183 172 217 206
rect 183 104 217 138
rect 339 1056 373 1090
rect 339 988 373 1022
rect 339 920 373 954
rect 339 852 373 886
rect 339 784 373 818
rect 339 716 373 750
rect 339 648 373 682
rect 339 580 373 614
rect 339 512 373 546
rect 339 444 373 478
rect 339 376 373 410
rect 339 308 373 342
rect 339 240 373 274
rect 339 172 373 206
rect 339 104 373 138
rect 495 1056 529 1090
rect 495 988 529 1022
rect 495 920 529 954
rect 495 852 529 886
rect 495 784 529 818
rect 495 716 529 750
rect 495 648 529 682
rect 495 580 529 614
rect 495 512 529 546
rect 495 444 529 478
rect 495 376 529 410
rect 495 308 529 342
rect 495 240 529 274
rect 495 172 529 206
rect 495 104 529 138
rect 651 1056 685 1090
rect 651 988 685 1022
rect 651 920 685 954
rect 651 852 685 886
rect 651 784 685 818
rect 651 716 685 750
rect 651 648 685 682
rect 651 580 685 614
rect 651 512 685 546
rect 651 444 685 478
rect 651 376 685 410
rect 651 308 685 342
rect 651 240 685 274
rect 651 172 685 206
rect 651 104 685 138
rect 807 1056 841 1090
rect 807 988 841 1022
rect 807 920 841 954
rect 807 852 841 886
rect 807 784 841 818
rect 807 716 841 750
rect 807 648 841 682
rect 807 580 841 614
rect 807 512 841 546
rect 807 444 841 478
rect 807 376 841 410
rect 807 308 841 342
rect 807 240 841 274
rect 807 172 841 206
rect 807 104 841 138
rect 963 1056 997 1090
rect 963 988 997 1022
rect 963 920 997 954
rect 963 852 997 886
rect 963 784 997 818
rect 963 716 997 750
rect 963 648 997 682
rect 963 580 997 614
rect 963 512 997 546
rect 963 444 997 478
rect 963 376 997 410
rect 963 308 997 342
rect 963 240 997 274
rect 963 172 997 206
rect 963 104 997 138
rect 1119 1056 1153 1090
rect 1119 988 1153 1022
rect 1119 920 1153 954
rect 1119 852 1153 886
rect 1119 784 1153 818
rect 1119 716 1153 750
rect 1119 648 1153 682
rect 1119 580 1153 614
rect 1119 512 1153 546
rect 1119 444 1153 478
rect 1119 376 1153 410
rect 1119 308 1153 342
rect 1119 240 1153 274
rect 1119 172 1153 206
rect 1119 104 1153 138
rect 1275 1056 1309 1090
rect 1275 988 1309 1022
rect 1275 920 1309 954
rect 1275 852 1309 886
rect 1275 784 1309 818
rect 1275 716 1309 750
rect 1275 648 1309 682
rect 1275 580 1309 614
rect 1275 512 1309 546
rect 1275 444 1309 478
rect 1275 376 1309 410
rect 1275 308 1309 342
rect 1275 240 1309 274
rect 1275 172 1309 206
rect 1275 104 1309 138
rect 1431 1056 1465 1090
rect 1431 988 1465 1022
rect 1431 920 1465 954
rect 1431 852 1465 886
rect 1431 784 1465 818
rect 1431 716 1465 750
rect 1431 648 1465 682
rect 1431 580 1465 614
rect 1431 512 1465 546
rect 1431 444 1465 478
rect 1431 376 1465 410
rect 1431 308 1465 342
rect 1431 240 1465 274
rect 1431 172 1465 206
rect 1431 104 1465 138
rect 1587 1056 1621 1090
rect 1587 988 1621 1022
rect 1587 920 1621 954
rect 1587 852 1621 886
rect 1587 784 1621 818
rect 1587 716 1621 750
rect 1587 648 1621 682
rect 1587 580 1621 614
rect 1587 512 1621 546
rect 1587 444 1621 478
rect 1587 376 1621 410
rect 1587 308 1621 342
rect 1587 240 1621 274
rect 1587 172 1621 206
rect 1587 104 1621 138
rect 1743 1056 1777 1090
rect 1743 988 1777 1022
rect 1743 920 1777 954
rect 1743 852 1777 886
rect 1743 784 1777 818
rect 1743 716 1777 750
rect 1743 648 1777 682
rect 1743 580 1777 614
rect 1743 512 1777 546
rect 1743 444 1777 478
rect 1743 376 1777 410
rect 1743 308 1777 342
rect 1743 240 1777 274
rect 1743 172 1777 206
rect 1743 104 1777 138
<< mvpsubdiff >>
rect 36 1056 94 1102
rect 36 1022 48 1056
rect 82 1022 94 1056
rect 36 988 94 1022
rect 36 954 48 988
rect 82 954 94 988
rect 36 920 94 954
rect 36 886 48 920
rect 82 886 94 920
rect 36 852 94 886
rect 36 818 48 852
rect 82 818 94 852
rect 36 784 94 818
rect 36 750 48 784
rect 82 750 94 784
rect 36 716 94 750
rect 36 682 48 716
rect 82 682 94 716
rect 36 648 94 682
rect 36 614 48 648
rect 82 614 94 648
rect 36 580 94 614
rect 36 546 48 580
rect 82 546 94 580
rect 36 512 94 546
rect 36 478 48 512
rect 82 478 94 512
rect 36 444 94 478
rect 36 410 48 444
rect 82 410 94 444
rect 36 376 94 410
rect 36 342 48 376
rect 82 342 94 376
rect 36 308 94 342
rect 36 274 48 308
rect 82 274 94 308
rect 36 240 94 274
rect 36 206 48 240
rect 82 206 94 240
rect 36 172 94 206
rect 36 138 48 172
rect 82 138 94 172
rect 36 92 94 138
rect 1866 1056 1924 1102
rect 1866 1022 1878 1056
rect 1912 1022 1924 1056
rect 1866 988 1924 1022
rect 1866 954 1878 988
rect 1912 954 1924 988
rect 1866 920 1924 954
rect 1866 886 1878 920
rect 1912 886 1924 920
rect 1866 852 1924 886
rect 1866 818 1878 852
rect 1912 818 1924 852
rect 1866 784 1924 818
rect 1866 750 1878 784
rect 1912 750 1924 784
rect 1866 716 1924 750
rect 1866 682 1878 716
rect 1912 682 1924 716
rect 1866 648 1924 682
rect 1866 614 1878 648
rect 1912 614 1924 648
rect 1866 580 1924 614
rect 1866 546 1878 580
rect 1912 546 1924 580
rect 1866 512 1924 546
rect 1866 478 1878 512
rect 1912 478 1924 512
rect 1866 444 1924 478
rect 1866 410 1878 444
rect 1912 410 1924 444
rect 1866 376 1924 410
rect 1866 342 1878 376
rect 1912 342 1924 376
rect 1866 308 1924 342
rect 1866 274 1878 308
rect 1912 274 1924 308
rect 1866 240 1924 274
rect 1866 206 1878 240
rect 1912 206 1924 240
rect 1866 172 1924 206
rect 1866 138 1878 172
rect 1912 138 1924 172
rect 1866 92 1924 138
<< mvpsubdiffcont >>
rect 48 1022 82 1056
rect 48 954 82 988
rect 48 886 82 920
rect 48 818 82 852
rect 48 750 82 784
rect 48 682 82 716
rect 48 614 82 648
rect 48 546 82 580
rect 48 478 82 512
rect 48 410 82 444
rect 48 342 82 376
rect 48 274 82 308
rect 48 206 82 240
rect 48 138 82 172
rect 1878 1022 1912 1056
rect 1878 954 1912 988
rect 1878 886 1912 920
rect 1878 818 1912 852
rect 1878 750 1912 784
rect 1878 682 1912 716
rect 1878 614 1912 648
rect 1878 546 1912 580
rect 1878 478 1912 512
rect 1878 410 1912 444
rect 1878 342 1912 376
rect 1878 274 1912 308
rect 1878 206 1912 240
rect 1878 138 1912 172
<< poly >>
rect 199 1174 1761 1194
rect 199 1140 215 1174
rect 249 1140 283 1174
rect 317 1140 351 1174
rect 385 1140 419 1174
rect 453 1140 487 1174
rect 521 1140 555 1174
rect 589 1140 623 1174
rect 657 1140 691 1174
rect 725 1140 759 1174
rect 793 1140 827 1174
rect 861 1140 895 1174
rect 929 1140 963 1174
rect 997 1140 1031 1174
rect 1065 1140 1099 1174
rect 1133 1140 1167 1174
rect 1201 1140 1235 1174
rect 1269 1140 1303 1174
rect 1337 1140 1371 1174
rect 1405 1140 1439 1174
rect 1473 1140 1507 1174
rect 1541 1140 1575 1174
rect 1609 1140 1643 1174
rect 1677 1140 1711 1174
rect 1745 1140 1761 1174
rect 199 1124 1761 1140
rect 228 1102 328 1124
rect 384 1102 484 1124
rect 540 1102 640 1124
rect 696 1102 796 1124
rect 852 1102 952 1124
rect 1008 1102 1108 1124
rect 1164 1102 1264 1124
rect 1320 1102 1420 1124
rect 1476 1102 1576 1124
rect 1632 1102 1732 1124
rect 228 70 328 92
rect 384 70 484 92
rect 540 70 640 92
rect 696 70 796 92
rect 852 70 952 92
rect 1008 70 1108 92
rect 1164 70 1264 92
rect 1320 70 1420 92
rect 1476 70 1576 92
rect 1632 70 1732 92
rect 199 54 1761 70
rect 199 20 215 54
rect 249 20 283 54
rect 317 20 351 54
rect 385 20 419 54
rect 453 20 487 54
rect 521 20 555 54
rect 589 20 623 54
rect 657 20 691 54
rect 725 20 759 54
rect 793 20 827 54
rect 861 20 895 54
rect 929 20 963 54
rect 997 20 1031 54
rect 1065 20 1099 54
rect 1133 20 1167 54
rect 1201 20 1235 54
rect 1269 20 1303 54
rect 1337 20 1371 54
rect 1405 20 1439 54
rect 1473 20 1507 54
rect 1541 20 1575 54
rect 1609 20 1643 54
rect 1677 20 1711 54
rect 1745 20 1761 54
rect 199 0 1761 20
<< polycont >>
rect 215 1140 249 1174
rect 283 1140 317 1174
rect 351 1140 385 1174
rect 419 1140 453 1174
rect 487 1140 521 1174
rect 555 1140 589 1174
rect 623 1140 657 1174
rect 691 1140 725 1174
rect 759 1140 793 1174
rect 827 1140 861 1174
rect 895 1140 929 1174
rect 963 1140 997 1174
rect 1031 1140 1065 1174
rect 1099 1140 1133 1174
rect 1167 1140 1201 1174
rect 1235 1140 1269 1174
rect 1303 1140 1337 1174
rect 1371 1140 1405 1174
rect 1439 1140 1473 1174
rect 1507 1140 1541 1174
rect 1575 1140 1609 1174
rect 1643 1140 1677 1174
rect 1711 1140 1745 1174
rect 215 20 249 54
rect 283 20 317 54
rect 351 20 385 54
rect 419 20 453 54
rect 487 20 521 54
rect 555 20 589 54
rect 623 20 657 54
rect 691 20 725 54
rect 759 20 793 54
rect 827 20 861 54
rect 895 20 929 54
rect 963 20 997 54
rect 1031 20 1065 54
rect 1099 20 1133 54
rect 1167 20 1201 54
rect 1235 20 1269 54
rect 1303 20 1337 54
rect 1371 20 1405 54
rect 1439 20 1473 54
rect 1507 20 1541 54
rect 1575 20 1609 54
rect 1643 20 1677 54
rect 1711 20 1745 54
<< locali >>
rect 199 1140 207 1174
rect 249 1140 279 1174
rect 317 1140 351 1174
rect 385 1140 419 1174
rect 457 1140 487 1174
rect 529 1140 555 1174
rect 601 1140 623 1174
rect 673 1140 691 1174
rect 745 1140 759 1174
rect 817 1140 827 1174
rect 889 1140 895 1174
rect 961 1140 963 1174
rect 997 1140 999 1174
rect 1065 1140 1071 1174
rect 1133 1140 1143 1174
rect 1201 1140 1215 1174
rect 1269 1140 1287 1174
rect 1337 1140 1359 1174
rect 1405 1140 1431 1174
rect 1473 1140 1503 1174
rect 1541 1140 1575 1174
rect 1609 1140 1643 1174
rect 1681 1140 1711 1174
rect 1753 1140 1761 1174
rect 183 1090 217 1106
rect 48 1010 82 1022
rect 48 938 82 954
rect 48 866 82 886
rect 48 794 82 818
rect 48 722 82 750
rect 48 650 82 682
rect 48 580 82 614
rect 48 512 82 544
rect 48 444 82 472
rect 48 376 82 400
rect 48 308 82 328
rect 48 240 82 256
rect 48 172 82 184
rect 183 1022 217 1048
rect 183 954 217 976
rect 183 886 217 904
rect 183 818 217 832
rect 183 750 217 760
rect 183 682 217 688
rect 183 614 217 616
rect 183 578 217 580
rect 183 506 217 512
rect 183 434 217 444
rect 183 362 217 376
rect 183 290 217 308
rect 183 218 217 240
rect 183 146 217 172
rect 183 88 217 104
rect 339 1090 373 1106
rect 339 1022 373 1048
rect 339 954 373 976
rect 339 886 373 904
rect 339 818 373 832
rect 339 750 373 760
rect 339 682 373 688
rect 339 614 373 616
rect 339 578 373 580
rect 339 506 373 512
rect 339 434 373 444
rect 339 362 373 376
rect 339 290 373 308
rect 339 218 373 240
rect 339 146 373 172
rect 339 88 373 104
rect 495 1090 529 1106
rect 495 1022 529 1048
rect 495 954 529 976
rect 495 886 529 904
rect 495 818 529 832
rect 495 750 529 760
rect 495 682 529 688
rect 495 614 529 616
rect 495 578 529 580
rect 495 506 529 512
rect 495 434 529 444
rect 495 362 529 376
rect 495 290 529 308
rect 495 218 529 240
rect 495 146 529 172
rect 495 88 529 104
rect 651 1090 685 1106
rect 651 1022 685 1048
rect 651 954 685 976
rect 651 886 685 904
rect 651 818 685 832
rect 651 750 685 760
rect 651 682 685 688
rect 651 614 685 616
rect 651 578 685 580
rect 651 506 685 512
rect 651 434 685 444
rect 651 362 685 376
rect 651 290 685 308
rect 651 218 685 240
rect 651 146 685 172
rect 651 88 685 104
rect 807 1090 841 1106
rect 807 1022 841 1048
rect 807 954 841 976
rect 807 886 841 904
rect 807 818 841 832
rect 807 750 841 760
rect 807 682 841 688
rect 807 614 841 616
rect 807 578 841 580
rect 807 506 841 512
rect 807 434 841 444
rect 807 362 841 376
rect 807 290 841 308
rect 807 218 841 240
rect 807 146 841 172
rect 807 88 841 104
rect 963 1090 997 1106
rect 963 1022 997 1048
rect 963 954 997 976
rect 963 886 997 904
rect 963 818 997 832
rect 963 750 997 760
rect 963 682 997 688
rect 963 614 997 616
rect 963 578 997 580
rect 963 506 997 512
rect 963 434 997 444
rect 963 362 997 376
rect 963 290 997 308
rect 963 218 997 240
rect 963 146 997 172
rect 963 88 997 104
rect 1119 1090 1153 1106
rect 1119 1022 1153 1048
rect 1119 954 1153 976
rect 1119 886 1153 904
rect 1119 818 1153 832
rect 1119 750 1153 760
rect 1119 682 1153 688
rect 1119 614 1153 616
rect 1119 578 1153 580
rect 1119 506 1153 512
rect 1119 434 1153 444
rect 1119 362 1153 376
rect 1119 290 1153 308
rect 1119 218 1153 240
rect 1119 146 1153 172
rect 1119 88 1153 104
rect 1275 1090 1309 1106
rect 1275 1022 1309 1048
rect 1275 954 1309 976
rect 1275 886 1309 904
rect 1275 818 1309 832
rect 1275 750 1309 760
rect 1275 682 1309 688
rect 1275 614 1309 616
rect 1275 578 1309 580
rect 1275 506 1309 512
rect 1275 434 1309 444
rect 1275 362 1309 376
rect 1275 290 1309 308
rect 1275 218 1309 240
rect 1275 146 1309 172
rect 1275 88 1309 104
rect 1431 1090 1465 1106
rect 1431 1022 1465 1048
rect 1431 954 1465 976
rect 1431 886 1465 904
rect 1431 818 1465 832
rect 1431 750 1465 760
rect 1431 682 1465 688
rect 1431 614 1465 616
rect 1431 578 1465 580
rect 1431 506 1465 512
rect 1431 434 1465 444
rect 1431 362 1465 376
rect 1431 290 1465 308
rect 1431 218 1465 240
rect 1431 146 1465 172
rect 1431 88 1465 104
rect 1587 1090 1621 1106
rect 1587 1022 1621 1048
rect 1587 954 1621 976
rect 1587 886 1621 904
rect 1587 818 1621 832
rect 1587 750 1621 760
rect 1587 682 1621 688
rect 1587 614 1621 616
rect 1587 578 1621 580
rect 1587 506 1621 512
rect 1587 434 1621 444
rect 1587 362 1621 376
rect 1587 290 1621 308
rect 1587 218 1621 240
rect 1587 146 1621 172
rect 1587 88 1621 104
rect 1743 1090 1777 1106
rect 1743 1022 1777 1048
rect 1743 954 1777 976
rect 1743 886 1777 904
rect 1743 818 1777 832
rect 1743 750 1777 760
rect 1743 682 1777 688
rect 1743 614 1777 616
rect 1743 578 1777 580
rect 1743 506 1777 512
rect 1743 434 1777 444
rect 1743 362 1777 376
rect 1743 290 1777 308
rect 1743 218 1777 240
rect 1743 146 1777 172
rect 1878 1010 1912 1022
rect 1878 938 1912 954
rect 1878 866 1912 886
rect 1878 794 1912 818
rect 1878 722 1912 750
rect 1878 650 1912 682
rect 1878 580 1912 614
rect 1878 512 1912 544
rect 1878 444 1912 472
rect 1878 376 1912 400
rect 1878 308 1912 328
rect 1878 240 1912 256
rect 1878 172 1912 184
rect 1743 88 1777 104
rect 199 20 207 54
rect 249 20 279 54
rect 317 20 351 54
rect 385 20 419 54
rect 457 20 487 54
rect 529 20 555 54
rect 601 20 623 54
rect 673 20 691 54
rect 745 20 759 54
rect 817 20 827 54
rect 889 20 895 54
rect 961 20 963 54
rect 997 20 999 54
rect 1065 20 1071 54
rect 1133 20 1143 54
rect 1201 20 1215 54
rect 1269 20 1287 54
rect 1337 20 1359 54
rect 1405 20 1431 54
rect 1473 20 1503 54
rect 1541 20 1575 54
rect 1609 20 1643 54
rect 1681 20 1711 54
rect 1753 20 1761 54
<< viali >>
rect 207 1140 215 1174
rect 215 1140 241 1174
rect 279 1140 283 1174
rect 283 1140 313 1174
rect 351 1140 385 1174
rect 423 1140 453 1174
rect 453 1140 457 1174
rect 495 1140 521 1174
rect 521 1140 529 1174
rect 567 1140 589 1174
rect 589 1140 601 1174
rect 639 1140 657 1174
rect 657 1140 673 1174
rect 711 1140 725 1174
rect 725 1140 745 1174
rect 783 1140 793 1174
rect 793 1140 817 1174
rect 855 1140 861 1174
rect 861 1140 889 1174
rect 927 1140 929 1174
rect 929 1140 961 1174
rect 999 1140 1031 1174
rect 1031 1140 1033 1174
rect 1071 1140 1099 1174
rect 1099 1140 1105 1174
rect 1143 1140 1167 1174
rect 1167 1140 1177 1174
rect 1215 1140 1235 1174
rect 1235 1140 1249 1174
rect 1287 1140 1303 1174
rect 1303 1140 1321 1174
rect 1359 1140 1371 1174
rect 1371 1140 1393 1174
rect 1431 1140 1439 1174
rect 1439 1140 1465 1174
rect 1503 1140 1507 1174
rect 1507 1140 1537 1174
rect 1575 1140 1609 1174
rect 1647 1140 1677 1174
rect 1677 1140 1681 1174
rect 1719 1140 1745 1174
rect 1745 1140 1753 1174
rect 48 1056 82 1082
rect 48 1048 82 1056
rect 48 988 82 1010
rect 48 976 82 988
rect 48 920 82 938
rect 48 904 82 920
rect 48 852 82 866
rect 48 832 82 852
rect 48 784 82 794
rect 48 760 82 784
rect 48 716 82 722
rect 48 688 82 716
rect 48 648 82 650
rect 48 616 82 648
rect 48 546 82 578
rect 48 544 82 546
rect 48 478 82 506
rect 48 472 82 478
rect 48 410 82 434
rect 48 400 82 410
rect 48 342 82 362
rect 48 328 82 342
rect 48 274 82 290
rect 48 256 82 274
rect 48 206 82 218
rect 48 184 82 206
rect 48 138 82 146
rect 48 112 82 138
rect 183 1056 217 1082
rect 183 1048 217 1056
rect 183 988 217 1010
rect 183 976 217 988
rect 183 920 217 938
rect 183 904 217 920
rect 183 852 217 866
rect 183 832 217 852
rect 183 784 217 794
rect 183 760 217 784
rect 183 716 217 722
rect 183 688 217 716
rect 183 648 217 650
rect 183 616 217 648
rect 183 546 217 578
rect 183 544 217 546
rect 183 478 217 506
rect 183 472 217 478
rect 183 410 217 434
rect 183 400 217 410
rect 183 342 217 362
rect 183 328 217 342
rect 183 274 217 290
rect 183 256 217 274
rect 183 206 217 218
rect 183 184 217 206
rect 183 138 217 146
rect 183 112 217 138
rect 339 1056 373 1082
rect 339 1048 373 1056
rect 339 988 373 1010
rect 339 976 373 988
rect 339 920 373 938
rect 339 904 373 920
rect 339 852 373 866
rect 339 832 373 852
rect 339 784 373 794
rect 339 760 373 784
rect 339 716 373 722
rect 339 688 373 716
rect 339 648 373 650
rect 339 616 373 648
rect 339 546 373 578
rect 339 544 373 546
rect 339 478 373 506
rect 339 472 373 478
rect 339 410 373 434
rect 339 400 373 410
rect 339 342 373 362
rect 339 328 373 342
rect 339 274 373 290
rect 339 256 373 274
rect 339 206 373 218
rect 339 184 373 206
rect 339 138 373 146
rect 339 112 373 138
rect 495 1056 529 1082
rect 495 1048 529 1056
rect 495 988 529 1010
rect 495 976 529 988
rect 495 920 529 938
rect 495 904 529 920
rect 495 852 529 866
rect 495 832 529 852
rect 495 784 529 794
rect 495 760 529 784
rect 495 716 529 722
rect 495 688 529 716
rect 495 648 529 650
rect 495 616 529 648
rect 495 546 529 578
rect 495 544 529 546
rect 495 478 529 506
rect 495 472 529 478
rect 495 410 529 434
rect 495 400 529 410
rect 495 342 529 362
rect 495 328 529 342
rect 495 274 529 290
rect 495 256 529 274
rect 495 206 529 218
rect 495 184 529 206
rect 495 138 529 146
rect 495 112 529 138
rect 651 1056 685 1082
rect 651 1048 685 1056
rect 651 988 685 1010
rect 651 976 685 988
rect 651 920 685 938
rect 651 904 685 920
rect 651 852 685 866
rect 651 832 685 852
rect 651 784 685 794
rect 651 760 685 784
rect 651 716 685 722
rect 651 688 685 716
rect 651 648 685 650
rect 651 616 685 648
rect 651 546 685 578
rect 651 544 685 546
rect 651 478 685 506
rect 651 472 685 478
rect 651 410 685 434
rect 651 400 685 410
rect 651 342 685 362
rect 651 328 685 342
rect 651 274 685 290
rect 651 256 685 274
rect 651 206 685 218
rect 651 184 685 206
rect 651 138 685 146
rect 651 112 685 138
rect 807 1056 841 1082
rect 807 1048 841 1056
rect 807 988 841 1010
rect 807 976 841 988
rect 807 920 841 938
rect 807 904 841 920
rect 807 852 841 866
rect 807 832 841 852
rect 807 784 841 794
rect 807 760 841 784
rect 807 716 841 722
rect 807 688 841 716
rect 807 648 841 650
rect 807 616 841 648
rect 807 546 841 578
rect 807 544 841 546
rect 807 478 841 506
rect 807 472 841 478
rect 807 410 841 434
rect 807 400 841 410
rect 807 342 841 362
rect 807 328 841 342
rect 807 274 841 290
rect 807 256 841 274
rect 807 206 841 218
rect 807 184 841 206
rect 807 138 841 146
rect 807 112 841 138
rect 963 1056 997 1082
rect 963 1048 997 1056
rect 963 988 997 1010
rect 963 976 997 988
rect 963 920 997 938
rect 963 904 997 920
rect 963 852 997 866
rect 963 832 997 852
rect 963 784 997 794
rect 963 760 997 784
rect 963 716 997 722
rect 963 688 997 716
rect 963 648 997 650
rect 963 616 997 648
rect 963 546 997 578
rect 963 544 997 546
rect 963 478 997 506
rect 963 472 997 478
rect 963 410 997 434
rect 963 400 997 410
rect 963 342 997 362
rect 963 328 997 342
rect 963 274 997 290
rect 963 256 997 274
rect 963 206 997 218
rect 963 184 997 206
rect 963 138 997 146
rect 963 112 997 138
rect 1119 1056 1153 1082
rect 1119 1048 1153 1056
rect 1119 988 1153 1010
rect 1119 976 1153 988
rect 1119 920 1153 938
rect 1119 904 1153 920
rect 1119 852 1153 866
rect 1119 832 1153 852
rect 1119 784 1153 794
rect 1119 760 1153 784
rect 1119 716 1153 722
rect 1119 688 1153 716
rect 1119 648 1153 650
rect 1119 616 1153 648
rect 1119 546 1153 578
rect 1119 544 1153 546
rect 1119 478 1153 506
rect 1119 472 1153 478
rect 1119 410 1153 434
rect 1119 400 1153 410
rect 1119 342 1153 362
rect 1119 328 1153 342
rect 1119 274 1153 290
rect 1119 256 1153 274
rect 1119 206 1153 218
rect 1119 184 1153 206
rect 1119 138 1153 146
rect 1119 112 1153 138
rect 1275 1056 1309 1082
rect 1275 1048 1309 1056
rect 1275 988 1309 1010
rect 1275 976 1309 988
rect 1275 920 1309 938
rect 1275 904 1309 920
rect 1275 852 1309 866
rect 1275 832 1309 852
rect 1275 784 1309 794
rect 1275 760 1309 784
rect 1275 716 1309 722
rect 1275 688 1309 716
rect 1275 648 1309 650
rect 1275 616 1309 648
rect 1275 546 1309 578
rect 1275 544 1309 546
rect 1275 478 1309 506
rect 1275 472 1309 478
rect 1275 410 1309 434
rect 1275 400 1309 410
rect 1275 342 1309 362
rect 1275 328 1309 342
rect 1275 274 1309 290
rect 1275 256 1309 274
rect 1275 206 1309 218
rect 1275 184 1309 206
rect 1275 138 1309 146
rect 1275 112 1309 138
rect 1431 1056 1465 1082
rect 1431 1048 1465 1056
rect 1431 988 1465 1010
rect 1431 976 1465 988
rect 1431 920 1465 938
rect 1431 904 1465 920
rect 1431 852 1465 866
rect 1431 832 1465 852
rect 1431 784 1465 794
rect 1431 760 1465 784
rect 1431 716 1465 722
rect 1431 688 1465 716
rect 1431 648 1465 650
rect 1431 616 1465 648
rect 1431 546 1465 578
rect 1431 544 1465 546
rect 1431 478 1465 506
rect 1431 472 1465 478
rect 1431 410 1465 434
rect 1431 400 1465 410
rect 1431 342 1465 362
rect 1431 328 1465 342
rect 1431 274 1465 290
rect 1431 256 1465 274
rect 1431 206 1465 218
rect 1431 184 1465 206
rect 1431 138 1465 146
rect 1431 112 1465 138
rect 1587 1056 1621 1082
rect 1587 1048 1621 1056
rect 1587 988 1621 1010
rect 1587 976 1621 988
rect 1587 920 1621 938
rect 1587 904 1621 920
rect 1587 852 1621 866
rect 1587 832 1621 852
rect 1587 784 1621 794
rect 1587 760 1621 784
rect 1587 716 1621 722
rect 1587 688 1621 716
rect 1587 648 1621 650
rect 1587 616 1621 648
rect 1587 546 1621 578
rect 1587 544 1621 546
rect 1587 478 1621 506
rect 1587 472 1621 478
rect 1587 410 1621 434
rect 1587 400 1621 410
rect 1587 342 1621 362
rect 1587 328 1621 342
rect 1587 274 1621 290
rect 1587 256 1621 274
rect 1587 206 1621 218
rect 1587 184 1621 206
rect 1587 138 1621 146
rect 1587 112 1621 138
rect 1743 1056 1777 1082
rect 1743 1048 1777 1056
rect 1743 988 1777 1010
rect 1743 976 1777 988
rect 1743 920 1777 938
rect 1743 904 1777 920
rect 1743 852 1777 866
rect 1743 832 1777 852
rect 1743 784 1777 794
rect 1743 760 1777 784
rect 1743 716 1777 722
rect 1743 688 1777 716
rect 1743 648 1777 650
rect 1743 616 1777 648
rect 1743 546 1777 578
rect 1743 544 1777 546
rect 1743 478 1777 506
rect 1743 472 1777 478
rect 1743 410 1777 434
rect 1743 400 1777 410
rect 1743 342 1777 362
rect 1743 328 1777 342
rect 1743 274 1777 290
rect 1743 256 1777 274
rect 1743 206 1777 218
rect 1743 184 1777 206
rect 1743 138 1777 146
rect 1743 112 1777 138
rect 1878 1056 1912 1082
rect 1878 1048 1912 1056
rect 1878 988 1912 1010
rect 1878 976 1912 988
rect 1878 920 1912 938
rect 1878 904 1912 920
rect 1878 852 1912 866
rect 1878 832 1912 852
rect 1878 784 1912 794
rect 1878 760 1912 784
rect 1878 716 1912 722
rect 1878 688 1912 716
rect 1878 648 1912 650
rect 1878 616 1912 648
rect 1878 546 1912 578
rect 1878 544 1912 546
rect 1878 478 1912 506
rect 1878 472 1912 478
rect 1878 410 1912 434
rect 1878 400 1912 410
rect 1878 342 1912 362
rect 1878 328 1912 342
rect 1878 274 1912 290
rect 1878 256 1912 274
rect 1878 206 1912 218
rect 1878 184 1912 206
rect 1878 138 1912 146
rect 1878 112 1912 138
rect 207 20 215 54
rect 215 20 241 54
rect 279 20 283 54
rect 283 20 313 54
rect 351 20 385 54
rect 423 20 453 54
rect 453 20 457 54
rect 495 20 521 54
rect 521 20 529 54
rect 567 20 589 54
rect 589 20 601 54
rect 639 20 657 54
rect 657 20 673 54
rect 711 20 725 54
rect 725 20 745 54
rect 783 20 793 54
rect 793 20 817 54
rect 855 20 861 54
rect 861 20 889 54
rect 927 20 929 54
rect 929 20 961 54
rect 999 20 1031 54
rect 1031 20 1033 54
rect 1071 20 1099 54
rect 1099 20 1105 54
rect 1143 20 1167 54
rect 1167 20 1177 54
rect 1215 20 1235 54
rect 1235 20 1249 54
rect 1287 20 1303 54
rect 1303 20 1321 54
rect 1359 20 1371 54
rect 1371 20 1393 54
rect 1431 20 1439 54
rect 1439 20 1465 54
rect 1503 20 1507 54
rect 1507 20 1537 54
rect 1575 20 1609 54
rect 1647 20 1677 54
rect 1677 20 1681 54
rect 1719 20 1745 54
rect 1745 20 1753 54
<< metal1 >>
rect 195 1174 1765 1194
rect 195 1140 207 1174
rect 241 1140 279 1174
rect 313 1140 351 1174
rect 385 1140 423 1174
rect 457 1140 495 1174
rect 529 1140 567 1174
rect 601 1140 639 1174
rect 673 1140 711 1174
rect 745 1140 783 1174
rect 817 1140 855 1174
rect 889 1140 927 1174
rect 961 1140 999 1174
rect 1033 1140 1071 1174
rect 1105 1140 1143 1174
rect 1177 1140 1215 1174
rect 1249 1140 1287 1174
rect 1321 1140 1359 1174
rect 1393 1140 1431 1174
rect 1465 1140 1503 1174
rect 1537 1140 1575 1174
rect 1609 1140 1647 1174
rect 1681 1140 1719 1174
rect 1753 1140 1765 1174
rect 195 1128 1765 1140
rect 36 1082 95 1094
rect 36 1048 48 1082
rect 82 1048 95 1082
rect 36 1010 95 1048
rect 36 976 48 1010
rect 82 976 95 1010
rect 36 938 95 976
rect 36 904 48 938
rect 82 904 95 938
rect 36 866 95 904
rect 36 832 48 866
rect 82 832 95 866
rect 36 794 95 832
rect 36 760 48 794
rect 82 760 95 794
rect 36 722 95 760
rect 36 688 48 722
rect 82 688 95 722
rect 36 650 95 688
rect 36 616 48 650
rect 82 616 95 650
rect 36 578 95 616
rect 36 544 48 578
rect 82 544 95 578
rect 36 506 95 544
rect 36 472 48 506
rect 82 472 95 506
rect 36 434 95 472
rect 36 400 48 434
rect 82 400 95 434
rect 36 362 95 400
rect 36 328 48 362
rect 82 328 95 362
rect 36 290 95 328
rect 36 256 48 290
rect 82 256 95 290
rect 36 218 95 256
rect 36 184 48 218
rect 82 184 95 218
rect 36 146 95 184
rect 36 112 48 146
rect 82 112 95 146
rect 36 100 95 112
rect 174 1082 226 1094
rect 174 1048 183 1082
rect 217 1048 226 1082
rect 174 1010 226 1048
rect 174 976 183 1010
rect 217 976 226 1010
rect 174 938 226 976
rect 174 904 183 938
rect 217 904 226 938
rect 174 866 226 904
rect 174 832 183 866
rect 217 832 226 866
rect 174 794 226 832
rect 174 760 183 794
rect 217 760 226 794
rect 174 722 226 760
rect 174 688 183 722
rect 217 688 226 722
rect 174 650 226 688
rect 174 616 183 650
rect 217 616 226 650
rect 174 578 226 616
rect 174 544 183 578
rect 217 544 226 578
rect 174 542 226 544
rect 174 478 183 490
rect 217 478 226 490
rect 174 414 183 426
rect 217 414 226 426
rect 174 350 183 362
rect 217 350 226 362
rect 174 290 226 298
rect 174 286 183 290
rect 217 286 226 290
rect 174 222 226 234
rect 174 158 226 170
rect 174 100 226 106
rect 330 1088 382 1094
rect 330 1024 382 1036
rect 330 960 382 972
rect 330 904 339 908
rect 373 904 382 908
rect 330 896 382 904
rect 330 832 339 844
rect 373 832 382 844
rect 330 768 339 780
rect 373 768 382 780
rect 330 704 339 716
rect 373 704 382 716
rect 330 650 382 652
rect 330 616 339 650
rect 373 616 382 650
rect 330 578 382 616
rect 330 544 339 578
rect 373 544 382 578
rect 330 506 382 544
rect 330 472 339 506
rect 373 472 382 506
rect 330 434 382 472
rect 330 400 339 434
rect 373 400 382 434
rect 330 362 382 400
rect 330 328 339 362
rect 373 328 382 362
rect 330 290 382 328
rect 330 256 339 290
rect 373 256 382 290
rect 330 218 382 256
rect 330 184 339 218
rect 373 184 382 218
rect 330 146 382 184
rect 330 112 339 146
rect 373 112 382 146
rect 330 100 382 112
rect 486 1082 538 1094
rect 486 1048 495 1082
rect 529 1048 538 1082
rect 486 1010 538 1048
rect 486 976 495 1010
rect 529 976 538 1010
rect 486 938 538 976
rect 486 904 495 938
rect 529 904 538 938
rect 486 866 538 904
rect 486 832 495 866
rect 529 832 538 866
rect 486 794 538 832
rect 486 760 495 794
rect 529 760 538 794
rect 486 722 538 760
rect 486 688 495 722
rect 529 688 538 722
rect 486 650 538 688
rect 486 616 495 650
rect 529 616 538 650
rect 486 578 538 616
rect 486 544 495 578
rect 529 544 538 578
rect 486 542 538 544
rect 486 478 495 490
rect 529 478 538 490
rect 486 414 495 426
rect 529 414 538 426
rect 486 350 495 362
rect 529 350 538 362
rect 486 290 538 298
rect 486 286 495 290
rect 529 286 538 290
rect 486 222 538 234
rect 486 158 538 170
rect 486 100 538 106
rect 642 1088 694 1094
rect 642 1024 694 1036
rect 642 960 694 972
rect 642 904 651 908
rect 685 904 694 908
rect 642 896 694 904
rect 642 832 651 844
rect 685 832 694 844
rect 642 768 651 780
rect 685 768 694 780
rect 642 704 651 716
rect 685 704 694 716
rect 642 650 694 652
rect 642 616 651 650
rect 685 616 694 650
rect 642 578 694 616
rect 642 544 651 578
rect 685 544 694 578
rect 642 506 694 544
rect 642 472 651 506
rect 685 472 694 506
rect 642 434 694 472
rect 642 400 651 434
rect 685 400 694 434
rect 642 362 694 400
rect 642 328 651 362
rect 685 328 694 362
rect 642 290 694 328
rect 642 256 651 290
rect 685 256 694 290
rect 642 218 694 256
rect 642 184 651 218
rect 685 184 694 218
rect 642 146 694 184
rect 642 112 651 146
rect 685 112 694 146
rect 642 100 694 112
rect 798 1082 850 1094
rect 798 1048 807 1082
rect 841 1048 850 1082
rect 798 1010 850 1048
rect 798 976 807 1010
rect 841 976 850 1010
rect 798 938 850 976
rect 798 904 807 938
rect 841 904 850 938
rect 798 866 850 904
rect 798 832 807 866
rect 841 832 850 866
rect 798 794 850 832
rect 798 760 807 794
rect 841 760 850 794
rect 798 722 850 760
rect 798 688 807 722
rect 841 688 850 722
rect 798 650 850 688
rect 798 616 807 650
rect 841 616 850 650
rect 798 578 850 616
rect 798 544 807 578
rect 841 544 850 578
rect 798 542 850 544
rect 798 478 807 490
rect 841 478 850 490
rect 798 414 807 426
rect 841 414 850 426
rect 798 350 807 362
rect 841 350 850 362
rect 798 290 850 298
rect 798 286 807 290
rect 841 286 850 290
rect 798 222 850 234
rect 798 158 850 170
rect 798 100 850 106
rect 954 1088 1006 1094
rect 954 1024 1006 1036
rect 954 960 1006 972
rect 954 904 963 908
rect 997 904 1006 908
rect 954 896 1006 904
rect 954 832 963 844
rect 997 832 1006 844
rect 954 768 963 780
rect 997 768 1006 780
rect 954 704 963 716
rect 997 704 1006 716
rect 954 650 1006 652
rect 954 616 963 650
rect 997 616 1006 650
rect 954 578 1006 616
rect 954 544 963 578
rect 997 544 1006 578
rect 954 506 1006 544
rect 954 472 963 506
rect 997 472 1006 506
rect 954 434 1006 472
rect 954 400 963 434
rect 997 400 1006 434
rect 954 362 1006 400
rect 954 328 963 362
rect 997 328 1006 362
rect 954 290 1006 328
rect 954 256 963 290
rect 997 256 1006 290
rect 954 218 1006 256
rect 954 184 963 218
rect 997 184 1006 218
rect 954 146 1006 184
rect 954 112 963 146
rect 997 112 1006 146
rect 954 100 1006 112
rect 1110 1082 1162 1094
rect 1110 1048 1119 1082
rect 1153 1048 1162 1082
rect 1110 1010 1162 1048
rect 1110 976 1119 1010
rect 1153 976 1162 1010
rect 1110 938 1162 976
rect 1110 904 1119 938
rect 1153 904 1162 938
rect 1110 866 1162 904
rect 1110 832 1119 866
rect 1153 832 1162 866
rect 1110 794 1162 832
rect 1110 760 1119 794
rect 1153 760 1162 794
rect 1110 722 1162 760
rect 1110 688 1119 722
rect 1153 688 1162 722
rect 1110 650 1162 688
rect 1110 616 1119 650
rect 1153 616 1162 650
rect 1110 578 1162 616
rect 1110 544 1119 578
rect 1153 544 1162 578
rect 1110 542 1162 544
rect 1110 478 1119 490
rect 1153 478 1162 490
rect 1110 414 1119 426
rect 1153 414 1162 426
rect 1110 350 1119 362
rect 1153 350 1162 362
rect 1110 290 1162 298
rect 1110 286 1119 290
rect 1153 286 1162 290
rect 1110 222 1162 234
rect 1110 158 1162 170
rect 1110 100 1162 106
rect 1266 1088 1318 1094
rect 1266 1024 1318 1036
rect 1266 960 1318 972
rect 1266 904 1275 908
rect 1309 904 1318 908
rect 1266 896 1318 904
rect 1266 832 1275 844
rect 1309 832 1318 844
rect 1266 768 1275 780
rect 1309 768 1318 780
rect 1266 704 1275 716
rect 1309 704 1318 716
rect 1266 650 1318 652
rect 1266 616 1275 650
rect 1309 616 1318 650
rect 1266 578 1318 616
rect 1266 544 1275 578
rect 1309 544 1318 578
rect 1266 506 1318 544
rect 1266 472 1275 506
rect 1309 472 1318 506
rect 1266 434 1318 472
rect 1266 400 1275 434
rect 1309 400 1318 434
rect 1266 362 1318 400
rect 1266 328 1275 362
rect 1309 328 1318 362
rect 1266 290 1318 328
rect 1266 256 1275 290
rect 1309 256 1318 290
rect 1266 218 1318 256
rect 1266 184 1275 218
rect 1309 184 1318 218
rect 1266 146 1318 184
rect 1266 112 1275 146
rect 1309 112 1318 146
rect 1266 100 1318 112
rect 1422 1082 1474 1094
rect 1422 1048 1431 1082
rect 1465 1048 1474 1082
rect 1422 1010 1474 1048
rect 1422 976 1431 1010
rect 1465 976 1474 1010
rect 1422 938 1474 976
rect 1422 904 1431 938
rect 1465 904 1474 938
rect 1422 866 1474 904
rect 1422 832 1431 866
rect 1465 832 1474 866
rect 1422 794 1474 832
rect 1422 760 1431 794
rect 1465 760 1474 794
rect 1422 722 1474 760
rect 1422 688 1431 722
rect 1465 688 1474 722
rect 1422 650 1474 688
rect 1422 616 1431 650
rect 1465 616 1474 650
rect 1422 578 1474 616
rect 1422 544 1431 578
rect 1465 544 1474 578
rect 1422 542 1474 544
rect 1422 478 1431 490
rect 1465 478 1474 490
rect 1422 414 1431 426
rect 1465 414 1474 426
rect 1422 350 1431 362
rect 1465 350 1474 362
rect 1422 290 1474 298
rect 1422 286 1431 290
rect 1465 286 1474 290
rect 1422 222 1474 234
rect 1422 158 1474 170
rect 1422 100 1474 106
rect 1578 1088 1630 1094
rect 1578 1024 1630 1036
rect 1578 960 1630 972
rect 1578 904 1587 908
rect 1621 904 1630 908
rect 1578 896 1630 904
rect 1578 832 1587 844
rect 1621 832 1630 844
rect 1578 768 1587 780
rect 1621 768 1630 780
rect 1578 704 1587 716
rect 1621 704 1630 716
rect 1578 650 1630 652
rect 1578 616 1587 650
rect 1621 616 1630 650
rect 1578 578 1630 616
rect 1578 544 1587 578
rect 1621 544 1630 578
rect 1578 506 1630 544
rect 1578 472 1587 506
rect 1621 472 1630 506
rect 1578 434 1630 472
rect 1578 400 1587 434
rect 1621 400 1630 434
rect 1578 362 1630 400
rect 1578 328 1587 362
rect 1621 328 1630 362
rect 1578 290 1630 328
rect 1578 256 1587 290
rect 1621 256 1630 290
rect 1578 218 1630 256
rect 1578 184 1587 218
rect 1621 184 1630 218
rect 1578 146 1630 184
rect 1578 112 1587 146
rect 1621 112 1630 146
rect 1578 100 1630 112
rect 1734 1082 1786 1094
rect 1734 1048 1743 1082
rect 1777 1048 1786 1082
rect 1734 1010 1786 1048
rect 1734 976 1743 1010
rect 1777 976 1786 1010
rect 1734 938 1786 976
rect 1734 904 1743 938
rect 1777 904 1786 938
rect 1734 866 1786 904
rect 1734 832 1743 866
rect 1777 832 1786 866
rect 1734 794 1786 832
rect 1734 760 1743 794
rect 1777 760 1786 794
rect 1734 722 1786 760
rect 1734 688 1743 722
rect 1777 688 1786 722
rect 1734 650 1786 688
rect 1734 616 1743 650
rect 1777 616 1786 650
rect 1734 578 1786 616
rect 1734 544 1743 578
rect 1777 544 1786 578
rect 1734 542 1786 544
rect 1734 478 1743 490
rect 1777 478 1786 490
rect 1734 414 1743 426
rect 1777 414 1786 426
rect 1734 350 1743 362
rect 1777 350 1786 362
rect 1734 290 1786 298
rect 1734 286 1743 290
rect 1777 286 1786 290
rect 1734 222 1786 234
rect 1734 158 1786 170
rect 1734 100 1786 106
rect 1866 1082 1925 1094
rect 1866 1048 1878 1082
rect 1912 1048 1925 1082
rect 1866 1010 1925 1048
rect 1866 976 1878 1010
rect 1912 976 1925 1010
rect 1866 938 1925 976
rect 1866 904 1878 938
rect 1912 904 1925 938
rect 1866 866 1925 904
rect 1866 832 1878 866
rect 1912 832 1925 866
rect 1866 794 1925 832
rect 1866 760 1878 794
rect 1912 760 1925 794
rect 1866 722 1925 760
rect 1866 688 1878 722
rect 1912 688 1925 722
rect 1866 650 1925 688
rect 1866 616 1878 650
rect 1912 616 1925 650
rect 1866 578 1925 616
rect 1866 544 1878 578
rect 1912 544 1925 578
rect 1866 506 1925 544
rect 1866 472 1878 506
rect 1912 472 1925 506
rect 1866 434 1925 472
rect 1866 400 1878 434
rect 1912 400 1925 434
rect 1866 362 1925 400
rect 1866 328 1878 362
rect 1912 328 1925 362
rect 1866 290 1925 328
rect 1866 256 1878 290
rect 1912 256 1925 290
rect 1866 218 1925 256
rect 1866 184 1878 218
rect 1912 184 1925 218
rect 1866 146 1925 184
rect 1866 112 1878 146
rect 1912 112 1925 146
rect 1866 100 1925 112
rect 195 54 1765 66
rect 195 20 207 54
rect 241 20 279 54
rect 313 20 351 54
rect 385 20 423 54
rect 457 20 495 54
rect 529 20 567 54
rect 601 20 639 54
rect 673 20 711 54
rect 745 20 783 54
rect 817 20 855 54
rect 889 20 927 54
rect 961 20 999 54
rect 1033 20 1071 54
rect 1105 20 1143 54
rect 1177 20 1215 54
rect 1249 20 1287 54
rect 1321 20 1359 54
rect 1393 20 1431 54
rect 1465 20 1503 54
rect 1537 20 1575 54
rect 1609 20 1647 54
rect 1681 20 1719 54
rect 1753 20 1765 54
rect 195 0 1765 20
<< via1 >>
rect 174 506 226 542
rect 174 490 183 506
rect 183 490 217 506
rect 217 490 226 506
rect 174 472 183 478
rect 183 472 217 478
rect 217 472 226 478
rect 174 434 226 472
rect 174 426 183 434
rect 183 426 217 434
rect 217 426 226 434
rect 174 400 183 414
rect 183 400 217 414
rect 217 400 226 414
rect 174 362 226 400
rect 174 328 183 350
rect 183 328 217 350
rect 217 328 226 350
rect 174 298 226 328
rect 174 256 183 286
rect 183 256 217 286
rect 217 256 226 286
rect 174 234 226 256
rect 174 218 226 222
rect 174 184 183 218
rect 183 184 217 218
rect 217 184 226 218
rect 174 170 226 184
rect 174 146 226 158
rect 174 112 183 146
rect 183 112 217 146
rect 217 112 226 146
rect 174 106 226 112
rect 330 1082 382 1088
rect 330 1048 339 1082
rect 339 1048 373 1082
rect 373 1048 382 1082
rect 330 1036 382 1048
rect 330 1010 382 1024
rect 330 976 339 1010
rect 339 976 373 1010
rect 373 976 382 1010
rect 330 972 382 976
rect 330 938 382 960
rect 330 908 339 938
rect 339 908 373 938
rect 373 908 382 938
rect 330 866 382 896
rect 330 844 339 866
rect 339 844 373 866
rect 373 844 382 866
rect 330 794 382 832
rect 330 780 339 794
rect 339 780 373 794
rect 373 780 382 794
rect 330 760 339 768
rect 339 760 373 768
rect 373 760 382 768
rect 330 722 382 760
rect 330 716 339 722
rect 339 716 373 722
rect 373 716 382 722
rect 330 688 339 704
rect 339 688 373 704
rect 373 688 382 704
rect 330 652 382 688
rect 486 506 538 542
rect 486 490 495 506
rect 495 490 529 506
rect 529 490 538 506
rect 486 472 495 478
rect 495 472 529 478
rect 529 472 538 478
rect 486 434 538 472
rect 486 426 495 434
rect 495 426 529 434
rect 529 426 538 434
rect 486 400 495 414
rect 495 400 529 414
rect 529 400 538 414
rect 486 362 538 400
rect 486 328 495 350
rect 495 328 529 350
rect 529 328 538 350
rect 486 298 538 328
rect 486 256 495 286
rect 495 256 529 286
rect 529 256 538 286
rect 486 234 538 256
rect 486 218 538 222
rect 486 184 495 218
rect 495 184 529 218
rect 529 184 538 218
rect 486 170 538 184
rect 486 146 538 158
rect 486 112 495 146
rect 495 112 529 146
rect 529 112 538 146
rect 486 106 538 112
rect 642 1082 694 1088
rect 642 1048 651 1082
rect 651 1048 685 1082
rect 685 1048 694 1082
rect 642 1036 694 1048
rect 642 1010 694 1024
rect 642 976 651 1010
rect 651 976 685 1010
rect 685 976 694 1010
rect 642 972 694 976
rect 642 938 694 960
rect 642 908 651 938
rect 651 908 685 938
rect 685 908 694 938
rect 642 866 694 896
rect 642 844 651 866
rect 651 844 685 866
rect 685 844 694 866
rect 642 794 694 832
rect 642 780 651 794
rect 651 780 685 794
rect 685 780 694 794
rect 642 760 651 768
rect 651 760 685 768
rect 685 760 694 768
rect 642 722 694 760
rect 642 716 651 722
rect 651 716 685 722
rect 685 716 694 722
rect 642 688 651 704
rect 651 688 685 704
rect 685 688 694 704
rect 642 652 694 688
rect 798 506 850 542
rect 798 490 807 506
rect 807 490 841 506
rect 841 490 850 506
rect 798 472 807 478
rect 807 472 841 478
rect 841 472 850 478
rect 798 434 850 472
rect 798 426 807 434
rect 807 426 841 434
rect 841 426 850 434
rect 798 400 807 414
rect 807 400 841 414
rect 841 400 850 414
rect 798 362 850 400
rect 798 328 807 350
rect 807 328 841 350
rect 841 328 850 350
rect 798 298 850 328
rect 798 256 807 286
rect 807 256 841 286
rect 841 256 850 286
rect 798 234 850 256
rect 798 218 850 222
rect 798 184 807 218
rect 807 184 841 218
rect 841 184 850 218
rect 798 170 850 184
rect 798 146 850 158
rect 798 112 807 146
rect 807 112 841 146
rect 841 112 850 146
rect 798 106 850 112
rect 954 1082 1006 1088
rect 954 1048 963 1082
rect 963 1048 997 1082
rect 997 1048 1006 1082
rect 954 1036 1006 1048
rect 954 1010 1006 1024
rect 954 976 963 1010
rect 963 976 997 1010
rect 997 976 1006 1010
rect 954 972 1006 976
rect 954 938 1006 960
rect 954 908 963 938
rect 963 908 997 938
rect 997 908 1006 938
rect 954 866 1006 896
rect 954 844 963 866
rect 963 844 997 866
rect 997 844 1006 866
rect 954 794 1006 832
rect 954 780 963 794
rect 963 780 997 794
rect 997 780 1006 794
rect 954 760 963 768
rect 963 760 997 768
rect 997 760 1006 768
rect 954 722 1006 760
rect 954 716 963 722
rect 963 716 997 722
rect 997 716 1006 722
rect 954 688 963 704
rect 963 688 997 704
rect 997 688 1006 704
rect 954 652 1006 688
rect 1110 506 1162 542
rect 1110 490 1119 506
rect 1119 490 1153 506
rect 1153 490 1162 506
rect 1110 472 1119 478
rect 1119 472 1153 478
rect 1153 472 1162 478
rect 1110 434 1162 472
rect 1110 426 1119 434
rect 1119 426 1153 434
rect 1153 426 1162 434
rect 1110 400 1119 414
rect 1119 400 1153 414
rect 1153 400 1162 414
rect 1110 362 1162 400
rect 1110 328 1119 350
rect 1119 328 1153 350
rect 1153 328 1162 350
rect 1110 298 1162 328
rect 1110 256 1119 286
rect 1119 256 1153 286
rect 1153 256 1162 286
rect 1110 234 1162 256
rect 1110 218 1162 222
rect 1110 184 1119 218
rect 1119 184 1153 218
rect 1153 184 1162 218
rect 1110 170 1162 184
rect 1110 146 1162 158
rect 1110 112 1119 146
rect 1119 112 1153 146
rect 1153 112 1162 146
rect 1110 106 1162 112
rect 1266 1082 1318 1088
rect 1266 1048 1275 1082
rect 1275 1048 1309 1082
rect 1309 1048 1318 1082
rect 1266 1036 1318 1048
rect 1266 1010 1318 1024
rect 1266 976 1275 1010
rect 1275 976 1309 1010
rect 1309 976 1318 1010
rect 1266 972 1318 976
rect 1266 938 1318 960
rect 1266 908 1275 938
rect 1275 908 1309 938
rect 1309 908 1318 938
rect 1266 866 1318 896
rect 1266 844 1275 866
rect 1275 844 1309 866
rect 1309 844 1318 866
rect 1266 794 1318 832
rect 1266 780 1275 794
rect 1275 780 1309 794
rect 1309 780 1318 794
rect 1266 760 1275 768
rect 1275 760 1309 768
rect 1309 760 1318 768
rect 1266 722 1318 760
rect 1266 716 1275 722
rect 1275 716 1309 722
rect 1309 716 1318 722
rect 1266 688 1275 704
rect 1275 688 1309 704
rect 1309 688 1318 704
rect 1266 652 1318 688
rect 1422 506 1474 542
rect 1422 490 1431 506
rect 1431 490 1465 506
rect 1465 490 1474 506
rect 1422 472 1431 478
rect 1431 472 1465 478
rect 1465 472 1474 478
rect 1422 434 1474 472
rect 1422 426 1431 434
rect 1431 426 1465 434
rect 1465 426 1474 434
rect 1422 400 1431 414
rect 1431 400 1465 414
rect 1465 400 1474 414
rect 1422 362 1474 400
rect 1422 328 1431 350
rect 1431 328 1465 350
rect 1465 328 1474 350
rect 1422 298 1474 328
rect 1422 256 1431 286
rect 1431 256 1465 286
rect 1465 256 1474 286
rect 1422 234 1474 256
rect 1422 218 1474 222
rect 1422 184 1431 218
rect 1431 184 1465 218
rect 1465 184 1474 218
rect 1422 170 1474 184
rect 1422 146 1474 158
rect 1422 112 1431 146
rect 1431 112 1465 146
rect 1465 112 1474 146
rect 1422 106 1474 112
rect 1578 1082 1630 1088
rect 1578 1048 1587 1082
rect 1587 1048 1621 1082
rect 1621 1048 1630 1082
rect 1578 1036 1630 1048
rect 1578 1010 1630 1024
rect 1578 976 1587 1010
rect 1587 976 1621 1010
rect 1621 976 1630 1010
rect 1578 972 1630 976
rect 1578 938 1630 960
rect 1578 908 1587 938
rect 1587 908 1621 938
rect 1621 908 1630 938
rect 1578 866 1630 896
rect 1578 844 1587 866
rect 1587 844 1621 866
rect 1621 844 1630 866
rect 1578 794 1630 832
rect 1578 780 1587 794
rect 1587 780 1621 794
rect 1621 780 1630 794
rect 1578 760 1587 768
rect 1587 760 1621 768
rect 1621 760 1630 768
rect 1578 722 1630 760
rect 1578 716 1587 722
rect 1587 716 1621 722
rect 1621 716 1630 722
rect 1578 688 1587 704
rect 1587 688 1621 704
rect 1621 688 1630 704
rect 1578 652 1630 688
rect 1734 506 1786 542
rect 1734 490 1743 506
rect 1743 490 1777 506
rect 1777 490 1786 506
rect 1734 472 1743 478
rect 1743 472 1777 478
rect 1777 472 1786 478
rect 1734 434 1786 472
rect 1734 426 1743 434
rect 1743 426 1777 434
rect 1777 426 1786 434
rect 1734 400 1743 414
rect 1743 400 1777 414
rect 1777 400 1786 414
rect 1734 362 1786 400
rect 1734 328 1743 350
rect 1743 328 1777 350
rect 1777 328 1786 350
rect 1734 298 1786 328
rect 1734 256 1743 286
rect 1743 256 1777 286
rect 1777 256 1786 286
rect 1734 234 1786 256
rect 1734 218 1786 222
rect 1734 184 1743 218
rect 1743 184 1777 218
rect 1777 184 1786 218
rect 1734 170 1786 184
rect 1734 146 1786 158
rect 1734 112 1743 146
rect 1743 112 1777 146
rect 1777 112 1786 146
rect 1734 106 1786 112
<< metal2 >>
rect 14 1088 1946 1094
rect 14 1036 330 1088
rect 382 1036 642 1088
rect 694 1036 954 1088
rect 1006 1036 1266 1088
rect 1318 1036 1578 1088
rect 1630 1036 1946 1088
rect 14 1024 1946 1036
rect 14 972 330 1024
rect 382 972 642 1024
rect 694 972 954 1024
rect 1006 972 1266 1024
rect 1318 972 1578 1024
rect 1630 972 1946 1024
rect 14 960 1946 972
rect 14 908 330 960
rect 382 908 642 960
rect 694 908 954 960
rect 1006 908 1266 960
rect 1318 908 1578 960
rect 1630 908 1946 960
rect 14 896 1946 908
rect 14 844 330 896
rect 382 844 642 896
rect 694 844 954 896
rect 1006 844 1266 896
rect 1318 844 1578 896
rect 1630 844 1946 896
rect 14 832 1946 844
rect 14 780 330 832
rect 382 780 642 832
rect 694 780 954 832
rect 1006 780 1266 832
rect 1318 780 1578 832
rect 1630 780 1946 832
rect 14 768 1946 780
rect 14 716 330 768
rect 382 716 642 768
rect 694 716 954 768
rect 1006 716 1266 768
rect 1318 716 1578 768
rect 1630 716 1946 768
rect 14 704 1946 716
rect 14 652 330 704
rect 382 652 642 704
rect 694 652 954 704
rect 1006 652 1266 704
rect 1318 652 1578 704
rect 1630 652 1946 704
rect 14 622 1946 652
rect 14 542 1946 572
rect 14 490 174 542
rect 226 490 486 542
rect 538 490 798 542
rect 850 490 1110 542
rect 1162 490 1422 542
rect 1474 490 1734 542
rect 1786 490 1946 542
rect 14 478 1946 490
rect 14 426 174 478
rect 226 426 486 478
rect 538 426 798 478
rect 850 426 1110 478
rect 1162 426 1422 478
rect 1474 426 1734 478
rect 1786 426 1946 478
rect 14 414 1946 426
rect 14 362 174 414
rect 226 362 486 414
rect 538 362 798 414
rect 850 362 1110 414
rect 1162 362 1422 414
rect 1474 362 1734 414
rect 1786 362 1946 414
rect 14 350 1946 362
rect 14 298 174 350
rect 226 298 486 350
rect 538 298 798 350
rect 850 298 1110 350
rect 1162 298 1422 350
rect 1474 298 1734 350
rect 1786 298 1946 350
rect 14 286 1946 298
rect 14 234 174 286
rect 226 234 486 286
rect 538 234 798 286
rect 850 234 1110 286
rect 1162 234 1422 286
rect 1474 234 1734 286
rect 1786 234 1946 286
rect 14 222 1946 234
rect 14 170 174 222
rect 226 170 486 222
rect 538 170 798 222
rect 850 170 1110 222
rect 1162 170 1422 222
rect 1474 170 1734 222
rect 1786 170 1946 222
rect 14 158 1946 170
rect 14 106 174 158
rect 226 106 486 158
rect 538 106 798 158
rect 850 106 1110 158
rect 1162 106 1422 158
rect 1474 106 1734 158
rect 1786 106 1946 158
rect 14 100 1946 106
<< labels >>
flabel metal1 s 46 554 72 621 0 FreeSans 400 90 0 0 SUBSTRATE
port 1 nsew
flabel metal1 s 933 1148 1019 1173 0 FreeSans 400 0 0 0 GATE
port 2 nsew
flabel metal1 s 1885 554 1911 621 0 FreeSans 400 90 0 0 SUBSTRATE
port 1 nsew
flabel metal2 s 122 128 198 153 0 FreeSans 400 0 0 0 SOURCE
port 3 nsew
flabel metal2 s 112 1047 201 1079 0 FreeSans 400 0 0 0 DRAIN
port 4 nsew
<< properties >>
string GDS_END 4422476
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 4379780
<< end >>
