magic
tech sky130A
magscale 1 2
timestamp 1666464484
<< nwell >>
rect 1231 8984 28211 9406
rect 1231 1044 1653 8984
rect 2067 2147 27387 8584
rect 27789 1044 28211 8984
rect 1231 742 28211 1044
<< pwell >>
rect 1779 8647 27708 8869
rect 1779 2022 2001 8647
rect 27486 2022 27708 8647
rect 1779 1276 27708 2022
<< mvpsubdiff >>
rect 1805 8775 1873 8843
rect 1839 8741 1873 8775
rect 27407 8809 27442 8843
rect 27476 8809 27511 8843
rect 27545 8809 27580 8843
rect 27614 8809 27682 8843
rect 27407 8775 27682 8809
rect 27407 8741 27442 8775
rect 27476 8741 27511 8775
rect 27545 8741 27580 8775
rect 1805 8706 1941 8741
rect 1839 8672 1873 8706
rect 1907 8673 1941 8706
rect 27339 8707 27580 8741
rect 27339 8673 27374 8707
rect 27408 8673 27443 8707
rect 27477 8673 27512 8707
rect 1907 8672 1975 8673
rect 1805 8638 1975 8672
rect 1805 8637 1941 8638
rect 1839 8603 1873 8637
rect 1907 8604 1941 8637
rect 1907 8603 1975 8604
rect 1805 8569 1975 8603
rect 1805 8568 1941 8569
rect 1839 8534 1873 8568
rect 1907 8535 1941 8568
rect 1907 8534 1975 8535
rect 1805 8500 1975 8534
rect 1805 8499 1941 8500
rect 1839 8465 1873 8499
rect 1907 8466 1941 8499
rect 1907 8465 1975 8466
rect 1805 8431 1975 8465
rect 1805 8430 1941 8431
rect 1839 8396 1873 8430
rect 1907 8397 1941 8430
rect 1907 8396 1975 8397
rect 1805 8362 1975 8396
rect 1805 8361 1941 8362
rect 1839 8327 1873 8361
rect 1907 8328 1941 8361
rect 1907 8327 1975 8328
rect 1805 8293 1975 8327
rect 1805 8292 1941 8293
rect 1839 8258 1873 8292
rect 1907 8259 1941 8292
rect 1907 8258 1975 8259
rect 1805 8224 1975 8258
rect 1805 8223 1941 8224
rect 1839 8189 1873 8223
rect 1907 8190 1941 8223
rect 1907 8189 1975 8190
rect 1805 8155 1975 8189
rect 1805 8154 1941 8155
rect 1839 8120 1873 8154
rect 1907 8121 1941 8154
rect 1907 8120 1975 8121
rect 1805 8086 1975 8120
rect 1805 8085 1941 8086
rect 1839 8051 1873 8085
rect 1907 8052 1941 8085
rect 1907 8051 1975 8052
rect 1805 8017 1975 8051
rect 1805 8016 1941 8017
rect 1839 7982 1873 8016
rect 1907 7983 1941 8016
rect 1907 7982 1975 7983
rect 1805 7948 1975 7982
rect 1805 7947 1941 7948
rect 1839 7913 1873 7947
rect 1907 7914 1941 7947
rect 1907 7913 1975 7914
rect 1805 7879 1975 7913
rect 1805 7878 1941 7879
rect 1839 7844 1873 7878
rect 1907 7845 1941 7878
rect 1907 7844 1975 7845
rect 1805 7810 1975 7844
rect 1805 7809 1941 7810
rect 1839 7775 1873 7809
rect 1907 7776 1941 7809
rect 1907 7775 1975 7776
rect 1805 7741 1975 7775
rect 1805 7740 1941 7741
rect 1839 7706 1873 7740
rect 1907 7707 1941 7740
rect 1907 7706 1975 7707
rect 1805 7672 1975 7706
rect 1805 7671 1941 7672
rect 1839 7637 1873 7671
rect 1907 7638 1941 7671
rect 1907 7637 1975 7638
rect 1805 7603 1975 7637
rect 1805 7602 1941 7603
rect 1839 7568 1873 7602
rect 1907 7569 1941 7602
rect 1907 7568 1975 7569
rect 1805 7534 1975 7568
rect 1805 7533 1941 7534
rect 1839 7499 1873 7533
rect 1907 7500 1941 7533
rect 1907 7499 1975 7500
rect 1805 7465 1975 7499
rect 1805 7464 1941 7465
rect 1839 7430 1873 7464
rect 1907 7431 1941 7464
rect 1907 7430 1975 7431
rect 1805 7396 1975 7430
rect 1805 7395 1941 7396
rect 1839 7361 1873 7395
rect 1907 7362 1941 7395
rect 1907 7361 1975 7362
rect 1805 7327 1975 7361
rect 1805 7326 1941 7327
rect 1839 7292 1873 7326
rect 1907 7293 1941 7326
rect 1907 7292 1975 7293
rect 1805 7258 1975 7292
rect 1805 7257 1941 7258
rect 1839 7223 1873 7257
rect 1907 7224 1941 7257
rect 1907 7223 1975 7224
rect 1805 7189 1975 7223
rect 1805 7188 1941 7189
rect 1839 7154 1873 7188
rect 1907 7155 1941 7188
rect 1907 7154 1975 7155
rect 1805 7120 1975 7154
rect 1805 7119 1941 7120
rect 1839 7085 1873 7119
rect 1907 7086 1941 7119
rect 1907 7085 1975 7086
rect 1805 7051 1975 7085
rect 1805 7050 1941 7051
rect 1839 7016 1873 7050
rect 1907 7017 1941 7050
rect 1907 7016 1975 7017
rect 1805 6982 1975 7016
rect 1805 6981 1941 6982
rect 1839 6947 1873 6981
rect 1907 6948 1941 6981
rect 1907 6947 1975 6948
rect 1805 6913 1975 6947
rect 1805 6912 1941 6913
rect 1839 6878 1873 6912
rect 1907 6879 1941 6912
rect 1907 6878 1975 6879
rect 1805 6844 1975 6878
rect 1805 6843 1941 6844
rect 1839 6809 1873 6843
rect 1907 6810 1941 6843
rect 1907 6809 1975 6810
rect 1805 6775 1975 6809
rect 1805 6774 1941 6775
rect 1839 6740 1873 6774
rect 1907 6741 1941 6774
rect 1907 6740 1975 6741
rect 1805 6706 1975 6740
rect 1805 6705 1941 6706
rect 1839 6671 1873 6705
rect 1907 6672 1941 6705
rect 1907 6671 1975 6672
rect 1805 6637 1975 6671
rect 1805 6636 1941 6637
rect 1839 6602 1873 6636
rect 1907 6603 1941 6636
rect 1907 6602 1975 6603
rect 1805 6568 1975 6602
rect 1805 6567 1941 6568
rect 1839 6533 1873 6567
rect 1907 6534 1941 6567
rect 1907 6533 1975 6534
rect 1805 6499 1975 6533
rect 1805 6498 1941 6499
rect 1839 6464 1873 6498
rect 1907 6465 1941 6498
rect 1907 6464 1975 6465
rect 1805 6430 1975 6464
rect 1805 6429 1941 6430
rect 1839 6395 1873 6429
rect 1907 6396 1941 6429
rect 1907 6395 1975 6396
rect 1805 6361 1975 6395
rect 1805 6360 1941 6361
rect 1839 6326 1873 6360
rect 1907 6327 1941 6360
rect 1907 6326 1975 6327
rect 1805 6292 1975 6326
rect 1805 6291 1941 6292
rect 1839 6257 1873 6291
rect 1907 6258 1941 6291
rect 1907 6257 1975 6258
rect 1805 6223 1975 6257
rect 1805 6222 1941 6223
rect 1839 6188 1873 6222
rect 1907 6189 1941 6222
rect 1907 6188 1975 6189
rect 1805 6154 1975 6188
rect 1805 6153 1941 6154
rect 1839 6119 1873 6153
rect 1907 6120 1941 6153
rect 1907 6119 1975 6120
rect 1805 6085 1975 6119
rect 1805 6084 1941 6085
rect 1839 6050 1873 6084
rect 1907 6051 1941 6084
rect 1907 6050 1975 6051
rect 1805 6016 1975 6050
rect 1805 6015 1941 6016
rect 1907 5982 1941 6015
rect 1907 5947 1975 5982
rect 1805 5369 1975 5437
rect 1839 5335 1873 5369
rect 1907 5335 1941 5369
rect 1805 5300 1975 5335
rect 1839 5266 1873 5300
rect 1907 5266 1941 5300
rect 1805 5231 1975 5266
rect 1839 5197 1873 5231
rect 1907 5197 1941 5231
rect 1805 5162 1975 5197
rect 1839 5128 1873 5162
rect 1907 5128 1941 5162
rect 1805 5093 1975 5128
rect 1839 5059 1873 5093
rect 1907 5059 1941 5093
rect 1805 5024 1975 5059
rect 1839 4990 1873 5024
rect 1907 4990 1941 5024
rect 1805 4955 1975 4990
rect 1839 4921 1873 4955
rect 1907 4921 1941 4955
rect 1805 4886 1975 4921
rect 1839 4852 1873 4886
rect 1907 4852 1941 4886
rect 1805 4817 1975 4852
rect 1839 4783 1873 4817
rect 1907 4783 1941 4817
rect 1805 4748 1975 4783
rect 1839 4714 1873 4748
rect 1907 4714 1941 4748
rect 1805 4679 1975 4714
rect 1839 4645 1873 4679
rect 1907 4645 1941 4679
rect 1805 4610 1975 4645
rect 1839 4576 1873 4610
rect 1907 4576 1941 4610
rect 1805 4541 1975 4576
rect 1839 4507 1873 4541
rect 1907 4507 1941 4541
rect 1805 4472 1975 4507
rect 1839 4438 1873 4472
rect 1907 4438 1941 4472
rect 1805 4403 1975 4438
rect 1839 4369 1873 4403
rect 1907 4369 1941 4403
rect 1805 4334 1975 4369
rect 1839 4300 1873 4334
rect 1907 4300 1941 4334
rect 1805 4265 1975 4300
rect 1839 4231 1873 4265
rect 1907 4231 1941 4265
rect 1805 4196 1975 4231
rect 1839 4162 1873 4196
rect 1907 4162 1941 4196
rect 1805 4127 1975 4162
rect 1839 4093 1873 4127
rect 1907 4093 1941 4127
rect 1805 4058 1975 4093
rect 1839 4024 1873 4058
rect 1907 4024 1941 4058
rect 1805 3989 1975 4024
rect 1839 3955 1873 3989
rect 1907 3955 1941 3989
rect 1805 3920 1975 3955
rect 27512 3266 27580 3301
rect 27546 3233 27580 3266
rect 27546 3232 27682 3233
rect 27512 3198 27682 3232
rect 27512 3197 27580 3198
rect 27546 3164 27580 3197
rect 27614 3164 27648 3198
rect 27546 3163 27682 3164
rect 27512 3129 27682 3163
rect 27512 3128 27580 3129
rect 27546 3095 27580 3128
rect 27614 3095 27648 3129
rect 27546 3094 27682 3095
rect 27512 3060 27682 3094
rect 27512 3059 27580 3060
rect 27546 3026 27580 3059
rect 27614 3026 27648 3060
rect 27546 3025 27682 3026
rect 27512 2991 27682 3025
rect 27512 2990 27580 2991
rect 27546 2957 27580 2990
rect 27614 2957 27648 2991
rect 27546 2956 27682 2957
rect 27512 2922 27682 2956
rect 27512 2921 27580 2922
rect 27546 2888 27580 2921
rect 27614 2888 27648 2922
rect 27546 2887 27682 2888
rect 27512 2853 27682 2887
rect 27512 2852 27580 2853
rect 27546 2819 27580 2852
rect 27614 2819 27648 2853
rect 27546 2818 27682 2819
rect 27512 2784 27682 2818
rect 27512 2783 27580 2784
rect 27546 2750 27580 2783
rect 27614 2750 27648 2784
rect 27546 2749 27682 2750
rect 27512 2715 27682 2749
rect 27512 2714 27580 2715
rect 27546 2681 27580 2714
rect 27614 2681 27648 2715
rect 27546 2680 27682 2681
rect 27512 2646 27682 2680
rect 27512 2645 27580 2646
rect 27546 2612 27580 2645
rect 27614 2612 27648 2646
rect 27546 2611 27682 2612
rect 27512 2577 27682 2611
rect 27512 2576 27580 2577
rect 27546 2543 27580 2576
rect 27614 2543 27648 2577
rect 27546 2542 27682 2543
rect 27512 2508 27682 2542
rect 27512 2507 27580 2508
rect 27546 2474 27580 2507
rect 27614 2474 27648 2508
rect 27546 2473 27682 2474
rect 27512 2439 27682 2473
rect 27512 2438 27580 2439
rect 27546 2405 27580 2438
rect 27614 2405 27648 2439
rect 27546 2404 27682 2405
rect 27512 2370 27682 2404
rect 27512 2369 27580 2370
rect 27546 2336 27580 2369
rect 27614 2336 27648 2370
rect 27546 2335 27682 2336
rect 27512 2301 27682 2335
rect 27512 2300 27580 2301
rect 27546 2267 27580 2300
rect 27614 2267 27648 2301
rect 27546 2266 27682 2267
rect 27512 2232 27682 2266
rect 27512 2231 27580 2232
rect 27546 2198 27580 2231
rect 27614 2198 27648 2232
rect 27546 2197 27682 2198
rect 27512 2163 27682 2197
rect 27512 2162 27580 2163
rect 27546 2129 27580 2162
rect 27614 2129 27648 2163
rect 27546 2128 27682 2129
rect 27512 2094 27682 2128
rect 27512 2093 27580 2094
rect 27546 2060 27580 2093
rect 27614 2060 27648 2094
rect 27546 2059 27682 2060
rect 27512 2025 27682 2059
rect 27512 2024 27580 2025
rect 1975 1995 27512 1996
rect 1975 1961 2009 1995
rect 2043 1961 2078 1995
rect 2112 1961 2147 1995
rect 2181 1961 2216 1995
rect 2250 1961 2284 1995
rect 2318 1961 2352 1995
rect 2386 1961 2420 1995
rect 2454 1961 2488 1995
rect 2522 1961 2556 1995
rect 2590 1961 2624 1995
rect 2658 1961 2692 1995
rect 2726 1961 2760 1995
rect 2794 1961 2828 1995
rect 2862 1961 2896 1995
rect 2930 1961 2964 1995
rect 2998 1961 3032 1995
rect 3066 1961 3100 1995
rect 3134 1961 3168 1995
rect 3202 1961 3236 1995
rect 3270 1961 3304 1995
rect 3338 1961 3372 1995
rect 3406 1961 3440 1995
rect 3474 1961 3508 1995
rect 3542 1961 3576 1995
rect 3610 1961 3644 1995
rect 3678 1961 3712 1995
rect 3746 1961 3780 1995
rect 3814 1961 3848 1995
rect 3882 1961 3916 1995
rect 3950 1961 3984 1995
rect 4018 1961 4052 1995
rect 4086 1961 4120 1995
rect 4154 1961 4188 1995
rect 4222 1961 4256 1995
rect 4290 1961 4324 1995
rect 4358 1961 4392 1995
rect 4426 1961 4460 1995
rect 4494 1961 4528 1995
rect 4562 1961 4596 1995
rect 4630 1961 4664 1995
rect 4698 1961 4732 1995
rect 4766 1961 4800 1995
rect 4834 1961 4868 1995
rect 4902 1961 4936 1995
rect 4970 1961 5004 1995
rect 5038 1961 5072 1995
rect 5106 1961 5140 1995
rect 5174 1961 5208 1995
rect 5242 1961 5276 1995
rect 5310 1961 5344 1995
rect 5378 1961 5412 1995
rect 5446 1961 5480 1995
rect 5514 1961 5548 1995
rect 5582 1961 5616 1995
rect 5650 1961 5684 1995
rect 5718 1961 5752 1995
rect 5786 1961 5820 1995
rect 5854 1961 5888 1995
rect 5922 1961 5956 1995
rect 5990 1961 6024 1995
rect 6058 1961 6092 1995
rect 6126 1961 6160 1995
rect 6194 1961 6228 1995
rect 6262 1961 6296 1995
rect 6330 1961 6364 1995
rect 6398 1961 6432 1995
rect 6466 1961 6500 1995
rect 6534 1961 6568 1995
rect 6602 1961 6636 1995
rect 6670 1961 6704 1995
rect 6738 1961 6772 1995
rect 6806 1961 6840 1995
rect 6874 1961 6908 1995
rect 6942 1961 6976 1995
rect 7010 1961 7044 1995
rect 7078 1961 7112 1995
rect 7146 1961 7180 1995
rect 7214 1961 7248 1995
rect 7282 1961 7316 1995
rect 7350 1961 7384 1995
rect 7418 1961 7452 1995
rect 7486 1961 7520 1995
rect 7554 1961 7588 1995
rect 7622 1961 7656 1995
rect 7690 1961 7724 1995
rect 7758 1961 7792 1995
rect 7826 1961 7860 1995
rect 7894 1961 7928 1995
rect 7962 1961 7996 1995
rect 8030 1961 8064 1995
rect 8098 1961 8132 1995
rect 8166 1961 8200 1995
rect 8234 1961 8268 1995
rect 8302 1961 8336 1995
rect 8370 1961 8404 1995
rect 8438 1961 8472 1995
rect 8506 1961 8540 1995
rect 8574 1961 8608 1995
rect 8642 1961 8676 1995
rect 8710 1961 8744 1995
rect 8778 1961 8812 1995
rect 8846 1961 8880 1995
rect 8914 1961 8948 1995
rect 8982 1961 9016 1995
rect 9050 1961 9084 1995
rect 9118 1961 9152 1995
rect 9186 1961 9220 1995
rect 9254 1961 9288 1995
rect 9322 1961 9356 1995
rect 9390 1961 9424 1995
rect 9458 1961 9492 1995
rect 9526 1961 9560 1995
rect 9594 1961 9628 1995
rect 9662 1961 9696 1995
rect 9730 1961 9764 1995
rect 9798 1961 9832 1995
rect 9866 1961 9900 1995
rect 9934 1961 9968 1995
rect 10002 1961 10036 1995
rect 10070 1961 10104 1995
rect 10138 1961 10172 1995
rect 10206 1961 10240 1995
rect 10274 1961 10308 1995
rect 10342 1961 10376 1995
rect 10410 1961 10444 1995
rect 10478 1961 10512 1995
rect 10546 1961 10580 1995
rect 10614 1961 10648 1995
rect 10682 1961 10716 1995
rect 10750 1961 10784 1995
rect 10818 1961 10852 1995
rect 10886 1961 10920 1995
rect 10954 1961 10988 1995
rect 11022 1961 11056 1995
rect 11090 1961 11124 1995
rect 11158 1961 11192 1995
rect 11226 1961 11260 1995
rect 11294 1961 11328 1995
rect 11362 1961 11396 1995
rect 11430 1961 11464 1995
rect 11498 1961 11532 1995
rect 11566 1961 11600 1995
rect 11634 1961 11668 1995
rect 11702 1961 11736 1995
rect 11770 1961 11804 1995
rect 11838 1961 11872 1995
rect 11906 1961 11940 1995
rect 11974 1961 12008 1995
rect 12042 1961 12076 1995
rect 12110 1961 12144 1995
rect 12178 1961 12212 1995
rect 12246 1961 12280 1995
rect 12314 1961 12348 1995
rect 12382 1961 12416 1995
rect 12450 1961 12484 1995
rect 12518 1961 12552 1995
rect 12586 1961 12620 1995
rect 12654 1961 12688 1995
rect 12722 1961 12756 1995
rect 12790 1961 12824 1995
rect 12858 1961 12892 1995
rect 12926 1961 12960 1995
rect 12994 1961 13028 1995
rect 13062 1961 13096 1995
rect 13130 1961 13164 1995
rect 13198 1961 13232 1995
rect 13266 1961 13300 1995
rect 13334 1961 13368 1995
rect 13402 1961 13436 1995
rect 13470 1961 13504 1995
rect 13538 1961 13572 1995
rect 13606 1961 13640 1995
rect 13674 1961 13708 1995
rect 13742 1961 13776 1995
rect 13810 1961 13844 1995
rect 13878 1961 13912 1995
rect 13946 1961 13980 1995
rect 14014 1961 14048 1995
rect 14082 1961 14116 1995
rect 14150 1961 14184 1995
rect 14218 1961 14252 1995
rect 14286 1961 14320 1995
rect 14354 1961 14388 1995
rect 14422 1961 14456 1995
rect 14490 1961 14524 1995
rect 14558 1961 14592 1995
rect 14626 1961 14660 1995
rect 14694 1961 14728 1995
rect 14762 1961 14796 1995
rect 14830 1961 14864 1995
rect 14898 1961 14932 1995
rect 14966 1961 15000 1995
rect 15034 1961 15068 1995
rect 15102 1961 15136 1995
rect 15170 1961 15204 1995
rect 15238 1961 15272 1995
rect 15306 1961 15340 1995
rect 15374 1961 15408 1995
rect 15442 1961 15476 1995
rect 15510 1961 15544 1995
rect 15578 1961 15612 1995
rect 15646 1961 15680 1995
rect 15714 1961 15748 1995
rect 15782 1961 15816 1995
rect 15850 1961 15884 1995
rect 15918 1961 15952 1995
rect 15986 1961 16020 1995
rect 16054 1961 16088 1995
rect 16122 1961 16156 1995
rect 16190 1961 16224 1995
rect 16258 1961 16292 1995
rect 16326 1961 16360 1995
rect 16394 1961 16428 1995
rect 16462 1961 16496 1995
rect 16530 1961 16564 1995
rect 16598 1961 16632 1995
rect 16666 1961 16700 1995
rect 16734 1961 16768 1995
rect 16802 1961 16836 1995
rect 16870 1961 16904 1995
rect 16938 1961 16972 1995
rect 17006 1961 17040 1995
rect 17074 1961 17108 1995
rect 17142 1961 17176 1995
rect 17210 1961 17244 1995
rect 17278 1961 17312 1995
rect 17346 1961 17380 1995
rect 17414 1961 17448 1995
rect 17482 1961 17516 1995
rect 17550 1961 17584 1995
rect 17618 1961 17652 1995
rect 17686 1961 17720 1995
rect 17754 1961 17788 1995
rect 17822 1961 17856 1995
rect 17890 1961 17924 1995
rect 17958 1961 17992 1995
rect 18026 1961 18060 1995
rect 18094 1961 18128 1995
rect 18162 1961 18196 1995
rect 18230 1961 18264 1995
rect 18298 1961 18332 1995
rect 18366 1961 18400 1995
rect 18434 1961 18468 1995
rect 18502 1961 18536 1995
rect 18570 1961 18604 1995
rect 18638 1961 18672 1995
rect 18706 1961 18740 1995
rect 18774 1961 18808 1995
rect 18842 1961 18876 1995
rect 18910 1961 18944 1995
rect 18978 1961 19012 1995
rect 19046 1961 19080 1995
rect 19114 1961 19148 1995
rect 19182 1961 19216 1995
rect 19250 1961 19284 1995
rect 19318 1961 19352 1995
rect 19386 1961 19420 1995
rect 19454 1961 19488 1995
rect 19522 1961 19556 1995
rect 19590 1961 19624 1995
rect 19658 1961 19692 1995
rect 19726 1961 19760 1995
rect 19794 1961 19828 1995
rect 19862 1961 19896 1995
rect 19930 1961 19964 1995
rect 19998 1961 20032 1995
rect 20066 1961 20100 1995
rect 20134 1961 20168 1995
rect 20202 1961 20236 1995
rect 20270 1961 20304 1995
rect 20338 1961 20372 1995
rect 20406 1961 20440 1995
rect 20474 1961 20508 1995
rect 20542 1961 20576 1995
rect 20610 1961 20644 1995
rect 20678 1961 20712 1995
rect 20746 1961 20780 1995
rect 20814 1961 20848 1995
rect 20882 1961 20916 1995
rect 20950 1961 20984 1995
rect 21018 1961 21052 1995
rect 21086 1961 21120 1995
rect 21154 1961 21188 1995
rect 21222 1961 21256 1995
rect 21290 1961 21324 1995
rect 21358 1961 21392 1995
rect 21426 1961 21460 1995
rect 21494 1961 21528 1995
rect 21562 1961 21596 1995
rect 21630 1961 21664 1995
rect 21698 1961 21732 1995
rect 21766 1961 21800 1995
rect 21834 1961 21868 1995
rect 21902 1961 21936 1995
rect 21970 1961 22004 1995
rect 22038 1961 22072 1995
rect 22106 1961 22140 1995
rect 22174 1961 22208 1995
rect 22242 1961 22276 1995
rect 22310 1961 22344 1995
rect 22378 1961 22412 1995
rect 22446 1961 22480 1995
rect 22514 1961 22548 1995
rect 22582 1961 22616 1995
rect 22650 1961 22684 1995
rect 22718 1961 22752 1995
rect 22786 1961 22820 1995
rect 22854 1961 22888 1995
rect 22922 1961 22956 1995
rect 22990 1961 23024 1995
rect 23058 1961 23092 1995
rect 23126 1961 23160 1995
rect 23194 1961 23228 1995
rect 23262 1961 23296 1995
rect 23330 1961 23364 1995
rect 23398 1961 23432 1995
rect 23466 1961 23500 1995
rect 23534 1961 23568 1995
rect 23602 1961 23636 1995
rect 23670 1961 23704 1995
rect 23738 1961 23772 1995
rect 23806 1961 23840 1995
rect 23874 1961 23908 1995
rect 23942 1961 23976 1995
rect 24010 1961 24044 1995
rect 24078 1961 24112 1995
rect 24146 1961 24180 1995
rect 24214 1961 24248 1995
rect 24282 1961 24316 1995
rect 24350 1961 24384 1995
rect 24418 1961 24452 1995
rect 24486 1961 24520 1995
rect 24554 1961 24588 1995
rect 24622 1961 24656 1995
rect 24690 1961 24724 1995
rect 24758 1961 24792 1995
rect 24826 1961 24860 1995
rect 24894 1961 24928 1995
rect 24962 1961 24996 1995
rect 25030 1961 25064 1995
rect 25098 1961 25132 1995
rect 25166 1961 25200 1995
rect 25234 1961 25268 1995
rect 25302 1961 25336 1995
rect 25370 1961 25404 1995
rect 25438 1961 25472 1995
rect 25506 1961 25540 1995
rect 25574 1961 25608 1995
rect 25642 1961 25676 1995
rect 25710 1961 25744 1995
rect 25778 1961 25812 1995
rect 25846 1961 25880 1995
rect 25914 1961 25948 1995
rect 25982 1961 26016 1995
rect 26050 1961 26084 1995
rect 26118 1961 26152 1995
rect 26186 1961 26220 1995
rect 26254 1961 26288 1995
rect 26322 1961 26356 1995
rect 26390 1961 26424 1995
rect 26458 1961 26492 1995
rect 26526 1961 26560 1995
rect 26594 1961 26628 1995
rect 26662 1961 26696 1995
rect 26730 1961 26764 1995
rect 26798 1961 26832 1995
rect 26866 1961 26900 1995
rect 26934 1961 26968 1995
rect 27002 1961 27036 1995
rect 27070 1961 27104 1995
rect 27138 1961 27172 1995
rect 27206 1961 27240 1995
rect 27274 1961 27308 1995
rect 27342 1961 27376 1995
rect 27410 1961 27444 1995
rect 27478 1990 27512 1995
rect 27546 1991 27580 2024
rect 27614 1991 27648 2025
rect 27546 1990 27682 1991
rect 27478 1961 27682 1990
rect 1975 1956 27682 1961
rect 1975 1955 27580 1956
rect 1975 1921 27512 1955
rect 27546 1922 27580 1955
rect 27614 1922 27648 1956
rect 27546 1921 27682 1922
rect 1975 1887 2009 1921
rect 2043 1887 2078 1921
rect 2112 1887 2147 1921
rect 2181 1887 2216 1921
rect 2250 1887 2284 1921
rect 2318 1887 2352 1921
rect 2386 1887 2420 1921
rect 2454 1887 2488 1921
rect 2522 1887 2556 1921
rect 2590 1887 2624 1921
rect 2658 1887 2692 1921
rect 2726 1887 2760 1921
rect 2794 1887 2828 1921
rect 2862 1887 2896 1921
rect 2930 1887 2964 1921
rect 2998 1887 3032 1921
rect 3066 1887 3100 1921
rect 3134 1887 3168 1921
rect 3202 1887 3236 1921
rect 3270 1887 3304 1921
rect 3338 1887 3372 1921
rect 3406 1887 3440 1921
rect 3474 1887 3508 1921
rect 3542 1887 3576 1921
rect 3610 1887 3644 1921
rect 3678 1887 3712 1921
rect 3746 1887 3780 1921
rect 3814 1887 3848 1921
rect 3882 1887 3916 1921
rect 3950 1887 3984 1921
rect 4018 1887 4052 1921
rect 4086 1887 4120 1921
rect 4154 1887 4188 1921
rect 4222 1887 4256 1921
rect 4290 1887 4324 1921
rect 4358 1887 4392 1921
rect 4426 1887 4460 1921
rect 4494 1887 4528 1921
rect 4562 1887 4596 1921
rect 4630 1887 4664 1921
rect 4698 1887 4732 1921
rect 4766 1887 4800 1921
rect 4834 1887 4868 1921
rect 4902 1887 4936 1921
rect 4970 1887 5004 1921
rect 5038 1887 5072 1921
rect 5106 1887 5140 1921
rect 5174 1887 5208 1921
rect 5242 1887 5276 1921
rect 5310 1887 5344 1921
rect 5378 1887 5412 1921
rect 5446 1887 5480 1921
rect 5514 1887 5548 1921
rect 5582 1887 5616 1921
rect 5650 1887 5684 1921
rect 5718 1887 5752 1921
rect 5786 1887 5820 1921
rect 5854 1887 5888 1921
rect 5922 1887 5956 1921
rect 5990 1887 6024 1921
rect 6058 1887 6092 1921
rect 6126 1887 6160 1921
rect 6194 1887 6228 1921
rect 6262 1887 6296 1921
rect 6330 1887 6364 1921
rect 6398 1887 6432 1921
rect 6466 1887 6500 1921
rect 6534 1887 6568 1921
rect 6602 1887 6636 1921
rect 6670 1887 6704 1921
rect 6738 1887 6772 1921
rect 6806 1887 6840 1921
rect 6874 1887 6908 1921
rect 6942 1887 6976 1921
rect 7010 1887 7044 1921
rect 7078 1887 7112 1921
rect 7146 1887 7180 1921
rect 7214 1887 7248 1921
rect 7282 1887 7316 1921
rect 7350 1887 7384 1921
rect 7418 1887 7452 1921
rect 7486 1887 7520 1921
rect 7554 1887 7588 1921
rect 7622 1887 7656 1921
rect 7690 1887 7724 1921
rect 7758 1887 7792 1921
rect 7826 1887 7860 1921
rect 7894 1887 7928 1921
rect 7962 1887 7996 1921
rect 8030 1887 8064 1921
rect 8098 1887 8132 1921
rect 8166 1887 8200 1921
rect 8234 1887 8268 1921
rect 8302 1887 8336 1921
rect 8370 1887 8404 1921
rect 8438 1887 8472 1921
rect 8506 1887 8540 1921
rect 8574 1887 8608 1921
rect 8642 1887 8676 1921
rect 8710 1887 8744 1921
rect 8778 1887 8812 1921
rect 8846 1887 8880 1921
rect 8914 1887 8948 1921
rect 8982 1887 9016 1921
rect 9050 1887 9084 1921
rect 9118 1887 9152 1921
rect 9186 1887 9220 1921
rect 9254 1887 9288 1921
rect 9322 1887 9356 1921
rect 9390 1887 9424 1921
rect 9458 1887 9492 1921
rect 9526 1887 9560 1921
rect 9594 1887 9628 1921
rect 9662 1887 9696 1921
rect 9730 1887 9764 1921
rect 9798 1887 9832 1921
rect 9866 1887 9900 1921
rect 9934 1887 9968 1921
rect 10002 1887 10036 1921
rect 10070 1887 10104 1921
rect 10138 1887 10172 1921
rect 10206 1887 10240 1921
rect 10274 1887 10308 1921
rect 10342 1887 10376 1921
rect 10410 1887 10444 1921
rect 10478 1887 10512 1921
rect 10546 1887 10580 1921
rect 10614 1887 10648 1921
rect 10682 1887 10716 1921
rect 10750 1887 10784 1921
rect 10818 1887 10852 1921
rect 10886 1887 10920 1921
rect 10954 1887 10988 1921
rect 11022 1887 11056 1921
rect 11090 1887 11124 1921
rect 11158 1887 11192 1921
rect 11226 1887 11260 1921
rect 11294 1887 11328 1921
rect 11362 1887 11396 1921
rect 11430 1887 11464 1921
rect 11498 1887 11532 1921
rect 11566 1887 11600 1921
rect 11634 1887 11668 1921
rect 11702 1887 11736 1921
rect 11770 1887 11804 1921
rect 11838 1887 11872 1921
rect 11906 1887 11940 1921
rect 11974 1887 12008 1921
rect 12042 1887 12076 1921
rect 12110 1887 12144 1921
rect 12178 1887 12212 1921
rect 12246 1887 12280 1921
rect 12314 1887 12348 1921
rect 12382 1887 12416 1921
rect 12450 1887 12484 1921
rect 12518 1887 12552 1921
rect 12586 1887 12620 1921
rect 12654 1887 12688 1921
rect 12722 1887 12756 1921
rect 12790 1887 12824 1921
rect 12858 1887 12892 1921
rect 12926 1887 12960 1921
rect 12994 1887 13028 1921
rect 13062 1887 13096 1921
rect 13130 1887 13164 1921
rect 13198 1887 13232 1921
rect 13266 1887 13300 1921
rect 13334 1887 13368 1921
rect 13402 1887 13436 1921
rect 13470 1887 13504 1921
rect 13538 1887 13572 1921
rect 13606 1887 13640 1921
rect 13674 1887 13708 1921
rect 13742 1887 13776 1921
rect 13810 1887 13844 1921
rect 13878 1887 13912 1921
rect 13946 1887 13980 1921
rect 14014 1887 14048 1921
rect 14082 1887 14116 1921
rect 14150 1887 14184 1921
rect 14218 1887 14252 1921
rect 14286 1887 14320 1921
rect 14354 1887 14388 1921
rect 14422 1887 14456 1921
rect 14490 1887 14524 1921
rect 14558 1887 14592 1921
rect 14626 1887 14660 1921
rect 14694 1887 14728 1921
rect 14762 1887 14796 1921
rect 14830 1887 14864 1921
rect 14898 1887 14932 1921
rect 14966 1887 15000 1921
rect 15034 1887 15068 1921
rect 15102 1887 15136 1921
rect 15170 1887 15204 1921
rect 15238 1887 15272 1921
rect 15306 1887 15340 1921
rect 15374 1887 15408 1921
rect 15442 1887 15476 1921
rect 15510 1887 15544 1921
rect 15578 1887 15612 1921
rect 15646 1887 15680 1921
rect 15714 1887 15748 1921
rect 15782 1887 15816 1921
rect 15850 1887 15884 1921
rect 15918 1887 15952 1921
rect 15986 1887 16020 1921
rect 16054 1887 16088 1921
rect 16122 1887 16156 1921
rect 16190 1887 16224 1921
rect 16258 1887 16292 1921
rect 16326 1887 16360 1921
rect 16394 1887 16428 1921
rect 16462 1887 16496 1921
rect 16530 1887 16564 1921
rect 16598 1887 16632 1921
rect 16666 1887 16700 1921
rect 16734 1887 16768 1921
rect 16802 1887 16836 1921
rect 16870 1887 16904 1921
rect 16938 1887 16972 1921
rect 17006 1887 17040 1921
rect 17074 1887 17108 1921
rect 17142 1887 17176 1921
rect 17210 1887 17244 1921
rect 17278 1887 17312 1921
rect 17346 1887 17380 1921
rect 17414 1887 17448 1921
rect 17482 1887 17516 1921
rect 17550 1887 17584 1921
rect 17618 1887 17652 1921
rect 17686 1887 17720 1921
rect 17754 1887 17788 1921
rect 17822 1887 17856 1921
rect 17890 1887 17924 1921
rect 17958 1887 17992 1921
rect 18026 1887 18060 1921
rect 18094 1887 18128 1921
rect 18162 1887 18196 1921
rect 18230 1887 18264 1921
rect 18298 1887 18332 1921
rect 18366 1887 18400 1921
rect 18434 1887 18468 1921
rect 18502 1887 18536 1921
rect 18570 1887 18604 1921
rect 18638 1887 18672 1921
rect 18706 1887 18740 1921
rect 18774 1887 18808 1921
rect 18842 1887 18876 1921
rect 18910 1887 18944 1921
rect 18978 1887 19012 1921
rect 19046 1887 19080 1921
rect 19114 1887 19148 1921
rect 19182 1887 19216 1921
rect 19250 1887 19284 1921
rect 19318 1887 19352 1921
rect 19386 1887 19420 1921
rect 19454 1887 19488 1921
rect 19522 1887 19556 1921
rect 19590 1887 19624 1921
rect 19658 1887 19692 1921
rect 19726 1887 19760 1921
rect 19794 1887 19828 1921
rect 19862 1887 19896 1921
rect 19930 1887 19964 1921
rect 19998 1887 20032 1921
rect 20066 1887 20100 1921
rect 20134 1887 20168 1921
rect 20202 1887 20236 1921
rect 20270 1887 20304 1921
rect 20338 1887 20372 1921
rect 20406 1887 20440 1921
rect 20474 1887 20508 1921
rect 20542 1887 20576 1921
rect 20610 1887 20644 1921
rect 20678 1887 20712 1921
rect 20746 1887 20780 1921
rect 20814 1887 20848 1921
rect 20882 1887 20916 1921
rect 20950 1887 20984 1921
rect 21018 1887 21052 1921
rect 21086 1887 21120 1921
rect 21154 1887 21188 1921
rect 21222 1887 21256 1921
rect 21290 1887 21324 1921
rect 21358 1887 21392 1921
rect 21426 1887 21460 1921
rect 21494 1887 21528 1921
rect 21562 1887 21596 1921
rect 21630 1887 21664 1921
rect 21698 1887 21732 1921
rect 21766 1887 21800 1921
rect 21834 1887 21868 1921
rect 21902 1887 21936 1921
rect 21970 1887 22004 1921
rect 22038 1887 22072 1921
rect 22106 1887 22140 1921
rect 22174 1887 22208 1921
rect 22242 1887 22276 1921
rect 22310 1887 22344 1921
rect 22378 1887 22412 1921
rect 22446 1887 22480 1921
rect 22514 1887 22548 1921
rect 22582 1887 22616 1921
rect 22650 1887 22684 1921
rect 22718 1887 22752 1921
rect 22786 1887 22820 1921
rect 22854 1887 22888 1921
rect 22922 1887 22956 1921
rect 22990 1887 23024 1921
rect 23058 1887 23092 1921
rect 23126 1887 23160 1921
rect 23194 1887 23228 1921
rect 23262 1887 23296 1921
rect 23330 1887 23364 1921
rect 23398 1887 23432 1921
rect 23466 1887 23500 1921
rect 23534 1887 23568 1921
rect 23602 1887 23636 1921
rect 23670 1887 23704 1921
rect 23738 1887 23772 1921
rect 23806 1887 23840 1921
rect 23874 1887 23908 1921
rect 23942 1887 23976 1921
rect 24010 1887 24044 1921
rect 24078 1887 24112 1921
rect 24146 1887 24180 1921
rect 24214 1887 24248 1921
rect 24282 1887 24316 1921
rect 24350 1887 24384 1921
rect 24418 1887 24452 1921
rect 24486 1887 24520 1921
rect 24554 1887 24588 1921
rect 24622 1887 24656 1921
rect 24690 1887 24724 1921
rect 24758 1887 24792 1921
rect 24826 1887 24860 1921
rect 24894 1887 24928 1921
rect 24962 1887 24996 1921
rect 25030 1887 25064 1921
rect 25098 1887 25132 1921
rect 25166 1887 25200 1921
rect 25234 1887 25268 1921
rect 25302 1887 25336 1921
rect 25370 1887 25404 1921
rect 25438 1887 25472 1921
rect 25506 1887 25540 1921
rect 25574 1887 25608 1921
rect 25642 1887 25676 1921
rect 25710 1887 25744 1921
rect 25778 1887 25812 1921
rect 25846 1887 25880 1921
rect 25914 1887 25948 1921
rect 25982 1887 26016 1921
rect 26050 1887 26084 1921
rect 26118 1887 26152 1921
rect 26186 1887 26220 1921
rect 26254 1887 26288 1921
rect 26322 1887 26356 1921
rect 26390 1887 26424 1921
rect 26458 1887 26492 1921
rect 26526 1887 26560 1921
rect 26594 1887 26628 1921
rect 26662 1887 26696 1921
rect 26730 1887 26764 1921
rect 26798 1887 26832 1921
rect 26866 1887 26900 1921
rect 26934 1887 26968 1921
rect 27002 1887 27036 1921
rect 27070 1887 27104 1921
rect 27138 1887 27172 1921
rect 27206 1887 27240 1921
rect 27274 1887 27308 1921
rect 27342 1887 27376 1921
rect 27410 1887 27444 1921
rect 27478 1887 27682 1921
rect 1975 1886 27580 1887
rect 1975 1852 27512 1886
rect 27546 1853 27580 1886
rect 27614 1853 27648 1887
rect 27546 1852 27682 1853
rect 1975 1847 27682 1852
rect 1975 1813 2009 1847
rect 2043 1813 2078 1847
rect 2112 1813 2147 1847
rect 2181 1813 2216 1847
rect 2250 1813 2284 1847
rect 2318 1813 2352 1847
rect 2386 1813 2420 1847
rect 2454 1813 2488 1847
rect 2522 1813 2556 1847
rect 2590 1813 2624 1847
rect 2658 1813 2692 1847
rect 2726 1813 2760 1847
rect 2794 1813 2828 1847
rect 2862 1813 2896 1847
rect 2930 1813 2964 1847
rect 2998 1813 3032 1847
rect 3066 1813 3100 1847
rect 3134 1813 3168 1847
rect 3202 1813 3236 1847
rect 3270 1813 3304 1847
rect 3338 1813 3372 1847
rect 3406 1813 3440 1847
rect 3474 1813 3508 1847
rect 3542 1813 3576 1847
rect 3610 1813 3644 1847
rect 3678 1813 3712 1847
rect 3746 1813 3780 1847
rect 3814 1813 3848 1847
rect 3882 1813 3916 1847
rect 3950 1813 3984 1847
rect 4018 1813 4052 1847
rect 4086 1813 4120 1847
rect 4154 1813 4188 1847
rect 4222 1813 4256 1847
rect 4290 1813 4324 1847
rect 4358 1813 4392 1847
rect 4426 1813 4460 1847
rect 4494 1813 4528 1847
rect 4562 1813 4596 1847
rect 4630 1813 4664 1847
rect 4698 1813 4732 1847
rect 4766 1813 4800 1847
rect 4834 1813 4868 1847
rect 4902 1813 4936 1847
rect 4970 1813 5004 1847
rect 5038 1813 5072 1847
rect 5106 1813 5140 1847
rect 5174 1813 5208 1847
rect 5242 1813 5276 1847
rect 5310 1813 5344 1847
rect 5378 1813 5412 1847
rect 5446 1813 5480 1847
rect 5514 1813 5548 1847
rect 5582 1813 5616 1847
rect 5650 1813 5684 1847
rect 5718 1813 5752 1847
rect 5786 1813 5820 1847
rect 5854 1813 5888 1847
rect 5922 1813 5956 1847
rect 5990 1813 6024 1847
rect 6058 1813 6092 1847
rect 6126 1813 6160 1847
rect 6194 1813 6228 1847
rect 6262 1813 6296 1847
rect 6330 1813 6364 1847
rect 6398 1813 6432 1847
rect 6466 1813 6500 1847
rect 6534 1813 6568 1847
rect 6602 1813 6636 1847
rect 6670 1813 6704 1847
rect 6738 1813 6772 1847
rect 6806 1813 6840 1847
rect 6874 1813 6908 1847
rect 6942 1813 6976 1847
rect 7010 1813 7044 1847
rect 7078 1813 7112 1847
rect 7146 1813 7180 1847
rect 7214 1813 7248 1847
rect 7282 1813 7316 1847
rect 7350 1813 7384 1847
rect 7418 1813 7452 1847
rect 7486 1813 7520 1847
rect 7554 1813 7588 1847
rect 7622 1813 7656 1847
rect 7690 1813 7724 1847
rect 7758 1813 7792 1847
rect 7826 1813 7860 1847
rect 7894 1813 7928 1847
rect 7962 1813 7996 1847
rect 8030 1813 8064 1847
rect 8098 1813 8132 1847
rect 8166 1813 8200 1847
rect 8234 1813 8268 1847
rect 8302 1813 8336 1847
rect 8370 1813 8404 1847
rect 8438 1813 8472 1847
rect 8506 1813 8540 1847
rect 8574 1813 8608 1847
rect 8642 1813 8676 1847
rect 8710 1813 8744 1847
rect 8778 1813 8812 1847
rect 8846 1813 8880 1847
rect 8914 1813 8948 1847
rect 8982 1813 9016 1847
rect 9050 1813 9084 1847
rect 9118 1813 9152 1847
rect 9186 1813 9220 1847
rect 9254 1813 9288 1847
rect 9322 1813 9356 1847
rect 9390 1813 9424 1847
rect 9458 1813 9492 1847
rect 9526 1813 9560 1847
rect 9594 1813 9628 1847
rect 9662 1813 9696 1847
rect 9730 1813 9764 1847
rect 9798 1813 9832 1847
rect 9866 1813 9900 1847
rect 9934 1813 9968 1847
rect 10002 1813 10036 1847
rect 10070 1813 10104 1847
rect 10138 1813 10172 1847
rect 10206 1813 10240 1847
rect 10274 1813 10308 1847
rect 10342 1813 10376 1847
rect 10410 1813 10444 1847
rect 10478 1813 10512 1847
rect 10546 1813 10580 1847
rect 10614 1813 10648 1847
rect 10682 1813 10716 1847
rect 10750 1813 10784 1847
rect 10818 1813 10852 1847
rect 10886 1813 10920 1847
rect 10954 1813 10988 1847
rect 11022 1813 11056 1847
rect 11090 1813 11124 1847
rect 11158 1813 11192 1847
rect 11226 1813 11260 1847
rect 11294 1813 11328 1847
rect 11362 1813 11396 1847
rect 11430 1813 11464 1847
rect 11498 1813 11532 1847
rect 11566 1813 11600 1847
rect 11634 1813 11668 1847
rect 11702 1813 11736 1847
rect 11770 1813 11804 1847
rect 11838 1813 11872 1847
rect 11906 1813 11940 1847
rect 11974 1813 12008 1847
rect 12042 1813 12076 1847
rect 12110 1813 12144 1847
rect 12178 1813 12212 1847
rect 12246 1813 12280 1847
rect 12314 1813 12348 1847
rect 12382 1813 12416 1847
rect 12450 1813 12484 1847
rect 12518 1813 12552 1847
rect 12586 1813 12620 1847
rect 12654 1813 12688 1847
rect 12722 1813 12756 1847
rect 12790 1813 12824 1847
rect 12858 1813 12892 1847
rect 12926 1813 12960 1847
rect 12994 1813 13028 1847
rect 13062 1813 13096 1847
rect 13130 1813 13164 1847
rect 13198 1813 13232 1847
rect 13266 1813 13300 1847
rect 13334 1813 13368 1847
rect 13402 1813 13436 1847
rect 13470 1813 13504 1847
rect 13538 1813 13572 1847
rect 13606 1813 13640 1847
rect 13674 1813 13708 1847
rect 13742 1813 13776 1847
rect 13810 1813 13844 1847
rect 13878 1813 13912 1847
rect 13946 1813 13980 1847
rect 14014 1813 14048 1847
rect 14082 1813 14116 1847
rect 14150 1813 14184 1847
rect 14218 1813 14252 1847
rect 14286 1813 14320 1847
rect 14354 1813 14388 1847
rect 14422 1813 14456 1847
rect 14490 1813 14524 1847
rect 14558 1813 14592 1847
rect 14626 1813 14660 1847
rect 14694 1813 14728 1847
rect 14762 1813 14796 1847
rect 14830 1813 14864 1847
rect 14898 1813 14932 1847
rect 14966 1813 15000 1847
rect 15034 1813 15068 1847
rect 15102 1813 15136 1847
rect 15170 1813 15204 1847
rect 15238 1813 15272 1847
rect 15306 1813 15340 1847
rect 15374 1813 15408 1847
rect 15442 1813 15476 1847
rect 15510 1813 15544 1847
rect 15578 1813 15612 1847
rect 15646 1813 15680 1847
rect 15714 1813 15748 1847
rect 15782 1813 15816 1847
rect 15850 1813 15884 1847
rect 15918 1813 15952 1847
rect 15986 1813 16020 1847
rect 16054 1813 16088 1847
rect 16122 1813 16156 1847
rect 16190 1813 16224 1847
rect 16258 1813 16292 1847
rect 16326 1813 16360 1847
rect 16394 1813 16428 1847
rect 16462 1813 16496 1847
rect 16530 1813 16564 1847
rect 16598 1813 16632 1847
rect 16666 1813 16700 1847
rect 16734 1813 16768 1847
rect 16802 1813 16836 1847
rect 16870 1813 16904 1847
rect 16938 1813 16972 1847
rect 17006 1813 17040 1847
rect 17074 1813 17108 1847
rect 17142 1813 17176 1847
rect 17210 1813 17244 1847
rect 17278 1813 17312 1847
rect 17346 1813 17380 1847
rect 17414 1813 17448 1847
rect 17482 1813 17516 1847
rect 17550 1813 17584 1847
rect 17618 1813 17652 1847
rect 17686 1813 17720 1847
rect 17754 1813 17788 1847
rect 17822 1813 17856 1847
rect 17890 1813 17924 1847
rect 17958 1813 17992 1847
rect 18026 1813 18060 1847
rect 18094 1813 18128 1847
rect 18162 1813 18196 1847
rect 18230 1813 18264 1847
rect 18298 1813 18332 1847
rect 18366 1813 18400 1847
rect 18434 1813 18468 1847
rect 18502 1813 18536 1847
rect 18570 1813 18604 1847
rect 18638 1813 18672 1847
rect 18706 1813 18740 1847
rect 18774 1813 18808 1847
rect 18842 1813 18876 1847
rect 18910 1813 18944 1847
rect 18978 1813 19012 1847
rect 19046 1813 19080 1847
rect 19114 1813 19148 1847
rect 19182 1813 19216 1847
rect 19250 1813 19284 1847
rect 19318 1813 19352 1847
rect 19386 1813 19420 1847
rect 19454 1813 19488 1847
rect 19522 1813 19556 1847
rect 19590 1813 19624 1847
rect 19658 1813 19692 1847
rect 19726 1813 19760 1847
rect 19794 1813 19828 1847
rect 19862 1813 19896 1847
rect 19930 1813 19964 1847
rect 19998 1813 20032 1847
rect 20066 1813 20100 1847
rect 20134 1813 20168 1847
rect 20202 1813 20236 1847
rect 20270 1813 20304 1847
rect 20338 1813 20372 1847
rect 20406 1813 20440 1847
rect 20474 1813 20508 1847
rect 20542 1813 20576 1847
rect 20610 1813 20644 1847
rect 20678 1813 20712 1847
rect 20746 1813 20780 1847
rect 20814 1813 20848 1847
rect 20882 1813 20916 1847
rect 20950 1813 20984 1847
rect 21018 1813 21052 1847
rect 21086 1813 21120 1847
rect 21154 1813 21188 1847
rect 21222 1813 21256 1847
rect 21290 1813 21324 1847
rect 21358 1813 21392 1847
rect 21426 1813 21460 1847
rect 21494 1813 21528 1847
rect 21562 1813 21596 1847
rect 21630 1813 21664 1847
rect 21698 1813 21732 1847
rect 21766 1813 21800 1847
rect 21834 1813 21868 1847
rect 21902 1813 21936 1847
rect 21970 1813 22004 1847
rect 22038 1813 22072 1847
rect 22106 1813 22140 1847
rect 22174 1813 22208 1847
rect 22242 1813 22276 1847
rect 22310 1813 22344 1847
rect 22378 1813 22412 1847
rect 22446 1813 22480 1847
rect 22514 1813 22548 1847
rect 22582 1813 22616 1847
rect 22650 1813 22684 1847
rect 22718 1813 22752 1847
rect 22786 1813 22820 1847
rect 22854 1813 22888 1847
rect 22922 1813 22956 1847
rect 22990 1813 23024 1847
rect 23058 1813 23092 1847
rect 23126 1813 23160 1847
rect 23194 1813 23228 1847
rect 23262 1813 23296 1847
rect 23330 1813 23364 1847
rect 23398 1813 23432 1847
rect 23466 1813 23500 1847
rect 23534 1813 23568 1847
rect 23602 1813 23636 1847
rect 23670 1813 23704 1847
rect 23738 1813 23772 1847
rect 23806 1813 23840 1847
rect 23874 1813 23908 1847
rect 23942 1813 23976 1847
rect 24010 1813 24044 1847
rect 24078 1813 24112 1847
rect 24146 1813 24180 1847
rect 24214 1813 24248 1847
rect 24282 1813 24316 1847
rect 24350 1813 24384 1847
rect 24418 1813 24452 1847
rect 24486 1813 24520 1847
rect 24554 1813 24588 1847
rect 24622 1813 24656 1847
rect 24690 1813 24724 1847
rect 24758 1813 24792 1847
rect 24826 1813 24860 1847
rect 24894 1813 24928 1847
rect 24962 1813 24996 1847
rect 25030 1813 25064 1847
rect 25098 1813 25132 1847
rect 25166 1813 25200 1847
rect 25234 1813 25268 1847
rect 25302 1813 25336 1847
rect 25370 1813 25404 1847
rect 25438 1813 25472 1847
rect 25506 1813 25540 1847
rect 25574 1813 25608 1847
rect 25642 1813 25676 1847
rect 25710 1813 25744 1847
rect 25778 1813 25812 1847
rect 25846 1813 25880 1847
rect 25914 1813 25948 1847
rect 25982 1813 26016 1847
rect 26050 1813 26084 1847
rect 26118 1813 26152 1847
rect 26186 1813 26220 1847
rect 26254 1813 26288 1847
rect 26322 1813 26356 1847
rect 26390 1813 26424 1847
rect 26458 1813 26492 1847
rect 26526 1813 26560 1847
rect 26594 1813 26628 1847
rect 26662 1813 26696 1847
rect 26730 1813 26764 1847
rect 26798 1813 26832 1847
rect 26866 1813 26900 1847
rect 26934 1813 26968 1847
rect 27002 1813 27036 1847
rect 27070 1813 27104 1847
rect 27138 1813 27172 1847
rect 27206 1813 27240 1847
rect 27274 1813 27308 1847
rect 27342 1813 27376 1847
rect 27410 1813 27444 1847
rect 27478 1818 27682 1847
rect 27478 1817 27580 1818
rect 27478 1813 27512 1817
rect 1975 1783 27512 1813
rect 27546 1784 27580 1817
rect 27614 1784 27648 1818
rect 27546 1783 27682 1784
rect 1975 1773 27682 1783
rect 1975 1739 2009 1773
rect 2043 1739 2078 1773
rect 2112 1739 2147 1773
rect 2181 1739 2216 1773
rect 2250 1739 2284 1773
rect 2318 1739 2352 1773
rect 2386 1739 2420 1773
rect 2454 1739 2488 1773
rect 2522 1739 2556 1773
rect 2590 1739 2624 1773
rect 2658 1739 2692 1773
rect 2726 1739 2760 1773
rect 2794 1739 2828 1773
rect 2862 1739 2896 1773
rect 2930 1739 2964 1773
rect 2998 1739 3032 1773
rect 3066 1739 3100 1773
rect 3134 1739 3168 1773
rect 3202 1739 3236 1773
rect 3270 1739 3304 1773
rect 3338 1739 3372 1773
rect 3406 1739 3440 1773
rect 3474 1739 3508 1773
rect 3542 1739 3576 1773
rect 3610 1739 3644 1773
rect 3678 1739 3712 1773
rect 3746 1739 3780 1773
rect 3814 1739 3848 1773
rect 3882 1739 3916 1773
rect 3950 1739 3984 1773
rect 4018 1739 4052 1773
rect 4086 1739 4120 1773
rect 4154 1739 4188 1773
rect 4222 1739 4256 1773
rect 4290 1739 4324 1773
rect 4358 1739 4392 1773
rect 4426 1739 4460 1773
rect 4494 1739 4528 1773
rect 4562 1739 4596 1773
rect 4630 1739 4664 1773
rect 4698 1739 4732 1773
rect 4766 1739 4800 1773
rect 4834 1739 4868 1773
rect 4902 1739 4936 1773
rect 4970 1739 5004 1773
rect 5038 1739 5072 1773
rect 5106 1739 5140 1773
rect 5174 1739 5208 1773
rect 5242 1739 5276 1773
rect 5310 1739 5344 1773
rect 5378 1739 5412 1773
rect 5446 1739 5480 1773
rect 5514 1739 5548 1773
rect 5582 1739 5616 1773
rect 5650 1739 5684 1773
rect 5718 1739 5752 1773
rect 5786 1739 5820 1773
rect 5854 1739 5888 1773
rect 5922 1739 5956 1773
rect 5990 1739 6024 1773
rect 6058 1739 6092 1773
rect 6126 1739 6160 1773
rect 6194 1739 6228 1773
rect 6262 1739 6296 1773
rect 6330 1739 6364 1773
rect 6398 1739 6432 1773
rect 6466 1739 6500 1773
rect 6534 1739 6568 1773
rect 6602 1739 6636 1773
rect 6670 1739 6704 1773
rect 6738 1739 6772 1773
rect 6806 1739 6840 1773
rect 6874 1739 6908 1773
rect 6942 1739 6976 1773
rect 7010 1739 7044 1773
rect 7078 1739 7112 1773
rect 7146 1739 7180 1773
rect 7214 1739 7248 1773
rect 7282 1739 7316 1773
rect 7350 1739 7384 1773
rect 7418 1739 7452 1773
rect 7486 1739 7520 1773
rect 7554 1739 7588 1773
rect 7622 1739 7656 1773
rect 7690 1739 7724 1773
rect 7758 1739 7792 1773
rect 7826 1739 7860 1773
rect 7894 1739 7928 1773
rect 7962 1739 7996 1773
rect 8030 1739 8064 1773
rect 8098 1739 8132 1773
rect 8166 1739 8200 1773
rect 8234 1739 8268 1773
rect 8302 1739 8336 1773
rect 8370 1739 8404 1773
rect 8438 1739 8472 1773
rect 8506 1739 8540 1773
rect 8574 1739 8608 1773
rect 8642 1739 8676 1773
rect 8710 1739 8744 1773
rect 8778 1739 8812 1773
rect 8846 1739 8880 1773
rect 8914 1739 8948 1773
rect 8982 1739 9016 1773
rect 9050 1739 9084 1773
rect 9118 1739 9152 1773
rect 9186 1739 9220 1773
rect 9254 1739 9288 1773
rect 9322 1739 9356 1773
rect 9390 1739 9424 1773
rect 9458 1739 9492 1773
rect 9526 1739 9560 1773
rect 9594 1739 9628 1773
rect 9662 1739 9696 1773
rect 9730 1739 9764 1773
rect 9798 1739 9832 1773
rect 9866 1739 9900 1773
rect 9934 1739 9968 1773
rect 10002 1739 10036 1773
rect 10070 1739 10104 1773
rect 10138 1739 10172 1773
rect 10206 1739 10240 1773
rect 10274 1739 10308 1773
rect 10342 1739 10376 1773
rect 10410 1739 10444 1773
rect 10478 1739 10512 1773
rect 10546 1739 10580 1773
rect 10614 1739 10648 1773
rect 10682 1739 10716 1773
rect 10750 1739 10784 1773
rect 10818 1739 10852 1773
rect 10886 1739 10920 1773
rect 10954 1739 10988 1773
rect 11022 1739 11056 1773
rect 11090 1739 11124 1773
rect 11158 1739 11192 1773
rect 11226 1739 11260 1773
rect 11294 1739 11328 1773
rect 11362 1739 11396 1773
rect 11430 1739 11464 1773
rect 11498 1739 11532 1773
rect 11566 1739 11600 1773
rect 11634 1739 11668 1773
rect 11702 1739 11736 1773
rect 11770 1739 11804 1773
rect 11838 1739 11872 1773
rect 11906 1739 11940 1773
rect 11974 1739 12008 1773
rect 12042 1739 12076 1773
rect 12110 1739 12144 1773
rect 12178 1739 12212 1773
rect 12246 1739 12280 1773
rect 12314 1739 12348 1773
rect 12382 1739 12416 1773
rect 12450 1739 12484 1773
rect 12518 1739 12552 1773
rect 12586 1739 12620 1773
rect 12654 1739 12688 1773
rect 12722 1739 12756 1773
rect 12790 1739 12824 1773
rect 12858 1739 12892 1773
rect 12926 1739 12960 1773
rect 12994 1739 13028 1773
rect 13062 1739 13096 1773
rect 13130 1739 13164 1773
rect 13198 1739 13232 1773
rect 13266 1739 13300 1773
rect 13334 1739 13368 1773
rect 13402 1739 13436 1773
rect 13470 1739 13504 1773
rect 13538 1739 13572 1773
rect 13606 1739 13640 1773
rect 13674 1739 13708 1773
rect 13742 1739 13776 1773
rect 13810 1739 13844 1773
rect 13878 1739 13912 1773
rect 13946 1739 13980 1773
rect 14014 1739 14048 1773
rect 14082 1739 14116 1773
rect 14150 1739 14184 1773
rect 14218 1739 14252 1773
rect 14286 1739 14320 1773
rect 14354 1739 14388 1773
rect 14422 1739 14456 1773
rect 14490 1739 14524 1773
rect 14558 1739 14592 1773
rect 14626 1739 14660 1773
rect 14694 1739 14728 1773
rect 14762 1739 14796 1773
rect 14830 1739 14864 1773
rect 14898 1739 14932 1773
rect 14966 1739 15000 1773
rect 15034 1739 15068 1773
rect 15102 1739 15136 1773
rect 15170 1739 15204 1773
rect 15238 1739 15272 1773
rect 15306 1739 15340 1773
rect 15374 1739 15408 1773
rect 15442 1739 15476 1773
rect 15510 1739 15544 1773
rect 15578 1739 15612 1773
rect 15646 1739 15680 1773
rect 15714 1739 15748 1773
rect 15782 1739 15816 1773
rect 15850 1739 15884 1773
rect 15918 1739 15952 1773
rect 15986 1739 16020 1773
rect 16054 1739 16088 1773
rect 16122 1739 16156 1773
rect 16190 1739 16224 1773
rect 16258 1739 16292 1773
rect 16326 1739 16360 1773
rect 16394 1739 16428 1773
rect 16462 1739 16496 1773
rect 16530 1739 16564 1773
rect 16598 1739 16632 1773
rect 16666 1739 16700 1773
rect 16734 1739 16768 1773
rect 16802 1739 16836 1773
rect 16870 1739 16904 1773
rect 16938 1739 16972 1773
rect 17006 1739 17040 1773
rect 17074 1739 17108 1773
rect 17142 1739 17176 1773
rect 17210 1739 17244 1773
rect 17278 1739 17312 1773
rect 17346 1739 17380 1773
rect 17414 1739 17448 1773
rect 17482 1739 17516 1773
rect 17550 1739 17584 1773
rect 17618 1739 17652 1773
rect 17686 1739 17720 1773
rect 17754 1739 17788 1773
rect 17822 1739 17856 1773
rect 17890 1739 17924 1773
rect 17958 1739 17992 1773
rect 18026 1739 18060 1773
rect 18094 1739 18128 1773
rect 18162 1739 18196 1773
rect 18230 1739 18264 1773
rect 18298 1739 18332 1773
rect 18366 1739 18400 1773
rect 18434 1739 18468 1773
rect 18502 1739 18536 1773
rect 18570 1739 18604 1773
rect 18638 1739 18672 1773
rect 18706 1739 18740 1773
rect 18774 1739 18808 1773
rect 18842 1739 18876 1773
rect 18910 1739 18944 1773
rect 18978 1739 19012 1773
rect 19046 1739 19080 1773
rect 19114 1739 19148 1773
rect 19182 1739 19216 1773
rect 19250 1739 19284 1773
rect 19318 1739 19352 1773
rect 19386 1739 19420 1773
rect 19454 1739 19488 1773
rect 19522 1739 19556 1773
rect 19590 1739 19624 1773
rect 19658 1739 19692 1773
rect 19726 1739 19760 1773
rect 19794 1739 19828 1773
rect 19862 1739 19896 1773
rect 19930 1739 19964 1773
rect 19998 1739 20032 1773
rect 20066 1739 20100 1773
rect 20134 1739 20168 1773
rect 20202 1739 20236 1773
rect 20270 1739 20304 1773
rect 20338 1739 20372 1773
rect 20406 1739 20440 1773
rect 20474 1739 20508 1773
rect 20542 1739 20576 1773
rect 20610 1739 20644 1773
rect 20678 1739 20712 1773
rect 20746 1739 20780 1773
rect 20814 1739 20848 1773
rect 20882 1739 20916 1773
rect 20950 1739 20984 1773
rect 21018 1739 21052 1773
rect 21086 1739 21120 1773
rect 21154 1739 21188 1773
rect 21222 1739 21256 1773
rect 21290 1739 21324 1773
rect 21358 1739 21392 1773
rect 21426 1739 21460 1773
rect 21494 1739 21528 1773
rect 21562 1739 21596 1773
rect 21630 1739 21664 1773
rect 21698 1739 21732 1773
rect 21766 1739 21800 1773
rect 21834 1739 21868 1773
rect 21902 1739 21936 1773
rect 21970 1739 22004 1773
rect 22038 1739 22072 1773
rect 22106 1739 22140 1773
rect 22174 1739 22208 1773
rect 22242 1739 22276 1773
rect 22310 1739 22344 1773
rect 22378 1739 22412 1773
rect 22446 1739 22480 1773
rect 22514 1739 22548 1773
rect 22582 1739 22616 1773
rect 22650 1739 22684 1773
rect 22718 1739 22752 1773
rect 22786 1739 22820 1773
rect 22854 1739 22888 1773
rect 22922 1739 22956 1773
rect 22990 1739 23024 1773
rect 23058 1739 23092 1773
rect 23126 1739 23160 1773
rect 23194 1739 23228 1773
rect 23262 1739 23296 1773
rect 23330 1739 23364 1773
rect 23398 1739 23432 1773
rect 23466 1739 23500 1773
rect 23534 1739 23568 1773
rect 23602 1739 23636 1773
rect 23670 1739 23704 1773
rect 23738 1739 23772 1773
rect 23806 1739 23840 1773
rect 23874 1739 23908 1773
rect 23942 1739 23976 1773
rect 24010 1739 24044 1773
rect 24078 1739 24112 1773
rect 24146 1739 24180 1773
rect 24214 1739 24248 1773
rect 24282 1739 24316 1773
rect 24350 1739 24384 1773
rect 24418 1739 24452 1773
rect 24486 1739 24520 1773
rect 24554 1739 24588 1773
rect 24622 1739 24656 1773
rect 24690 1739 24724 1773
rect 24758 1739 24792 1773
rect 24826 1739 24860 1773
rect 24894 1739 24928 1773
rect 24962 1739 24996 1773
rect 25030 1739 25064 1773
rect 25098 1739 25132 1773
rect 25166 1739 25200 1773
rect 25234 1739 25268 1773
rect 25302 1739 25336 1773
rect 25370 1739 25404 1773
rect 25438 1739 25472 1773
rect 25506 1739 25540 1773
rect 25574 1739 25608 1773
rect 25642 1739 25676 1773
rect 25710 1739 25744 1773
rect 25778 1739 25812 1773
rect 25846 1739 25880 1773
rect 25914 1739 25948 1773
rect 25982 1739 26016 1773
rect 26050 1739 26084 1773
rect 26118 1739 26152 1773
rect 26186 1739 26220 1773
rect 26254 1739 26288 1773
rect 26322 1739 26356 1773
rect 26390 1739 26424 1773
rect 26458 1739 26492 1773
rect 26526 1739 26560 1773
rect 26594 1739 26628 1773
rect 26662 1739 26696 1773
rect 26730 1739 26764 1773
rect 26798 1739 26832 1773
rect 26866 1739 26900 1773
rect 26934 1739 26968 1773
rect 27002 1739 27036 1773
rect 27070 1739 27104 1773
rect 27138 1739 27172 1773
rect 27206 1739 27240 1773
rect 27274 1739 27308 1773
rect 27342 1739 27376 1773
rect 27410 1739 27444 1773
rect 27478 1749 27682 1773
rect 27478 1748 27580 1749
rect 27478 1739 27512 1748
rect 1975 1714 27512 1739
rect 27546 1715 27580 1748
rect 27614 1715 27648 1749
rect 27546 1714 27682 1715
rect 1975 1699 27682 1714
rect 1975 1665 2009 1699
rect 2043 1665 2078 1699
rect 2112 1665 2147 1699
rect 2181 1665 2216 1699
rect 2250 1665 2284 1699
rect 2318 1665 2352 1699
rect 2386 1665 2420 1699
rect 2454 1665 2488 1699
rect 2522 1665 2556 1699
rect 2590 1665 2624 1699
rect 2658 1665 2692 1699
rect 2726 1665 2760 1699
rect 2794 1665 2828 1699
rect 2862 1665 2896 1699
rect 2930 1665 2964 1699
rect 2998 1665 3032 1699
rect 3066 1665 3100 1699
rect 3134 1665 3168 1699
rect 3202 1665 3236 1699
rect 3270 1665 3304 1699
rect 3338 1665 3372 1699
rect 3406 1665 3440 1699
rect 3474 1665 3508 1699
rect 3542 1665 3576 1699
rect 3610 1665 3644 1699
rect 3678 1665 3712 1699
rect 3746 1665 3780 1699
rect 3814 1665 3848 1699
rect 3882 1665 3916 1699
rect 3950 1665 3984 1699
rect 4018 1665 4052 1699
rect 4086 1665 4120 1699
rect 4154 1665 4188 1699
rect 4222 1665 4256 1699
rect 4290 1665 4324 1699
rect 4358 1665 4392 1699
rect 4426 1665 4460 1699
rect 4494 1665 4528 1699
rect 4562 1665 4596 1699
rect 4630 1665 4664 1699
rect 4698 1665 4732 1699
rect 4766 1665 4800 1699
rect 4834 1665 4868 1699
rect 4902 1665 4936 1699
rect 4970 1665 5004 1699
rect 5038 1665 5072 1699
rect 5106 1665 5140 1699
rect 5174 1665 5208 1699
rect 5242 1665 5276 1699
rect 5310 1665 5344 1699
rect 5378 1665 5412 1699
rect 5446 1665 5480 1699
rect 5514 1665 5548 1699
rect 5582 1665 5616 1699
rect 5650 1665 5684 1699
rect 5718 1665 5752 1699
rect 5786 1665 5820 1699
rect 5854 1665 5888 1699
rect 5922 1665 5956 1699
rect 5990 1665 6024 1699
rect 6058 1665 6092 1699
rect 6126 1665 6160 1699
rect 6194 1665 6228 1699
rect 6262 1665 6296 1699
rect 6330 1665 6364 1699
rect 6398 1665 6432 1699
rect 6466 1665 6500 1699
rect 6534 1665 6568 1699
rect 6602 1665 6636 1699
rect 6670 1665 6704 1699
rect 6738 1665 6772 1699
rect 6806 1665 6840 1699
rect 6874 1665 6908 1699
rect 6942 1665 6976 1699
rect 7010 1665 7044 1699
rect 7078 1665 7112 1699
rect 7146 1665 7180 1699
rect 7214 1665 7248 1699
rect 7282 1665 7316 1699
rect 7350 1665 7384 1699
rect 7418 1665 7452 1699
rect 7486 1665 7520 1699
rect 7554 1665 7588 1699
rect 7622 1665 7656 1699
rect 7690 1665 7724 1699
rect 7758 1665 7792 1699
rect 7826 1665 7860 1699
rect 7894 1665 7928 1699
rect 7962 1665 7996 1699
rect 8030 1665 8064 1699
rect 8098 1665 8132 1699
rect 8166 1665 8200 1699
rect 8234 1665 8268 1699
rect 8302 1665 8336 1699
rect 8370 1665 8404 1699
rect 8438 1665 8472 1699
rect 8506 1665 8540 1699
rect 8574 1665 8608 1699
rect 8642 1665 8676 1699
rect 8710 1665 8744 1699
rect 8778 1665 8812 1699
rect 8846 1665 8880 1699
rect 8914 1665 8948 1699
rect 8982 1665 9016 1699
rect 9050 1665 9084 1699
rect 9118 1665 9152 1699
rect 9186 1665 9220 1699
rect 9254 1665 9288 1699
rect 9322 1665 9356 1699
rect 9390 1665 9424 1699
rect 9458 1665 9492 1699
rect 9526 1665 9560 1699
rect 9594 1665 9628 1699
rect 9662 1665 9696 1699
rect 9730 1665 9764 1699
rect 9798 1665 9832 1699
rect 9866 1665 9900 1699
rect 9934 1665 9968 1699
rect 10002 1665 10036 1699
rect 10070 1665 10104 1699
rect 10138 1665 10172 1699
rect 10206 1665 10240 1699
rect 10274 1665 10308 1699
rect 10342 1665 10376 1699
rect 10410 1665 10444 1699
rect 10478 1665 10512 1699
rect 10546 1665 10580 1699
rect 10614 1665 10648 1699
rect 10682 1665 10716 1699
rect 10750 1665 10784 1699
rect 10818 1665 10852 1699
rect 10886 1665 10920 1699
rect 10954 1665 10988 1699
rect 11022 1665 11056 1699
rect 11090 1665 11124 1699
rect 11158 1665 11192 1699
rect 11226 1665 11260 1699
rect 11294 1665 11328 1699
rect 11362 1665 11396 1699
rect 11430 1665 11464 1699
rect 11498 1665 11532 1699
rect 11566 1665 11600 1699
rect 11634 1665 11668 1699
rect 11702 1665 11736 1699
rect 11770 1665 11804 1699
rect 11838 1665 11872 1699
rect 11906 1665 11940 1699
rect 11974 1665 12008 1699
rect 12042 1665 12076 1699
rect 12110 1665 12144 1699
rect 12178 1665 12212 1699
rect 12246 1665 12280 1699
rect 12314 1665 12348 1699
rect 12382 1665 12416 1699
rect 12450 1665 12484 1699
rect 12518 1665 12552 1699
rect 12586 1665 12620 1699
rect 12654 1665 12688 1699
rect 12722 1665 12756 1699
rect 12790 1665 12824 1699
rect 12858 1665 12892 1699
rect 12926 1665 12960 1699
rect 12994 1665 13028 1699
rect 13062 1665 13096 1699
rect 13130 1665 13164 1699
rect 13198 1665 13232 1699
rect 13266 1665 13300 1699
rect 13334 1665 13368 1699
rect 13402 1665 13436 1699
rect 13470 1665 13504 1699
rect 13538 1665 13572 1699
rect 13606 1665 13640 1699
rect 13674 1665 13708 1699
rect 13742 1665 13776 1699
rect 13810 1665 13844 1699
rect 13878 1665 13912 1699
rect 13946 1665 13980 1699
rect 14014 1665 14048 1699
rect 14082 1665 14116 1699
rect 14150 1665 14184 1699
rect 14218 1665 14252 1699
rect 14286 1665 14320 1699
rect 14354 1665 14388 1699
rect 14422 1665 14456 1699
rect 14490 1665 14524 1699
rect 14558 1665 14592 1699
rect 14626 1665 14660 1699
rect 14694 1665 14728 1699
rect 14762 1665 14796 1699
rect 14830 1665 14864 1699
rect 14898 1665 14932 1699
rect 14966 1665 15000 1699
rect 15034 1665 15068 1699
rect 15102 1665 15136 1699
rect 15170 1665 15204 1699
rect 15238 1665 15272 1699
rect 15306 1665 15340 1699
rect 15374 1665 15408 1699
rect 15442 1665 15476 1699
rect 15510 1665 15544 1699
rect 15578 1665 15612 1699
rect 15646 1665 15680 1699
rect 15714 1665 15748 1699
rect 15782 1665 15816 1699
rect 15850 1665 15884 1699
rect 15918 1665 15952 1699
rect 15986 1665 16020 1699
rect 16054 1665 16088 1699
rect 16122 1665 16156 1699
rect 16190 1665 16224 1699
rect 16258 1665 16292 1699
rect 16326 1665 16360 1699
rect 16394 1665 16428 1699
rect 16462 1665 16496 1699
rect 16530 1665 16564 1699
rect 16598 1665 16632 1699
rect 16666 1665 16700 1699
rect 16734 1665 16768 1699
rect 16802 1665 16836 1699
rect 16870 1665 16904 1699
rect 16938 1665 16972 1699
rect 17006 1665 17040 1699
rect 17074 1665 17108 1699
rect 17142 1665 17176 1699
rect 17210 1665 17244 1699
rect 17278 1665 17312 1699
rect 17346 1665 17380 1699
rect 17414 1665 17448 1699
rect 17482 1665 17516 1699
rect 17550 1665 17584 1699
rect 17618 1665 17652 1699
rect 17686 1665 17720 1699
rect 17754 1665 17788 1699
rect 17822 1665 17856 1699
rect 17890 1665 17924 1699
rect 17958 1665 17992 1699
rect 18026 1665 18060 1699
rect 18094 1665 18128 1699
rect 18162 1665 18196 1699
rect 18230 1665 18264 1699
rect 18298 1665 18332 1699
rect 18366 1665 18400 1699
rect 18434 1665 18468 1699
rect 18502 1665 18536 1699
rect 18570 1665 18604 1699
rect 18638 1665 18672 1699
rect 18706 1665 18740 1699
rect 18774 1665 18808 1699
rect 18842 1665 18876 1699
rect 18910 1665 18944 1699
rect 18978 1665 19012 1699
rect 19046 1665 19080 1699
rect 19114 1665 19148 1699
rect 19182 1665 19216 1699
rect 19250 1665 19284 1699
rect 19318 1665 19352 1699
rect 19386 1665 19420 1699
rect 19454 1665 19488 1699
rect 19522 1665 19556 1699
rect 19590 1665 19624 1699
rect 19658 1665 19692 1699
rect 19726 1665 19760 1699
rect 19794 1665 19828 1699
rect 19862 1665 19896 1699
rect 19930 1665 19964 1699
rect 19998 1665 20032 1699
rect 20066 1665 20100 1699
rect 20134 1665 20168 1699
rect 20202 1665 20236 1699
rect 20270 1665 20304 1699
rect 20338 1665 20372 1699
rect 20406 1665 20440 1699
rect 20474 1665 20508 1699
rect 20542 1665 20576 1699
rect 20610 1665 20644 1699
rect 20678 1665 20712 1699
rect 20746 1665 20780 1699
rect 20814 1665 20848 1699
rect 20882 1665 20916 1699
rect 20950 1665 20984 1699
rect 21018 1665 21052 1699
rect 21086 1665 21120 1699
rect 21154 1665 21188 1699
rect 21222 1665 21256 1699
rect 21290 1665 21324 1699
rect 21358 1665 21392 1699
rect 21426 1665 21460 1699
rect 21494 1665 21528 1699
rect 21562 1665 21596 1699
rect 21630 1665 21664 1699
rect 21698 1665 21732 1699
rect 21766 1665 21800 1699
rect 21834 1665 21868 1699
rect 21902 1665 21936 1699
rect 21970 1665 22004 1699
rect 22038 1665 22072 1699
rect 22106 1665 22140 1699
rect 22174 1665 22208 1699
rect 22242 1665 22276 1699
rect 22310 1665 22344 1699
rect 22378 1665 22412 1699
rect 22446 1665 22480 1699
rect 22514 1665 22548 1699
rect 22582 1665 22616 1699
rect 22650 1665 22684 1699
rect 22718 1665 22752 1699
rect 22786 1665 22820 1699
rect 22854 1665 22888 1699
rect 22922 1665 22956 1699
rect 22990 1665 23024 1699
rect 23058 1665 23092 1699
rect 23126 1665 23160 1699
rect 23194 1665 23228 1699
rect 23262 1665 23296 1699
rect 23330 1665 23364 1699
rect 23398 1665 23432 1699
rect 23466 1665 23500 1699
rect 23534 1665 23568 1699
rect 23602 1665 23636 1699
rect 23670 1665 23704 1699
rect 23738 1665 23772 1699
rect 23806 1665 23840 1699
rect 23874 1665 23908 1699
rect 23942 1665 23976 1699
rect 24010 1665 24044 1699
rect 24078 1665 24112 1699
rect 24146 1665 24180 1699
rect 24214 1665 24248 1699
rect 24282 1665 24316 1699
rect 24350 1665 24384 1699
rect 24418 1665 24452 1699
rect 24486 1665 24520 1699
rect 24554 1665 24588 1699
rect 24622 1665 24656 1699
rect 24690 1665 24724 1699
rect 24758 1665 24792 1699
rect 24826 1665 24860 1699
rect 24894 1665 24928 1699
rect 24962 1665 24996 1699
rect 25030 1665 25064 1699
rect 25098 1665 25132 1699
rect 25166 1665 25200 1699
rect 25234 1665 25268 1699
rect 25302 1665 25336 1699
rect 25370 1665 25404 1699
rect 25438 1665 25472 1699
rect 25506 1665 25540 1699
rect 25574 1665 25608 1699
rect 25642 1665 25676 1699
rect 25710 1665 25744 1699
rect 25778 1665 25812 1699
rect 25846 1665 25880 1699
rect 25914 1665 25948 1699
rect 25982 1665 26016 1699
rect 26050 1665 26084 1699
rect 26118 1665 26152 1699
rect 26186 1665 26220 1699
rect 26254 1665 26288 1699
rect 26322 1665 26356 1699
rect 26390 1665 26424 1699
rect 26458 1665 26492 1699
rect 26526 1665 26560 1699
rect 26594 1665 26628 1699
rect 26662 1665 26696 1699
rect 26730 1665 26764 1699
rect 26798 1665 26832 1699
rect 26866 1665 26900 1699
rect 26934 1665 26968 1699
rect 27002 1665 27036 1699
rect 27070 1665 27104 1699
rect 27138 1665 27172 1699
rect 27206 1665 27240 1699
rect 27274 1665 27308 1699
rect 27342 1665 27376 1699
rect 27410 1665 27444 1699
rect 27478 1680 27682 1699
rect 27478 1679 27580 1680
rect 27478 1665 27512 1679
rect 1975 1645 27512 1665
rect 27546 1646 27580 1679
rect 27614 1646 27648 1680
rect 27546 1645 27682 1646
rect 1975 1625 27682 1645
rect 1975 1591 2009 1625
rect 2043 1591 2078 1625
rect 2112 1591 2147 1625
rect 2181 1591 2216 1625
rect 2250 1591 2284 1625
rect 2318 1591 2352 1625
rect 2386 1591 2420 1625
rect 2454 1591 2488 1625
rect 2522 1591 2556 1625
rect 2590 1591 2624 1625
rect 2658 1591 2692 1625
rect 2726 1591 2760 1625
rect 2794 1591 2828 1625
rect 2862 1591 2896 1625
rect 2930 1591 2964 1625
rect 2998 1591 3032 1625
rect 3066 1591 3100 1625
rect 3134 1591 3168 1625
rect 3202 1591 3236 1625
rect 3270 1591 3304 1625
rect 3338 1591 3372 1625
rect 3406 1591 3440 1625
rect 3474 1591 3508 1625
rect 3542 1591 3576 1625
rect 3610 1591 3644 1625
rect 3678 1591 3712 1625
rect 3746 1591 3780 1625
rect 3814 1591 3848 1625
rect 3882 1591 3916 1625
rect 3950 1591 3984 1625
rect 4018 1591 4052 1625
rect 4086 1591 4120 1625
rect 4154 1591 4188 1625
rect 4222 1591 4256 1625
rect 4290 1591 4324 1625
rect 4358 1591 4392 1625
rect 4426 1591 4460 1625
rect 4494 1591 4528 1625
rect 4562 1591 4596 1625
rect 4630 1591 4664 1625
rect 4698 1591 4732 1625
rect 4766 1591 4800 1625
rect 4834 1591 4868 1625
rect 4902 1591 4936 1625
rect 4970 1591 5004 1625
rect 5038 1591 5072 1625
rect 5106 1591 5140 1625
rect 5174 1591 5208 1625
rect 5242 1591 5276 1625
rect 5310 1591 5344 1625
rect 5378 1591 5412 1625
rect 5446 1591 5480 1625
rect 5514 1591 5548 1625
rect 5582 1591 5616 1625
rect 5650 1591 5684 1625
rect 5718 1591 5752 1625
rect 5786 1591 5820 1625
rect 5854 1591 5888 1625
rect 5922 1591 5956 1625
rect 5990 1591 6024 1625
rect 6058 1591 6092 1625
rect 6126 1591 6160 1625
rect 6194 1591 6228 1625
rect 6262 1591 6296 1625
rect 6330 1591 6364 1625
rect 6398 1591 6432 1625
rect 6466 1591 6500 1625
rect 6534 1591 6568 1625
rect 6602 1591 6636 1625
rect 6670 1591 6704 1625
rect 6738 1591 6772 1625
rect 6806 1591 6840 1625
rect 6874 1591 6908 1625
rect 6942 1591 6976 1625
rect 7010 1591 7044 1625
rect 7078 1591 7112 1625
rect 7146 1591 7180 1625
rect 7214 1591 7248 1625
rect 7282 1591 7316 1625
rect 7350 1591 7384 1625
rect 7418 1591 7452 1625
rect 7486 1591 7520 1625
rect 7554 1591 7588 1625
rect 7622 1591 7656 1625
rect 7690 1591 7724 1625
rect 7758 1591 7792 1625
rect 7826 1591 7860 1625
rect 7894 1591 7928 1625
rect 7962 1591 7996 1625
rect 8030 1591 8064 1625
rect 8098 1591 8132 1625
rect 8166 1591 8200 1625
rect 8234 1591 8268 1625
rect 8302 1591 8336 1625
rect 8370 1591 8404 1625
rect 8438 1591 8472 1625
rect 8506 1591 8540 1625
rect 8574 1591 8608 1625
rect 8642 1591 8676 1625
rect 8710 1591 8744 1625
rect 8778 1591 8812 1625
rect 8846 1591 8880 1625
rect 8914 1591 8948 1625
rect 8982 1591 9016 1625
rect 9050 1591 9084 1625
rect 9118 1591 9152 1625
rect 9186 1591 9220 1625
rect 9254 1591 9288 1625
rect 9322 1591 9356 1625
rect 9390 1591 9424 1625
rect 9458 1591 9492 1625
rect 9526 1591 9560 1625
rect 9594 1591 9628 1625
rect 9662 1591 9696 1625
rect 9730 1591 9764 1625
rect 9798 1591 9832 1625
rect 9866 1591 9900 1625
rect 9934 1591 9968 1625
rect 10002 1591 10036 1625
rect 10070 1591 10104 1625
rect 10138 1591 10172 1625
rect 10206 1591 10240 1625
rect 10274 1591 10308 1625
rect 10342 1591 10376 1625
rect 10410 1591 10444 1625
rect 10478 1591 10512 1625
rect 10546 1591 10580 1625
rect 10614 1591 10648 1625
rect 10682 1591 10716 1625
rect 10750 1591 10784 1625
rect 10818 1591 10852 1625
rect 10886 1591 10920 1625
rect 10954 1591 10988 1625
rect 11022 1591 11056 1625
rect 11090 1591 11124 1625
rect 11158 1591 11192 1625
rect 11226 1591 11260 1625
rect 11294 1591 11328 1625
rect 11362 1591 11396 1625
rect 11430 1591 11464 1625
rect 11498 1591 11532 1625
rect 11566 1591 11600 1625
rect 11634 1591 11668 1625
rect 11702 1591 11736 1625
rect 11770 1591 11804 1625
rect 11838 1591 11872 1625
rect 11906 1591 11940 1625
rect 11974 1591 12008 1625
rect 12042 1591 12076 1625
rect 12110 1591 12144 1625
rect 12178 1591 12212 1625
rect 12246 1591 12280 1625
rect 12314 1591 12348 1625
rect 12382 1591 12416 1625
rect 12450 1591 12484 1625
rect 12518 1591 12552 1625
rect 12586 1591 12620 1625
rect 12654 1591 12688 1625
rect 12722 1591 12756 1625
rect 12790 1591 12824 1625
rect 12858 1591 12892 1625
rect 12926 1591 12960 1625
rect 12994 1591 13028 1625
rect 13062 1591 13096 1625
rect 13130 1591 13164 1625
rect 13198 1591 13232 1625
rect 13266 1591 13300 1625
rect 13334 1591 13368 1625
rect 13402 1591 13436 1625
rect 13470 1591 13504 1625
rect 13538 1591 13572 1625
rect 13606 1591 13640 1625
rect 13674 1591 13708 1625
rect 13742 1591 13776 1625
rect 13810 1591 13844 1625
rect 13878 1591 13912 1625
rect 13946 1591 13980 1625
rect 14014 1591 14048 1625
rect 14082 1591 14116 1625
rect 14150 1591 14184 1625
rect 14218 1591 14252 1625
rect 14286 1591 14320 1625
rect 14354 1591 14388 1625
rect 14422 1591 14456 1625
rect 14490 1591 14524 1625
rect 14558 1591 14592 1625
rect 14626 1591 14660 1625
rect 14694 1591 14728 1625
rect 14762 1591 14796 1625
rect 14830 1591 14864 1625
rect 14898 1591 14932 1625
rect 14966 1591 15000 1625
rect 15034 1591 15068 1625
rect 15102 1591 15136 1625
rect 15170 1591 15204 1625
rect 15238 1591 15272 1625
rect 15306 1591 15340 1625
rect 15374 1591 15408 1625
rect 15442 1591 15476 1625
rect 15510 1591 15544 1625
rect 15578 1591 15612 1625
rect 15646 1591 15680 1625
rect 15714 1591 15748 1625
rect 15782 1591 15816 1625
rect 15850 1591 15884 1625
rect 15918 1591 15952 1625
rect 15986 1591 16020 1625
rect 16054 1591 16088 1625
rect 16122 1591 16156 1625
rect 16190 1591 16224 1625
rect 16258 1591 16292 1625
rect 16326 1591 16360 1625
rect 16394 1591 16428 1625
rect 16462 1591 16496 1625
rect 16530 1591 16564 1625
rect 16598 1591 16632 1625
rect 16666 1591 16700 1625
rect 16734 1591 16768 1625
rect 16802 1591 16836 1625
rect 16870 1591 16904 1625
rect 16938 1591 16972 1625
rect 17006 1591 17040 1625
rect 17074 1591 17108 1625
rect 17142 1591 17176 1625
rect 17210 1591 17244 1625
rect 17278 1591 17312 1625
rect 17346 1591 17380 1625
rect 17414 1591 17448 1625
rect 17482 1591 17516 1625
rect 17550 1591 17584 1625
rect 17618 1591 17652 1625
rect 17686 1591 17720 1625
rect 17754 1591 17788 1625
rect 17822 1591 17856 1625
rect 17890 1591 17924 1625
rect 17958 1591 17992 1625
rect 18026 1591 18060 1625
rect 18094 1591 18128 1625
rect 18162 1591 18196 1625
rect 18230 1591 18264 1625
rect 18298 1591 18332 1625
rect 18366 1591 18400 1625
rect 18434 1591 18468 1625
rect 18502 1591 18536 1625
rect 18570 1591 18604 1625
rect 18638 1591 18672 1625
rect 18706 1591 18740 1625
rect 18774 1591 18808 1625
rect 18842 1591 18876 1625
rect 18910 1591 18944 1625
rect 18978 1591 19012 1625
rect 19046 1591 19080 1625
rect 19114 1591 19148 1625
rect 19182 1591 19216 1625
rect 19250 1591 19284 1625
rect 19318 1591 19352 1625
rect 19386 1591 19420 1625
rect 19454 1591 19488 1625
rect 19522 1591 19556 1625
rect 19590 1591 19624 1625
rect 19658 1591 19692 1625
rect 19726 1591 19760 1625
rect 19794 1591 19828 1625
rect 19862 1591 19896 1625
rect 19930 1591 19964 1625
rect 19998 1591 20032 1625
rect 20066 1591 20100 1625
rect 20134 1591 20168 1625
rect 20202 1591 20236 1625
rect 20270 1591 20304 1625
rect 20338 1591 20372 1625
rect 20406 1591 20440 1625
rect 20474 1591 20508 1625
rect 20542 1591 20576 1625
rect 20610 1591 20644 1625
rect 20678 1591 20712 1625
rect 20746 1591 20780 1625
rect 20814 1591 20848 1625
rect 20882 1591 20916 1625
rect 20950 1591 20984 1625
rect 21018 1591 21052 1625
rect 21086 1591 21120 1625
rect 21154 1591 21188 1625
rect 21222 1591 21256 1625
rect 21290 1591 21324 1625
rect 21358 1591 21392 1625
rect 21426 1591 21460 1625
rect 21494 1591 21528 1625
rect 21562 1591 21596 1625
rect 21630 1591 21664 1625
rect 21698 1591 21732 1625
rect 21766 1591 21800 1625
rect 21834 1591 21868 1625
rect 21902 1591 21936 1625
rect 21970 1591 22004 1625
rect 22038 1591 22072 1625
rect 22106 1591 22140 1625
rect 22174 1591 22208 1625
rect 22242 1591 22276 1625
rect 22310 1591 22344 1625
rect 22378 1591 22412 1625
rect 22446 1591 22480 1625
rect 22514 1591 22548 1625
rect 22582 1591 22616 1625
rect 22650 1591 22684 1625
rect 22718 1591 22752 1625
rect 22786 1591 22820 1625
rect 22854 1591 22888 1625
rect 22922 1591 22956 1625
rect 22990 1591 23024 1625
rect 23058 1591 23092 1625
rect 23126 1591 23160 1625
rect 23194 1591 23228 1625
rect 23262 1591 23296 1625
rect 23330 1591 23364 1625
rect 23398 1591 23432 1625
rect 23466 1591 23500 1625
rect 23534 1591 23568 1625
rect 23602 1591 23636 1625
rect 23670 1591 23704 1625
rect 23738 1591 23772 1625
rect 23806 1591 23840 1625
rect 23874 1591 23908 1625
rect 23942 1591 23976 1625
rect 24010 1591 24044 1625
rect 24078 1591 24112 1625
rect 24146 1591 24180 1625
rect 24214 1591 24248 1625
rect 24282 1591 24316 1625
rect 24350 1591 24384 1625
rect 24418 1591 24452 1625
rect 24486 1591 24520 1625
rect 24554 1591 24588 1625
rect 24622 1591 24656 1625
rect 24690 1591 24724 1625
rect 24758 1591 24792 1625
rect 24826 1591 24860 1625
rect 24894 1591 24928 1625
rect 24962 1591 24996 1625
rect 25030 1591 25064 1625
rect 25098 1591 25132 1625
rect 25166 1591 25200 1625
rect 25234 1591 25268 1625
rect 25302 1591 25336 1625
rect 25370 1591 25404 1625
rect 25438 1591 25472 1625
rect 25506 1591 25540 1625
rect 25574 1591 25608 1625
rect 25642 1591 25676 1625
rect 25710 1591 25744 1625
rect 25778 1591 25812 1625
rect 25846 1591 25880 1625
rect 25914 1591 25948 1625
rect 25982 1591 26016 1625
rect 26050 1591 26084 1625
rect 26118 1591 26152 1625
rect 26186 1591 26220 1625
rect 26254 1591 26288 1625
rect 26322 1591 26356 1625
rect 26390 1591 26424 1625
rect 26458 1591 26492 1625
rect 26526 1591 26560 1625
rect 26594 1591 26628 1625
rect 26662 1591 26696 1625
rect 26730 1591 26764 1625
rect 26798 1591 26832 1625
rect 26866 1591 26900 1625
rect 26934 1591 26968 1625
rect 27002 1591 27036 1625
rect 27070 1591 27104 1625
rect 27138 1591 27172 1625
rect 27206 1591 27240 1625
rect 27274 1591 27308 1625
rect 27342 1591 27376 1625
rect 27410 1591 27444 1625
rect 27478 1611 27682 1625
rect 27478 1610 27580 1611
rect 27478 1591 27512 1610
rect 1975 1576 27512 1591
rect 27546 1577 27580 1610
rect 27614 1577 27648 1611
rect 27546 1576 27682 1577
rect 1975 1551 27682 1576
rect 1975 1517 2009 1551
rect 2043 1517 2078 1551
rect 2112 1517 2147 1551
rect 2181 1517 2216 1551
rect 2250 1517 2284 1551
rect 2318 1517 2352 1551
rect 2386 1517 2420 1551
rect 2454 1517 2488 1551
rect 2522 1517 2556 1551
rect 2590 1517 2624 1551
rect 2658 1517 2692 1551
rect 2726 1517 2760 1551
rect 2794 1517 2828 1551
rect 2862 1517 2896 1551
rect 2930 1517 2964 1551
rect 2998 1517 3032 1551
rect 3066 1517 3100 1551
rect 3134 1517 3168 1551
rect 3202 1517 3236 1551
rect 3270 1517 3304 1551
rect 3338 1517 3372 1551
rect 3406 1517 3440 1551
rect 3474 1517 3508 1551
rect 3542 1517 3576 1551
rect 3610 1517 3644 1551
rect 3678 1517 3712 1551
rect 3746 1517 3780 1551
rect 3814 1517 3848 1551
rect 3882 1517 3916 1551
rect 3950 1517 3984 1551
rect 4018 1517 4052 1551
rect 4086 1517 4120 1551
rect 4154 1517 4188 1551
rect 4222 1517 4256 1551
rect 4290 1517 4324 1551
rect 4358 1517 4392 1551
rect 4426 1517 4460 1551
rect 4494 1517 4528 1551
rect 4562 1517 4596 1551
rect 4630 1517 4664 1551
rect 4698 1517 4732 1551
rect 4766 1517 4800 1551
rect 4834 1517 4868 1551
rect 4902 1517 4936 1551
rect 4970 1517 5004 1551
rect 5038 1517 5072 1551
rect 5106 1517 5140 1551
rect 5174 1517 5208 1551
rect 5242 1517 5276 1551
rect 5310 1517 5344 1551
rect 5378 1517 5412 1551
rect 5446 1517 5480 1551
rect 5514 1517 5548 1551
rect 5582 1517 5616 1551
rect 5650 1517 5684 1551
rect 5718 1517 5752 1551
rect 5786 1517 5820 1551
rect 5854 1517 5888 1551
rect 5922 1517 5956 1551
rect 5990 1517 6024 1551
rect 6058 1517 6092 1551
rect 6126 1517 6160 1551
rect 6194 1517 6228 1551
rect 6262 1517 6296 1551
rect 6330 1517 6364 1551
rect 6398 1517 6432 1551
rect 6466 1517 6500 1551
rect 6534 1517 6568 1551
rect 6602 1517 6636 1551
rect 6670 1517 6704 1551
rect 6738 1517 6772 1551
rect 6806 1517 6840 1551
rect 6874 1517 6908 1551
rect 6942 1517 6976 1551
rect 7010 1517 7044 1551
rect 7078 1517 7112 1551
rect 7146 1517 7180 1551
rect 7214 1517 7248 1551
rect 7282 1517 7316 1551
rect 7350 1517 7384 1551
rect 7418 1517 7452 1551
rect 7486 1517 7520 1551
rect 7554 1517 7588 1551
rect 7622 1517 7656 1551
rect 7690 1517 7724 1551
rect 7758 1517 7792 1551
rect 7826 1517 7860 1551
rect 7894 1517 7928 1551
rect 7962 1517 7996 1551
rect 8030 1517 8064 1551
rect 8098 1517 8132 1551
rect 8166 1517 8200 1551
rect 8234 1517 8268 1551
rect 8302 1517 8336 1551
rect 8370 1517 8404 1551
rect 8438 1517 8472 1551
rect 8506 1517 8540 1551
rect 8574 1517 8608 1551
rect 8642 1517 8676 1551
rect 8710 1517 8744 1551
rect 8778 1517 8812 1551
rect 8846 1517 8880 1551
rect 8914 1517 8948 1551
rect 8982 1517 9016 1551
rect 9050 1517 9084 1551
rect 9118 1517 9152 1551
rect 9186 1517 9220 1551
rect 9254 1517 9288 1551
rect 9322 1517 9356 1551
rect 9390 1517 9424 1551
rect 9458 1517 9492 1551
rect 9526 1517 9560 1551
rect 9594 1517 9628 1551
rect 9662 1517 9696 1551
rect 9730 1517 9764 1551
rect 9798 1517 9832 1551
rect 9866 1517 9900 1551
rect 9934 1517 9968 1551
rect 10002 1517 10036 1551
rect 10070 1517 10104 1551
rect 10138 1517 10172 1551
rect 10206 1517 10240 1551
rect 10274 1517 10308 1551
rect 10342 1517 10376 1551
rect 10410 1517 10444 1551
rect 10478 1517 10512 1551
rect 10546 1517 10580 1551
rect 10614 1517 10648 1551
rect 10682 1517 10716 1551
rect 10750 1517 10784 1551
rect 10818 1517 10852 1551
rect 10886 1517 10920 1551
rect 10954 1517 10988 1551
rect 11022 1517 11056 1551
rect 11090 1517 11124 1551
rect 11158 1517 11192 1551
rect 11226 1517 11260 1551
rect 11294 1517 11328 1551
rect 11362 1517 11396 1551
rect 11430 1517 11464 1551
rect 11498 1517 11532 1551
rect 11566 1517 11600 1551
rect 11634 1517 11668 1551
rect 11702 1517 11736 1551
rect 11770 1517 11804 1551
rect 11838 1517 11872 1551
rect 11906 1517 11940 1551
rect 11974 1517 12008 1551
rect 12042 1517 12076 1551
rect 12110 1517 12144 1551
rect 12178 1517 12212 1551
rect 12246 1517 12280 1551
rect 12314 1517 12348 1551
rect 12382 1517 12416 1551
rect 12450 1517 12484 1551
rect 12518 1517 12552 1551
rect 12586 1517 12620 1551
rect 12654 1517 12688 1551
rect 12722 1517 12756 1551
rect 12790 1517 12824 1551
rect 12858 1517 12892 1551
rect 12926 1517 12960 1551
rect 12994 1517 13028 1551
rect 13062 1517 13096 1551
rect 13130 1517 13164 1551
rect 13198 1517 13232 1551
rect 13266 1517 13300 1551
rect 13334 1517 13368 1551
rect 13402 1517 13436 1551
rect 13470 1517 13504 1551
rect 13538 1517 13572 1551
rect 13606 1517 13640 1551
rect 13674 1517 13708 1551
rect 13742 1517 13776 1551
rect 13810 1517 13844 1551
rect 13878 1517 13912 1551
rect 13946 1517 13980 1551
rect 14014 1517 14048 1551
rect 14082 1517 14116 1551
rect 14150 1517 14184 1551
rect 14218 1517 14252 1551
rect 14286 1517 14320 1551
rect 14354 1517 14388 1551
rect 14422 1517 14456 1551
rect 14490 1517 14524 1551
rect 14558 1517 14592 1551
rect 14626 1517 14660 1551
rect 14694 1517 14728 1551
rect 14762 1517 14796 1551
rect 14830 1517 14864 1551
rect 14898 1517 14932 1551
rect 14966 1517 15000 1551
rect 15034 1517 15068 1551
rect 15102 1517 15136 1551
rect 15170 1517 15204 1551
rect 15238 1517 15272 1551
rect 15306 1517 15340 1551
rect 15374 1517 15408 1551
rect 15442 1517 15476 1551
rect 15510 1517 15544 1551
rect 15578 1517 15612 1551
rect 15646 1517 15680 1551
rect 15714 1517 15748 1551
rect 15782 1517 15816 1551
rect 15850 1517 15884 1551
rect 15918 1517 15952 1551
rect 15986 1517 16020 1551
rect 16054 1517 16088 1551
rect 16122 1517 16156 1551
rect 16190 1517 16224 1551
rect 16258 1517 16292 1551
rect 16326 1517 16360 1551
rect 16394 1517 16428 1551
rect 16462 1517 16496 1551
rect 16530 1517 16564 1551
rect 16598 1517 16632 1551
rect 16666 1517 16700 1551
rect 16734 1517 16768 1551
rect 16802 1517 16836 1551
rect 16870 1517 16904 1551
rect 16938 1517 16972 1551
rect 17006 1517 17040 1551
rect 17074 1517 17108 1551
rect 17142 1517 17176 1551
rect 17210 1517 17244 1551
rect 17278 1517 17312 1551
rect 17346 1517 17380 1551
rect 17414 1517 17448 1551
rect 17482 1517 17516 1551
rect 17550 1517 17584 1551
rect 17618 1517 17652 1551
rect 17686 1517 17720 1551
rect 17754 1517 17788 1551
rect 17822 1517 17856 1551
rect 17890 1517 17924 1551
rect 17958 1517 17992 1551
rect 18026 1517 18060 1551
rect 18094 1517 18128 1551
rect 18162 1517 18196 1551
rect 18230 1517 18264 1551
rect 18298 1517 18332 1551
rect 18366 1517 18400 1551
rect 18434 1517 18468 1551
rect 18502 1517 18536 1551
rect 18570 1517 18604 1551
rect 18638 1517 18672 1551
rect 18706 1517 18740 1551
rect 18774 1517 18808 1551
rect 18842 1517 18876 1551
rect 18910 1517 18944 1551
rect 18978 1517 19012 1551
rect 19046 1517 19080 1551
rect 19114 1517 19148 1551
rect 19182 1517 19216 1551
rect 19250 1517 19284 1551
rect 19318 1517 19352 1551
rect 19386 1517 19420 1551
rect 19454 1517 19488 1551
rect 19522 1517 19556 1551
rect 19590 1517 19624 1551
rect 19658 1517 19692 1551
rect 19726 1517 19760 1551
rect 19794 1517 19828 1551
rect 19862 1517 19896 1551
rect 19930 1517 19964 1551
rect 19998 1517 20032 1551
rect 20066 1517 20100 1551
rect 20134 1517 20168 1551
rect 20202 1517 20236 1551
rect 20270 1517 20304 1551
rect 20338 1517 20372 1551
rect 20406 1517 20440 1551
rect 20474 1517 20508 1551
rect 20542 1517 20576 1551
rect 20610 1517 20644 1551
rect 20678 1517 20712 1551
rect 20746 1517 20780 1551
rect 20814 1517 20848 1551
rect 20882 1517 20916 1551
rect 20950 1517 20984 1551
rect 21018 1517 21052 1551
rect 21086 1517 21120 1551
rect 21154 1517 21188 1551
rect 21222 1517 21256 1551
rect 21290 1517 21324 1551
rect 21358 1517 21392 1551
rect 21426 1517 21460 1551
rect 21494 1517 21528 1551
rect 21562 1517 21596 1551
rect 21630 1517 21664 1551
rect 21698 1517 21732 1551
rect 21766 1517 21800 1551
rect 21834 1517 21868 1551
rect 21902 1517 21936 1551
rect 21970 1517 22004 1551
rect 22038 1517 22072 1551
rect 22106 1517 22140 1551
rect 22174 1517 22208 1551
rect 22242 1517 22276 1551
rect 22310 1517 22344 1551
rect 22378 1517 22412 1551
rect 22446 1517 22480 1551
rect 22514 1517 22548 1551
rect 22582 1517 22616 1551
rect 22650 1517 22684 1551
rect 22718 1517 22752 1551
rect 22786 1517 22820 1551
rect 22854 1517 22888 1551
rect 22922 1517 22956 1551
rect 22990 1517 23024 1551
rect 23058 1517 23092 1551
rect 23126 1517 23160 1551
rect 23194 1517 23228 1551
rect 23262 1517 23296 1551
rect 23330 1517 23364 1551
rect 23398 1517 23432 1551
rect 23466 1517 23500 1551
rect 23534 1517 23568 1551
rect 23602 1517 23636 1551
rect 23670 1517 23704 1551
rect 23738 1517 23772 1551
rect 23806 1517 23840 1551
rect 23874 1517 23908 1551
rect 23942 1517 23976 1551
rect 24010 1517 24044 1551
rect 24078 1517 24112 1551
rect 24146 1517 24180 1551
rect 24214 1517 24248 1551
rect 24282 1517 24316 1551
rect 24350 1517 24384 1551
rect 24418 1517 24452 1551
rect 24486 1517 24520 1551
rect 24554 1517 24588 1551
rect 24622 1517 24656 1551
rect 24690 1517 24724 1551
rect 24758 1517 24792 1551
rect 24826 1517 24860 1551
rect 24894 1517 24928 1551
rect 24962 1517 24996 1551
rect 25030 1517 25064 1551
rect 25098 1517 25132 1551
rect 25166 1517 25200 1551
rect 25234 1517 25268 1551
rect 25302 1517 25336 1551
rect 25370 1517 25404 1551
rect 25438 1517 25472 1551
rect 25506 1517 25540 1551
rect 25574 1517 25608 1551
rect 25642 1517 25676 1551
rect 25710 1517 25744 1551
rect 25778 1517 25812 1551
rect 25846 1517 25880 1551
rect 25914 1517 25948 1551
rect 25982 1517 26016 1551
rect 26050 1517 26084 1551
rect 26118 1517 26152 1551
rect 26186 1517 26220 1551
rect 26254 1517 26288 1551
rect 26322 1517 26356 1551
rect 26390 1517 26424 1551
rect 26458 1517 26492 1551
rect 26526 1517 26560 1551
rect 26594 1517 26628 1551
rect 26662 1517 26696 1551
rect 26730 1517 26764 1551
rect 26798 1517 26832 1551
rect 26866 1517 26900 1551
rect 26934 1517 26968 1551
rect 27002 1517 27036 1551
rect 27070 1517 27104 1551
rect 27138 1517 27172 1551
rect 27206 1517 27240 1551
rect 27274 1517 27308 1551
rect 27342 1517 27376 1551
rect 27410 1517 27444 1551
rect 27478 1542 27682 1551
rect 27478 1541 27580 1542
rect 27478 1517 27512 1541
rect 1975 1507 27512 1517
rect 27546 1508 27580 1541
rect 27614 1508 27648 1542
rect 27546 1507 27682 1508
rect 1975 1473 27682 1507
rect 1975 1472 27580 1473
rect 1975 1438 2010 1472
rect 2044 1438 2079 1472
rect 2113 1438 2148 1472
rect 1907 1404 2148 1438
rect 27546 1439 27580 1472
rect 27614 1439 27648 1473
rect 27546 1404 27682 1439
rect 1907 1370 1942 1404
rect 1976 1370 2011 1404
rect 2045 1370 2080 1404
rect 1805 1336 2080 1370
rect 1805 1302 1873 1336
rect 1907 1302 1942 1336
rect 1976 1302 2011 1336
rect 2045 1302 2080 1336
rect 27614 1370 27648 1404
rect 27614 1302 27682 1370
<< mvnsubdiff >>
rect 1357 9246 1480 9280
rect 1514 9246 1548 9280
rect 1357 9212 1548 9246
rect 1459 9178 1548 9212
rect 1459 9144 1616 9178
rect 1527 9110 1616 9144
rect 27966 9110 28085 9280
rect 27915 9036 28085 9110
rect 2191 8424 2273 8458
rect 2307 8424 2341 8458
rect 2191 8390 2341 8424
rect 2293 8356 2341 8390
rect 27195 8357 27263 8458
rect 27195 8356 27229 8357
rect 2293 8322 2409 8356
rect 2361 8288 2409 8322
rect 27127 8323 27229 8356
rect 27127 8289 27263 8323
rect 27127 8288 27161 8289
rect 2191 2790 2361 2916
rect 2293 2441 2361 2484
rect 27093 8221 27161 8288
rect 2293 2416 2327 2441
rect 2191 2382 2327 2416
rect 2225 2373 2327 2382
rect 27045 2407 27093 2441
rect 27045 2373 27161 2407
rect 2225 2348 2259 2373
rect 2191 2271 2259 2348
rect 27113 2339 27161 2373
rect 27113 2305 27263 2339
rect 27113 2271 27147 2305
rect 27181 2271 27263 2305
rect 1595 944 1630 978
rect 1664 944 1699 978
rect 1733 944 1768 978
rect 1802 944 1837 978
rect 1871 944 1906 978
rect 1940 944 1975 978
rect 2009 944 2044 978
rect 2078 944 2113 978
rect 2147 944 2182 978
rect 2216 944 2251 978
rect 2285 944 2320 978
rect 2354 944 2389 978
rect 2423 944 2458 978
rect 2492 944 2527 978
rect 2561 944 2596 978
rect 2630 944 2665 978
rect 2699 944 2734 978
rect 2768 944 2803 978
rect 2837 944 2872 978
rect 2906 944 2941 978
rect 2975 944 3010 978
rect 3044 944 3079 978
rect 3113 944 3148 978
rect 3182 944 3217 978
rect 3251 944 3286 978
rect 3320 944 3355 978
rect 3389 944 3424 978
rect 3458 944 3493 978
rect 3527 944 3562 978
rect 3596 944 3631 978
rect 3665 944 3700 978
rect 3734 944 3769 978
rect 3803 944 3838 978
rect 3872 944 3907 978
rect 3941 944 3976 978
rect 4010 944 4045 978
rect 4079 944 4114 978
rect 4148 944 4183 978
rect 1595 910 4183 944
rect 1357 876 1561 882
rect 1595 876 1630 910
rect 1664 876 1699 910
rect 1733 876 1768 910
rect 1802 876 1837 910
rect 1871 876 1906 910
rect 1940 876 1975 910
rect 2009 876 2044 910
rect 2078 876 2113 910
rect 2147 876 2182 910
rect 2216 876 2251 910
rect 2285 876 2320 910
rect 2354 876 2389 910
rect 2423 876 2458 910
rect 2492 876 2527 910
rect 2561 876 2596 910
rect 2630 876 2665 910
rect 2699 876 2734 910
rect 2768 876 2803 910
rect 2837 876 2872 910
rect 2906 876 2941 910
rect 2975 876 3010 910
rect 3044 876 3079 910
rect 3113 876 3148 910
rect 3182 876 3217 910
rect 3251 876 3286 910
rect 3320 876 3355 910
rect 3389 876 3424 910
rect 3458 876 3493 910
rect 3527 876 3562 910
rect 3596 876 3631 910
rect 3665 876 3700 910
rect 3734 876 3769 910
rect 3803 876 3838 910
rect 3872 876 3907 910
rect 3941 876 3976 910
rect 4010 876 4045 910
rect 4079 876 4114 910
rect 4148 876 4183 910
rect 1357 842 4183 876
rect 1357 808 1561 842
rect 1595 808 1630 842
rect 1664 808 1699 842
rect 1733 808 1768 842
rect 1802 808 1837 842
rect 1871 808 1906 842
rect 1940 808 1975 842
rect 2009 808 2044 842
rect 2078 808 2113 842
rect 2147 808 2182 842
rect 2216 808 2251 842
rect 2285 808 2320 842
rect 2354 808 2389 842
rect 2423 808 2458 842
rect 2492 808 2527 842
rect 2561 808 2596 842
rect 2630 808 2665 842
rect 2699 808 2734 842
rect 2768 808 2803 842
rect 2837 808 2872 842
rect 2906 808 2941 842
rect 2975 808 3010 842
rect 3044 808 3079 842
rect 3113 808 3148 842
rect 3182 808 3217 842
rect 3251 808 3286 842
rect 3320 808 3355 842
rect 3389 808 3424 842
rect 3458 808 3493 842
rect 3527 808 3562 842
rect 3596 808 3631 842
rect 3665 808 3700 842
rect 3734 808 3769 842
rect 3803 808 3838 842
rect 3872 808 3907 842
rect 3941 808 3976 842
rect 4010 808 4045 842
rect 4079 808 4114 842
rect 4148 808 4183 842
rect 27881 808 28085 842
<< mvpsubdiffcont >>
rect 1805 8741 1839 8775
rect 1873 8741 27407 8843
rect 27442 8809 27476 8843
rect 27511 8809 27545 8843
rect 27580 8809 27614 8843
rect 27442 8741 27476 8775
rect 27511 8741 27545 8775
rect 1805 8672 1839 8706
rect 1873 8672 1907 8706
rect 1941 8673 27339 8741
rect 27580 8707 27682 8775
rect 27374 8673 27408 8707
rect 27443 8673 27477 8707
rect 1805 8603 1839 8637
rect 1873 8603 1907 8637
rect 1941 8604 1975 8638
rect 1805 8534 1839 8568
rect 1873 8534 1907 8568
rect 1941 8535 1975 8569
rect 1805 8465 1839 8499
rect 1873 8465 1907 8499
rect 1941 8466 1975 8500
rect 1805 8396 1839 8430
rect 1873 8396 1907 8430
rect 1941 8397 1975 8431
rect 1805 8327 1839 8361
rect 1873 8327 1907 8361
rect 1941 8328 1975 8362
rect 1805 8258 1839 8292
rect 1873 8258 1907 8292
rect 1941 8259 1975 8293
rect 1805 8189 1839 8223
rect 1873 8189 1907 8223
rect 1941 8190 1975 8224
rect 1805 8120 1839 8154
rect 1873 8120 1907 8154
rect 1941 8121 1975 8155
rect 1805 8051 1839 8085
rect 1873 8051 1907 8085
rect 1941 8052 1975 8086
rect 1805 7982 1839 8016
rect 1873 7982 1907 8016
rect 1941 7983 1975 8017
rect 1805 7913 1839 7947
rect 1873 7913 1907 7947
rect 1941 7914 1975 7948
rect 1805 7844 1839 7878
rect 1873 7844 1907 7878
rect 1941 7845 1975 7879
rect 1805 7775 1839 7809
rect 1873 7775 1907 7809
rect 1941 7776 1975 7810
rect 1805 7706 1839 7740
rect 1873 7706 1907 7740
rect 1941 7707 1975 7741
rect 1805 7637 1839 7671
rect 1873 7637 1907 7671
rect 1941 7638 1975 7672
rect 1805 7568 1839 7602
rect 1873 7568 1907 7602
rect 1941 7569 1975 7603
rect 1805 7499 1839 7533
rect 1873 7499 1907 7533
rect 1941 7500 1975 7534
rect 1805 7430 1839 7464
rect 1873 7430 1907 7464
rect 1941 7431 1975 7465
rect 1805 7361 1839 7395
rect 1873 7361 1907 7395
rect 1941 7362 1975 7396
rect 1805 7292 1839 7326
rect 1873 7292 1907 7326
rect 1941 7293 1975 7327
rect 1805 7223 1839 7257
rect 1873 7223 1907 7257
rect 1941 7224 1975 7258
rect 1805 7154 1839 7188
rect 1873 7154 1907 7188
rect 1941 7155 1975 7189
rect 1805 7085 1839 7119
rect 1873 7085 1907 7119
rect 1941 7086 1975 7120
rect 1805 7016 1839 7050
rect 1873 7016 1907 7050
rect 1941 7017 1975 7051
rect 1805 6947 1839 6981
rect 1873 6947 1907 6981
rect 1941 6948 1975 6982
rect 1805 6878 1839 6912
rect 1873 6878 1907 6912
rect 1941 6879 1975 6913
rect 1805 6809 1839 6843
rect 1873 6809 1907 6843
rect 1941 6810 1975 6844
rect 1805 6740 1839 6774
rect 1873 6740 1907 6774
rect 1941 6741 1975 6775
rect 1805 6671 1839 6705
rect 1873 6671 1907 6705
rect 1941 6672 1975 6706
rect 1805 6602 1839 6636
rect 1873 6602 1907 6636
rect 1941 6603 1975 6637
rect 1805 6533 1839 6567
rect 1873 6533 1907 6567
rect 1941 6534 1975 6568
rect 1805 6464 1839 6498
rect 1873 6464 1907 6498
rect 1941 6465 1975 6499
rect 1805 6395 1839 6429
rect 1873 6395 1907 6429
rect 1941 6396 1975 6430
rect 1805 6326 1839 6360
rect 1873 6326 1907 6360
rect 1941 6327 1975 6361
rect 1805 6257 1839 6291
rect 1873 6257 1907 6291
rect 1941 6258 1975 6292
rect 1805 6188 1839 6222
rect 1873 6188 1907 6222
rect 1941 6189 1975 6223
rect 1805 6119 1839 6153
rect 1873 6119 1907 6153
rect 1941 6120 1975 6154
rect 1805 6050 1839 6084
rect 1873 6050 1907 6084
rect 1941 6051 1975 6085
rect 1805 5947 1907 6015
rect 1941 5982 1975 6016
rect 1805 5437 1975 5947
rect 1805 5335 1839 5369
rect 1873 5335 1907 5369
rect 1941 5335 1975 5369
rect 1805 5266 1839 5300
rect 1873 5266 1907 5300
rect 1941 5266 1975 5300
rect 1805 5197 1839 5231
rect 1873 5197 1907 5231
rect 1941 5197 1975 5231
rect 1805 5128 1839 5162
rect 1873 5128 1907 5162
rect 1941 5128 1975 5162
rect 1805 5059 1839 5093
rect 1873 5059 1907 5093
rect 1941 5059 1975 5093
rect 1805 4990 1839 5024
rect 1873 4990 1907 5024
rect 1941 4990 1975 5024
rect 1805 4921 1839 4955
rect 1873 4921 1907 4955
rect 1941 4921 1975 4955
rect 1805 4852 1839 4886
rect 1873 4852 1907 4886
rect 1941 4852 1975 4886
rect 1805 4783 1839 4817
rect 1873 4783 1907 4817
rect 1941 4783 1975 4817
rect 1805 4714 1839 4748
rect 1873 4714 1907 4748
rect 1941 4714 1975 4748
rect 1805 4645 1839 4679
rect 1873 4645 1907 4679
rect 1941 4645 1975 4679
rect 1805 4576 1839 4610
rect 1873 4576 1907 4610
rect 1941 4576 1975 4610
rect 1805 4507 1839 4541
rect 1873 4507 1907 4541
rect 1941 4507 1975 4541
rect 1805 4438 1839 4472
rect 1873 4438 1907 4472
rect 1941 4438 1975 4472
rect 1805 4369 1839 4403
rect 1873 4369 1907 4403
rect 1941 4369 1975 4403
rect 1805 4300 1839 4334
rect 1873 4300 1907 4334
rect 1941 4300 1975 4334
rect 1805 4231 1839 4265
rect 1873 4231 1907 4265
rect 1941 4231 1975 4265
rect 1805 4162 1839 4196
rect 1873 4162 1907 4196
rect 1941 4162 1975 4196
rect 1805 4093 1839 4127
rect 1873 4093 1907 4127
rect 1941 4093 1975 4127
rect 1805 4024 1839 4058
rect 1873 4024 1907 4058
rect 1941 4024 1975 4058
rect 1805 3955 1839 3989
rect 1873 3955 1907 3989
rect 1941 3955 1975 3989
rect 1805 1438 1975 3920
rect 27512 3301 27682 8707
rect 27512 3232 27546 3266
rect 27580 3233 27682 3301
rect 27512 3163 27546 3197
rect 27580 3164 27614 3198
rect 27648 3164 27682 3198
rect 27512 3094 27546 3128
rect 27580 3095 27614 3129
rect 27648 3095 27682 3129
rect 27512 3025 27546 3059
rect 27580 3026 27614 3060
rect 27648 3026 27682 3060
rect 27512 2956 27546 2990
rect 27580 2957 27614 2991
rect 27648 2957 27682 2991
rect 27512 2887 27546 2921
rect 27580 2888 27614 2922
rect 27648 2888 27682 2922
rect 27512 2818 27546 2852
rect 27580 2819 27614 2853
rect 27648 2819 27682 2853
rect 27512 2749 27546 2783
rect 27580 2750 27614 2784
rect 27648 2750 27682 2784
rect 27512 2680 27546 2714
rect 27580 2681 27614 2715
rect 27648 2681 27682 2715
rect 27512 2611 27546 2645
rect 27580 2612 27614 2646
rect 27648 2612 27682 2646
rect 27512 2542 27546 2576
rect 27580 2543 27614 2577
rect 27648 2543 27682 2577
rect 27512 2473 27546 2507
rect 27580 2474 27614 2508
rect 27648 2474 27682 2508
rect 27512 2404 27546 2438
rect 27580 2405 27614 2439
rect 27648 2405 27682 2439
rect 27512 2335 27546 2369
rect 27580 2336 27614 2370
rect 27648 2336 27682 2370
rect 27512 2266 27546 2300
rect 27580 2267 27614 2301
rect 27648 2267 27682 2301
rect 27512 2197 27546 2231
rect 27580 2198 27614 2232
rect 27648 2198 27682 2232
rect 27512 2128 27546 2162
rect 27580 2129 27614 2163
rect 27648 2129 27682 2163
rect 27512 2059 27546 2093
rect 27580 2060 27614 2094
rect 27648 2060 27682 2094
rect 2009 1961 2043 1995
rect 2078 1961 2112 1995
rect 2147 1961 2181 1995
rect 2216 1961 2250 1995
rect 2284 1961 2318 1995
rect 2352 1961 2386 1995
rect 2420 1961 2454 1995
rect 2488 1961 2522 1995
rect 2556 1961 2590 1995
rect 2624 1961 2658 1995
rect 2692 1961 2726 1995
rect 2760 1961 2794 1995
rect 2828 1961 2862 1995
rect 2896 1961 2930 1995
rect 2964 1961 2998 1995
rect 3032 1961 3066 1995
rect 3100 1961 3134 1995
rect 3168 1961 3202 1995
rect 3236 1961 3270 1995
rect 3304 1961 3338 1995
rect 3372 1961 3406 1995
rect 3440 1961 3474 1995
rect 3508 1961 3542 1995
rect 3576 1961 3610 1995
rect 3644 1961 3678 1995
rect 3712 1961 3746 1995
rect 3780 1961 3814 1995
rect 3848 1961 3882 1995
rect 3916 1961 3950 1995
rect 3984 1961 4018 1995
rect 4052 1961 4086 1995
rect 4120 1961 4154 1995
rect 4188 1961 4222 1995
rect 4256 1961 4290 1995
rect 4324 1961 4358 1995
rect 4392 1961 4426 1995
rect 4460 1961 4494 1995
rect 4528 1961 4562 1995
rect 4596 1961 4630 1995
rect 4664 1961 4698 1995
rect 4732 1961 4766 1995
rect 4800 1961 4834 1995
rect 4868 1961 4902 1995
rect 4936 1961 4970 1995
rect 5004 1961 5038 1995
rect 5072 1961 5106 1995
rect 5140 1961 5174 1995
rect 5208 1961 5242 1995
rect 5276 1961 5310 1995
rect 5344 1961 5378 1995
rect 5412 1961 5446 1995
rect 5480 1961 5514 1995
rect 5548 1961 5582 1995
rect 5616 1961 5650 1995
rect 5684 1961 5718 1995
rect 5752 1961 5786 1995
rect 5820 1961 5854 1995
rect 5888 1961 5922 1995
rect 5956 1961 5990 1995
rect 6024 1961 6058 1995
rect 6092 1961 6126 1995
rect 6160 1961 6194 1995
rect 6228 1961 6262 1995
rect 6296 1961 6330 1995
rect 6364 1961 6398 1995
rect 6432 1961 6466 1995
rect 6500 1961 6534 1995
rect 6568 1961 6602 1995
rect 6636 1961 6670 1995
rect 6704 1961 6738 1995
rect 6772 1961 6806 1995
rect 6840 1961 6874 1995
rect 6908 1961 6942 1995
rect 6976 1961 7010 1995
rect 7044 1961 7078 1995
rect 7112 1961 7146 1995
rect 7180 1961 7214 1995
rect 7248 1961 7282 1995
rect 7316 1961 7350 1995
rect 7384 1961 7418 1995
rect 7452 1961 7486 1995
rect 7520 1961 7554 1995
rect 7588 1961 7622 1995
rect 7656 1961 7690 1995
rect 7724 1961 7758 1995
rect 7792 1961 7826 1995
rect 7860 1961 7894 1995
rect 7928 1961 7962 1995
rect 7996 1961 8030 1995
rect 8064 1961 8098 1995
rect 8132 1961 8166 1995
rect 8200 1961 8234 1995
rect 8268 1961 8302 1995
rect 8336 1961 8370 1995
rect 8404 1961 8438 1995
rect 8472 1961 8506 1995
rect 8540 1961 8574 1995
rect 8608 1961 8642 1995
rect 8676 1961 8710 1995
rect 8744 1961 8778 1995
rect 8812 1961 8846 1995
rect 8880 1961 8914 1995
rect 8948 1961 8982 1995
rect 9016 1961 9050 1995
rect 9084 1961 9118 1995
rect 9152 1961 9186 1995
rect 9220 1961 9254 1995
rect 9288 1961 9322 1995
rect 9356 1961 9390 1995
rect 9424 1961 9458 1995
rect 9492 1961 9526 1995
rect 9560 1961 9594 1995
rect 9628 1961 9662 1995
rect 9696 1961 9730 1995
rect 9764 1961 9798 1995
rect 9832 1961 9866 1995
rect 9900 1961 9934 1995
rect 9968 1961 10002 1995
rect 10036 1961 10070 1995
rect 10104 1961 10138 1995
rect 10172 1961 10206 1995
rect 10240 1961 10274 1995
rect 10308 1961 10342 1995
rect 10376 1961 10410 1995
rect 10444 1961 10478 1995
rect 10512 1961 10546 1995
rect 10580 1961 10614 1995
rect 10648 1961 10682 1995
rect 10716 1961 10750 1995
rect 10784 1961 10818 1995
rect 10852 1961 10886 1995
rect 10920 1961 10954 1995
rect 10988 1961 11022 1995
rect 11056 1961 11090 1995
rect 11124 1961 11158 1995
rect 11192 1961 11226 1995
rect 11260 1961 11294 1995
rect 11328 1961 11362 1995
rect 11396 1961 11430 1995
rect 11464 1961 11498 1995
rect 11532 1961 11566 1995
rect 11600 1961 11634 1995
rect 11668 1961 11702 1995
rect 11736 1961 11770 1995
rect 11804 1961 11838 1995
rect 11872 1961 11906 1995
rect 11940 1961 11974 1995
rect 12008 1961 12042 1995
rect 12076 1961 12110 1995
rect 12144 1961 12178 1995
rect 12212 1961 12246 1995
rect 12280 1961 12314 1995
rect 12348 1961 12382 1995
rect 12416 1961 12450 1995
rect 12484 1961 12518 1995
rect 12552 1961 12586 1995
rect 12620 1961 12654 1995
rect 12688 1961 12722 1995
rect 12756 1961 12790 1995
rect 12824 1961 12858 1995
rect 12892 1961 12926 1995
rect 12960 1961 12994 1995
rect 13028 1961 13062 1995
rect 13096 1961 13130 1995
rect 13164 1961 13198 1995
rect 13232 1961 13266 1995
rect 13300 1961 13334 1995
rect 13368 1961 13402 1995
rect 13436 1961 13470 1995
rect 13504 1961 13538 1995
rect 13572 1961 13606 1995
rect 13640 1961 13674 1995
rect 13708 1961 13742 1995
rect 13776 1961 13810 1995
rect 13844 1961 13878 1995
rect 13912 1961 13946 1995
rect 13980 1961 14014 1995
rect 14048 1961 14082 1995
rect 14116 1961 14150 1995
rect 14184 1961 14218 1995
rect 14252 1961 14286 1995
rect 14320 1961 14354 1995
rect 14388 1961 14422 1995
rect 14456 1961 14490 1995
rect 14524 1961 14558 1995
rect 14592 1961 14626 1995
rect 14660 1961 14694 1995
rect 14728 1961 14762 1995
rect 14796 1961 14830 1995
rect 14864 1961 14898 1995
rect 14932 1961 14966 1995
rect 15000 1961 15034 1995
rect 15068 1961 15102 1995
rect 15136 1961 15170 1995
rect 15204 1961 15238 1995
rect 15272 1961 15306 1995
rect 15340 1961 15374 1995
rect 15408 1961 15442 1995
rect 15476 1961 15510 1995
rect 15544 1961 15578 1995
rect 15612 1961 15646 1995
rect 15680 1961 15714 1995
rect 15748 1961 15782 1995
rect 15816 1961 15850 1995
rect 15884 1961 15918 1995
rect 15952 1961 15986 1995
rect 16020 1961 16054 1995
rect 16088 1961 16122 1995
rect 16156 1961 16190 1995
rect 16224 1961 16258 1995
rect 16292 1961 16326 1995
rect 16360 1961 16394 1995
rect 16428 1961 16462 1995
rect 16496 1961 16530 1995
rect 16564 1961 16598 1995
rect 16632 1961 16666 1995
rect 16700 1961 16734 1995
rect 16768 1961 16802 1995
rect 16836 1961 16870 1995
rect 16904 1961 16938 1995
rect 16972 1961 17006 1995
rect 17040 1961 17074 1995
rect 17108 1961 17142 1995
rect 17176 1961 17210 1995
rect 17244 1961 17278 1995
rect 17312 1961 17346 1995
rect 17380 1961 17414 1995
rect 17448 1961 17482 1995
rect 17516 1961 17550 1995
rect 17584 1961 17618 1995
rect 17652 1961 17686 1995
rect 17720 1961 17754 1995
rect 17788 1961 17822 1995
rect 17856 1961 17890 1995
rect 17924 1961 17958 1995
rect 17992 1961 18026 1995
rect 18060 1961 18094 1995
rect 18128 1961 18162 1995
rect 18196 1961 18230 1995
rect 18264 1961 18298 1995
rect 18332 1961 18366 1995
rect 18400 1961 18434 1995
rect 18468 1961 18502 1995
rect 18536 1961 18570 1995
rect 18604 1961 18638 1995
rect 18672 1961 18706 1995
rect 18740 1961 18774 1995
rect 18808 1961 18842 1995
rect 18876 1961 18910 1995
rect 18944 1961 18978 1995
rect 19012 1961 19046 1995
rect 19080 1961 19114 1995
rect 19148 1961 19182 1995
rect 19216 1961 19250 1995
rect 19284 1961 19318 1995
rect 19352 1961 19386 1995
rect 19420 1961 19454 1995
rect 19488 1961 19522 1995
rect 19556 1961 19590 1995
rect 19624 1961 19658 1995
rect 19692 1961 19726 1995
rect 19760 1961 19794 1995
rect 19828 1961 19862 1995
rect 19896 1961 19930 1995
rect 19964 1961 19998 1995
rect 20032 1961 20066 1995
rect 20100 1961 20134 1995
rect 20168 1961 20202 1995
rect 20236 1961 20270 1995
rect 20304 1961 20338 1995
rect 20372 1961 20406 1995
rect 20440 1961 20474 1995
rect 20508 1961 20542 1995
rect 20576 1961 20610 1995
rect 20644 1961 20678 1995
rect 20712 1961 20746 1995
rect 20780 1961 20814 1995
rect 20848 1961 20882 1995
rect 20916 1961 20950 1995
rect 20984 1961 21018 1995
rect 21052 1961 21086 1995
rect 21120 1961 21154 1995
rect 21188 1961 21222 1995
rect 21256 1961 21290 1995
rect 21324 1961 21358 1995
rect 21392 1961 21426 1995
rect 21460 1961 21494 1995
rect 21528 1961 21562 1995
rect 21596 1961 21630 1995
rect 21664 1961 21698 1995
rect 21732 1961 21766 1995
rect 21800 1961 21834 1995
rect 21868 1961 21902 1995
rect 21936 1961 21970 1995
rect 22004 1961 22038 1995
rect 22072 1961 22106 1995
rect 22140 1961 22174 1995
rect 22208 1961 22242 1995
rect 22276 1961 22310 1995
rect 22344 1961 22378 1995
rect 22412 1961 22446 1995
rect 22480 1961 22514 1995
rect 22548 1961 22582 1995
rect 22616 1961 22650 1995
rect 22684 1961 22718 1995
rect 22752 1961 22786 1995
rect 22820 1961 22854 1995
rect 22888 1961 22922 1995
rect 22956 1961 22990 1995
rect 23024 1961 23058 1995
rect 23092 1961 23126 1995
rect 23160 1961 23194 1995
rect 23228 1961 23262 1995
rect 23296 1961 23330 1995
rect 23364 1961 23398 1995
rect 23432 1961 23466 1995
rect 23500 1961 23534 1995
rect 23568 1961 23602 1995
rect 23636 1961 23670 1995
rect 23704 1961 23738 1995
rect 23772 1961 23806 1995
rect 23840 1961 23874 1995
rect 23908 1961 23942 1995
rect 23976 1961 24010 1995
rect 24044 1961 24078 1995
rect 24112 1961 24146 1995
rect 24180 1961 24214 1995
rect 24248 1961 24282 1995
rect 24316 1961 24350 1995
rect 24384 1961 24418 1995
rect 24452 1961 24486 1995
rect 24520 1961 24554 1995
rect 24588 1961 24622 1995
rect 24656 1961 24690 1995
rect 24724 1961 24758 1995
rect 24792 1961 24826 1995
rect 24860 1961 24894 1995
rect 24928 1961 24962 1995
rect 24996 1961 25030 1995
rect 25064 1961 25098 1995
rect 25132 1961 25166 1995
rect 25200 1961 25234 1995
rect 25268 1961 25302 1995
rect 25336 1961 25370 1995
rect 25404 1961 25438 1995
rect 25472 1961 25506 1995
rect 25540 1961 25574 1995
rect 25608 1961 25642 1995
rect 25676 1961 25710 1995
rect 25744 1961 25778 1995
rect 25812 1961 25846 1995
rect 25880 1961 25914 1995
rect 25948 1961 25982 1995
rect 26016 1961 26050 1995
rect 26084 1961 26118 1995
rect 26152 1961 26186 1995
rect 26220 1961 26254 1995
rect 26288 1961 26322 1995
rect 26356 1961 26390 1995
rect 26424 1961 26458 1995
rect 26492 1961 26526 1995
rect 26560 1961 26594 1995
rect 26628 1961 26662 1995
rect 26696 1961 26730 1995
rect 26764 1961 26798 1995
rect 26832 1961 26866 1995
rect 26900 1961 26934 1995
rect 26968 1961 27002 1995
rect 27036 1961 27070 1995
rect 27104 1961 27138 1995
rect 27172 1961 27206 1995
rect 27240 1961 27274 1995
rect 27308 1961 27342 1995
rect 27376 1961 27410 1995
rect 27444 1961 27478 1995
rect 27512 1990 27546 2024
rect 27580 1991 27614 2025
rect 27648 1991 27682 2025
rect 27512 1921 27546 1955
rect 27580 1922 27614 1956
rect 27648 1922 27682 1956
rect 2009 1887 2043 1921
rect 2078 1887 2112 1921
rect 2147 1887 2181 1921
rect 2216 1887 2250 1921
rect 2284 1887 2318 1921
rect 2352 1887 2386 1921
rect 2420 1887 2454 1921
rect 2488 1887 2522 1921
rect 2556 1887 2590 1921
rect 2624 1887 2658 1921
rect 2692 1887 2726 1921
rect 2760 1887 2794 1921
rect 2828 1887 2862 1921
rect 2896 1887 2930 1921
rect 2964 1887 2998 1921
rect 3032 1887 3066 1921
rect 3100 1887 3134 1921
rect 3168 1887 3202 1921
rect 3236 1887 3270 1921
rect 3304 1887 3338 1921
rect 3372 1887 3406 1921
rect 3440 1887 3474 1921
rect 3508 1887 3542 1921
rect 3576 1887 3610 1921
rect 3644 1887 3678 1921
rect 3712 1887 3746 1921
rect 3780 1887 3814 1921
rect 3848 1887 3882 1921
rect 3916 1887 3950 1921
rect 3984 1887 4018 1921
rect 4052 1887 4086 1921
rect 4120 1887 4154 1921
rect 4188 1887 4222 1921
rect 4256 1887 4290 1921
rect 4324 1887 4358 1921
rect 4392 1887 4426 1921
rect 4460 1887 4494 1921
rect 4528 1887 4562 1921
rect 4596 1887 4630 1921
rect 4664 1887 4698 1921
rect 4732 1887 4766 1921
rect 4800 1887 4834 1921
rect 4868 1887 4902 1921
rect 4936 1887 4970 1921
rect 5004 1887 5038 1921
rect 5072 1887 5106 1921
rect 5140 1887 5174 1921
rect 5208 1887 5242 1921
rect 5276 1887 5310 1921
rect 5344 1887 5378 1921
rect 5412 1887 5446 1921
rect 5480 1887 5514 1921
rect 5548 1887 5582 1921
rect 5616 1887 5650 1921
rect 5684 1887 5718 1921
rect 5752 1887 5786 1921
rect 5820 1887 5854 1921
rect 5888 1887 5922 1921
rect 5956 1887 5990 1921
rect 6024 1887 6058 1921
rect 6092 1887 6126 1921
rect 6160 1887 6194 1921
rect 6228 1887 6262 1921
rect 6296 1887 6330 1921
rect 6364 1887 6398 1921
rect 6432 1887 6466 1921
rect 6500 1887 6534 1921
rect 6568 1887 6602 1921
rect 6636 1887 6670 1921
rect 6704 1887 6738 1921
rect 6772 1887 6806 1921
rect 6840 1887 6874 1921
rect 6908 1887 6942 1921
rect 6976 1887 7010 1921
rect 7044 1887 7078 1921
rect 7112 1887 7146 1921
rect 7180 1887 7214 1921
rect 7248 1887 7282 1921
rect 7316 1887 7350 1921
rect 7384 1887 7418 1921
rect 7452 1887 7486 1921
rect 7520 1887 7554 1921
rect 7588 1887 7622 1921
rect 7656 1887 7690 1921
rect 7724 1887 7758 1921
rect 7792 1887 7826 1921
rect 7860 1887 7894 1921
rect 7928 1887 7962 1921
rect 7996 1887 8030 1921
rect 8064 1887 8098 1921
rect 8132 1887 8166 1921
rect 8200 1887 8234 1921
rect 8268 1887 8302 1921
rect 8336 1887 8370 1921
rect 8404 1887 8438 1921
rect 8472 1887 8506 1921
rect 8540 1887 8574 1921
rect 8608 1887 8642 1921
rect 8676 1887 8710 1921
rect 8744 1887 8778 1921
rect 8812 1887 8846 1921
rect 8880 1887 8914 1921
rect 8948 1887 8982 1921
rect 9016 1887 9050 1921
rect 9084 1887 9118 1921
rect 9152 1887 9186 1921
rect 9220 1887 9254 1921
rect 9288 1887 9322 1921
rect 9356 1887 9390 1921
rect 9424 1887 9458 1921
rect 9492 1887 9526 1921
rect 9560 1887 9594 1921
rect 9628 1887 9662 1921
rect 9696 1887 9730 1921
rect 9764 1887 9798 1921
rect 9832 1887 9866 1921
rect 9900 1887 9934 1921
rect 9968 1887 10002 1921
rect 10036 1887 10070 1921
rect 10104 1887 10138 1921
rect 10172 1887 10206 1921
rect 10240 1887 10274 1921
rect 10308 1887 10342 1921
rect 10376 1887 10410 1921
rect 10444 1887 10478 1921
rect 10512 1887 10546 1921
rect 10580 1887 10614 1921
rect 10648 1887 10682 1921
rect 10716 1887 10750 1921
rect 10784 1887 10818 1921
rect 10852 1887 10886 1921
rect 10920 1887 10954 1921
rect 10988 1887 11022 1921
rect 11056 1887 11090 1921
rect 11124 1887 11158 1921
rect 11192 1887 11226 1921
rect 11260 1887 11294 1921
rect 11328 1887 11362 1921
rect 11396 1887 11430 1921
rect 11464 1887 11498 1921
rect 11532 1887 11566 1921
rect 11600 1887 11634 1921
rect 11668 1887 11702 1921
rect 11736 1887 11770 1921
rect 11804 1887 11838 1921
rect 11872 1887 11906 1921
rect 11940 1887 11974 1921
rect 12008 1887 12042 1921
rect 12076 1887 12110 1921
rect 12144 1887 12178 1921
rect 12212 1887 12246 1921
rect 12280 1887 12314 1921
rect 12348 1887 12382 1921
rect 12416 1887 12450 1921
rect 12484 1887 12518 1921
rect 12552 1887 12586 1921
rect 12620 1887 12654 1921
rect 12688 1887 12722 1921
rect 12756 1887 12790 1921
rect 12824 1887 12858 1921
rect 12892 1887 12926 1921
rect 12960 1887 12994 1921
rect 13028 1887 13062 1921
rect 13096 1887 13130 1921
rect 13164 1887 13198 1921
rect 13232 1887 13266 1921
rect 13300 1887 13334 1921
rect 13368 1887 13402 1921
rect 13436 1887 13470 1921
rect 13504 1887 13538 1921
rect 13572 1887 13606 1921
rect 13640 1887 13674 1921
rect 13708 1887 13742 1921
rect 13776 1887 13810 1921
rect 13844 1887 13878 1921
rect 13912 1887 13946 1921
rect 13980 1887 14014 1921
rect 14048 1887 14082 1921
rect 14116 1887 14150 1921
rect 14184 1887 14218 1921
rect 14252 1887 14286 1921
rect 14320 1887 14354 1921
rect 14388 1887 14422 1921
rect 14456 1887 14490 1921
rect 14524 1887 14558 1921
rect 14592 1887 14626 1921
rect 14660 1887 14694 1921
rect 14728 1887 14762 1921
rect 14796 1887 14830 1921
rect 14864 1887 14898 1921
rect 14932 1887 14966 1921
rect 15000 1887 15034 1921
rect 15068 1887 15102 1921
rect 15136 1887 15170 1921
rect 15204 1887 15238 1921
rect 15272 1887 15306 1921
rect 15340 1887 15374 1921
rect 15408 1887 15442 1921
rect 15476 1887 15510 1921
rect 15544 1887 15578 1921
rect 15612 1887 15646 1921
rect 15680 1887 15714 1921
rect 15748 1887 15782 1921
rect 15816 1887 15850 1921
rect 15884 1887 15918 1921
rect 15952 1887 15986 1921
rect 16020 1887 16054 1921
rect 16088 1887 16122 1921
rect 16156 1887 16190 1921
rect 16224 1887 16258 1921
rect 16292 1887 16326 1921
rect 16360 1887 16394 1921
rect 16428 1887 16462 1921
rect 16496 1887 16530 1921
rect 16564 1887 16598 1921
rect 16632 1887 16666 1921
rect 16700 1887 16734 1921
rect 16768 1887 16802 1921
rect 16836 1887 16870 1921
rect 16904 1887 16938 1921
rect 16972 1887 17006 1921
rect 17040 1887 17074 1921
rect 17108 1887 17142 1921
rect 17176 1887 17210 1921
rect 17244 1887 17278 1921
rect 17312 1887 17346 1921
rect 17380 1887 17414 1921
rect 17448 1887 17482 1921
rect 17516 1887 17550 1921
rect 17584 1887 17618 1921
rect 17652 1887 17686 1921
rect 17720 1887 17754 1921
rect 17788 1887 17822 1921
rect 17856 1887 17890 1921
rect 17924 1887 17958 1921
rect 17992 1887 18026 1921
rect 18060 1887 18094 1921
rect 18128 1887 18162 1921
rect 18196 1887 18230 1921
rect 18264 1887 18298 1921
rect 18332 1887 18366 1921
rect 18400 1887 18434 1921
rect 18468 1887 18502 1921
rect 18536 1887 18570 1921
rect 18604 1887 18638 1921
rect 18672 1887 18706 1921
rect 18740 1887 18774 1921
rect 18808 1887 18842 1921
rect 18876 1887 18910 1921
rect 18944 1887 18978 1921
rect 19012 1887 19046 1921
rect 19080 1887 19114 1921
rect 19148 1887 19182 1921
rect 19216 1887 19250 1921
rect 19284 1887 19318 1921
rect 19352 1887 19386 1921
rect 19420 1887 19454 1921
rect 19488 1887 19522 1921
rect 19556 1887 19590 1921
rect 19624 1887 19658 1921
rect 19692 1887 19726 1921
rect 19760 1887 19794 1921
rect 19828 1887 19862 1921
rect 19896 1887 19930 1921
rect 19964 1887 19998 1921
rect 20032 1887 20066 1921
rect 20100 1887 20134 1921
rect 20168 1887 20202 1921
rect 20236 1887 20270 1921
rect 20304 1887 20338 1921
rect 20372 1887 20406 1921
rect 20440 1887 20474 1921
rect 20508 1887 20542 1921
rect 20576 1887 20610 1921
rect 20644 1887 20678 1921
rect 20712 1887 20746 1921
rect 20780 1887 20814 1921
rect 20848 1887 20882 1921
rect 20916 1887 20950 1921
rect 20984 1887 21018 1921
rect 21052 1887 21086 1921
rect 21120 1887 21154 1921
rect 21188 1887 21222 1921
rect 21256 1887 21290 1921
rect 21324 1887 21358 1921
rect 21392 1887 21426 1921
rect 21460 1887 21494 1921
rect 21528 1887 21562 1921
rect 21596 1887 21630 1921
rect 21664 1887 21698 1921
rect 21732 1887 21766 1921
rect 21800 1887 21834 1921
rect 21868 1887 21902 1921
rect 21936 1887 21970 1921
rect 22004 1887 22038 1921
rect 22072 1887 22106 1921
rect 22140 1887 22174 1921
rect 22208 1887 22242 1921
rect 22276 1887 22310 1921
rect 22344 1887 22378 1921
rect 22412 1887 22446 1921
rect 22480 1887 22514 1921
rect 22548 1887 22582 1921
rect 22616 1887 22650 1921
rect 22684 1887 22718 1921
rect 22752 1887 22786 1921
rect 22820 1887 22854 1921
rect 22888 1887 22922 1921
rect 22956 1887 22990 1921
rect 23024 1887 23058 1921
rect 23092 1887 23126 1921
rect 23160 1887 23194 1921
rect 23228 1887 23262 1921
rect 23296 1887 23330 1921
rect 23364 1887 23398 1921
rect 23432 1887 23466 1921
rect 23500 1887 23534 1921
rect 23568 1887 23602 1921
rect 23636 1887 23670 1921
rect 23704 1887 23738 1921
rect 23772 1887 23806 1921
rect 23840 1887 23874 1921
rect 23908 1887 23942 1921
rect 23976 1887 24010 1921
rect 24044 1887 24078 1921
rect 24112 1887 24146 1921
rect 24180 1887 24214 1921
rect 24248 1887 24282 1921
rect 24316 1887 24350 1921
rect 24384 1887 24418 1921
rect 24452 1887 24486 1921
rect 24520 1887 24554 1921
rect 24588 1887 24622 1921
rect 24656 1887 24690 1921
rect 24724 1887 24758 1921
rect 24792 1887 24826 1921
rect 24860 1887 24894 1921
rect 24928 1887 24962 1921
rect 24996 1887 25030 1921
rect 25064 1887 25098 1921
rect 25132 1887 25166 1921
rect 25200 1887 25234 1921
rect 25268 1887 25302 1921
rect 25336 1887 25370 1921
rect 25404 1887 25438 1921
rect 25472 1887 25506 1921
rect 25540 1887 25574 1921
rect 25608 1887 25642 1921
rect 25676 1887 25710 1921
rect 25744 1887 25778 1921
rect 25812 1887 25846 1921
rect 25880 1887 25914 1921
rect 25948 1887 25982 1921
rect 26016 1887 26050 1921
rect 26084 1887 26118 1921
rect 26152 1887 26186 1921
rect 26220 1887 26254 1921
rect 26288 1887 26322 1921
rect 26356 1887 26390 1921
rect 26424 1887 26458 1921
rect 26492 1887 26526 1921
rect 26560 1887 26594 1921
rect 26628 1887 26662 1921
rect 26696 1887 26730 1921
rect 26764 1887 26798 1921
rect 26832 1887 26866 1921
rect 26900 1887 26934 1921
rect 26968 1887 27002 1921
rect 27036 1887 27070 1921
rect 27104 1887 27138 1921
rect 27172 1887 27206 1921
rect 27240 1887 27274 1921
rect 27308 1887 27342 1921
rect 27376 1887 27410 1921
rect 27444 1887 27478 1921
rect 27512 1852 27546 1886
rect 27580 1853 27614 1887
rect 27648 1853 27682 1887
rect 2009 1813 2043 1847
rect 2078 1813 2112 1847
rect 2147 1813 2181 1847
rect 2216 1813 2250 1847
rect 2284 1813 2318 1847
rect 2352 1813 2386 1847
rect 2420 1813 2454 1847
rect 2488 1813 2522 1847
rect 2556 1813 2590 1847
rect 2624 1813 2658 1847
rect 2692 1813 2726 1847
rect 2760 1813 2794 1847
rect 2828 1813 2862 1847
rect 2896 1813 2930 1847
rect 2964 1813 2998 1847
rect 3032 1813 3066 1847
rect 3100 1813 3134 1847
rect 3168 1813 3202 1847
rect 3236 1813 3270 1847
rect 3304 1813 3338 1847
rect 3372 1813 3406 1847
rect 3440 1813 3474 1847
rect 3508 1813 3542 1847
rect 3576 1813 3610 1847
rect 3644 1813 3678 1847
rect 3712 1813 3746 1847
rect 3780 1813 3814 1847
rect 3848 1813 3882 1847
rect 3916 1813 3950 1847
rect 3984 1813 4018 1847
rect 4052 1813 4086 1847
rect 4120 1813 4154 1847
rect 4188 1813 4222 1847
rect 4256 1813 4290 1847
rect 4324 1813 4358 1847
rect 4392 1813 4426 1847
rect 4460 1813 4494 1847
rect 4528 1813 4562 1847
rect 4596 1813 4630 1847
rect 4664 1813 4698 1847
rect 4732 1813 4766 1847
rect 4800 1813 4834 1847
rect 4868 1813 4902 1847
rect 4936 1813 4970 1847
rect 5004 1813 5038 1847
rect 5072 1813 5106 1847
rect 5140 1813 5174 1847
rect 5208 1813 5242 1847
rect 5276 1813 5310 1847
rect 5344 1813 5378 1847
rect 5412 1813 5446 1847
rect 5480 1813 5514 1847
rect 5548 1813 5582 1847
rect 5616 1813 5650 1847
rect 5684 1813 5718 1847
rect 5752 1813 5786 1847
rect 5820 1813 5854 1847
rect 5888 1813 5922 1847
rect 5956 1813 5990 1847
rect 6024 1813 6058 1847
rect 6092 1813 6126 1847
rect 6160 1813 6194 1847
rect 6228 1813 6262 1847
rect 6296 1813 6330 1847
rect 6364 1813 6398 1847
rect 6432 1813 6466 1847
rect 6500 1813 6534 1847
rect 6568 1813 6602 1847
rect 6636 1813 6670 1847
rect 6704 1813 6738 1847
rect 6772 1813 6806 1847
rect 6840 1813 6874 1847
rect 6908 1813 6942 1847
rect 6976 1813 7010 1847
rect 7044 1813 7078 1847
rect 7112 1813 7146 1847
rect 7180 1813 7214 1847
rect 7248 1813 7282 1847
rect 7316 1813 7350 1847
rect 7384 1813 7418 1847
rect 7452 1813 7486 1847
rect 7520 1813 7554 1847
rect 7588 1813 7622 1847
rect 7656 1813 7690 1847
rect 7724 1813 7758 1847
rect 7792 1813 7826 1847
rect 7860 1813 7894 1847
rect 7928 1813 7962 1847
rect 7996 1813 8030 1847
rect 8064 1813 8098 1847
rect 8132 1813 8166 1847
rect 8200 1813 8234 1847
rect 8268 1813 8302 1847
rect 8336 1813 8370 1847
rect 8404 1813 8438 1847
rect 8472 1813 8506 1847
rect 8540 1813 8574 1847
rect 8608 1813 8642 1847
rect 8676 1813 8710 1847
rect 8744 1813 8778 1847
rect 8812 1813 8846 1847
rect 8880 1813 8914 1847
rect 8948 1813 8982 1847
rect 9016 1813 9050 1847
rect 9084 1813 9118 1847
rect 9152 1813 9186 1847
rect 9220 1813 9254 1847
rect 9288 1813 9322 1847
rect 9356 1813 9390 1847
rect 9424 1813 9458 1847
rect 9492 1813 9526 1847
rect 9560 1813 9594 1847
rect 9628 1813 9662 1847
rect 9696 1813 9730 1847
rect 9764 1813 9798 1847
rect 9832 1813 9866 1847
rect 9900 1813 9934 1847
rect 9968 1813 10002 1847
rect 10036 1813 10070 1847
rect 10104 1813 10138 1847
rect 10172 1813 10206 1847
rect 10240 1813 10274 1847
rect 10308 1813 10342 1847
rect 10376 1813 10410 1847
rect 10444 1813 10478 1847
rect 10512 1813 10546 1847
rect 10580 1813 10614 1847
rect 10648 1813 10682 1847
rect 10716 1813 10750 1847
rect 10784 1813 10818 1847
rect 10852 1813 10886 1847
rect 10920 1813 10954 1847
rect 10988 1813 11022 1847
rect 11056 1813 11090 1847
rect 11124 1813 11158 1847
rect 11192 1813 11226 1847
rect 11260 1813 11294 1847
rect 11328 1813 11362 1847
rect 11396 1813 11430 1847
rect 11464 1813 11498 1847
rect 11532 1813 11566 1847
rect 11600 1813 11634 1847
rect 11668 1813 11702 1847
rect 11736 1813 11770 1847
rect 11804 1813 11838 1847
rect 11872 1813 11906 1847
rect 11940 1813 11974 1847
rect 12008 1813 12042 1847
rect 12076 1813 12110 1847
rect 12144 1813 12178 1847
rect 12212 1813 12246 1847
rect 12280 1813 12314 1847
rect 12348 1813 12382 1847
rect 12416 1813 12450 1847
rect 12484 1813 12518 1847
rect 12552 1813 12586 1847
rect 12620 1813 12654 1847
rect 12688 1813 12722 1847
rect 12756 1813 12790 1847
rect 12824 1813 12858 1847
rect 12892 1813 12926 1847
rect 12960 1813 12994 1847
rect 13028 1813 13062 1847
rect 13096 1813 13130 1847
rect 13164 1813 13198 1847
rect 13232 1813 13266 1847
rect 13300 1813 13334 1847
rect 13368 1813 13402 1847
rect 13436 1813 13470 1847
rect 13504 1813 13538 1847
rect 13572 1813 13606 1847
rect 13640 1813 13674 1847
rect 13708 1813 13742 1847
rect 13776 1813 13810 1847
rect 13844 1813 13878 1847
rect 13912 1813 13946 1847
rect 13980 1813 14014 1847
rect 14048 1813 14082 1847
rect 14116 1813 14150 1847
rect 14184 1813 14218 1847
rect 14252 1813 14286 1847
rect 14320 1813 14354 1847
rect 14388 1813 14422 1847
rect 14456 1813 14490 1847
rect 14524 1813 14558 1847
rect 14592 1813 14626 1847
rect 14660 1813 14694 1847
rect 14728 1813 14762 1847
rect 14796 1813 14830 1847
rect 14864 1813 14898 1847
rect 14932 1813 14966 1847
rect 15000 1813 15034 1847
rect 15068 1813 15102 1847
rect 15136 1813 15170 1847
rect 15204 1813 15238 1847
rect 15272 1813 15306 1847
rect 15340 1813 15374 1847
rect 15408 1813 15442 1847
rect 15476 1813 15510 1847
rect 15544 1813 15578 1847
rect 15612 1813 15646 1847
rect 15680 1813 15714 1847
rect 15748 1813 15782 1847
rect 15816 1813 15850 1847
rect 15884 1813 15918 1847
rect 15952 1813 15986 1847
rect 16020 1813 16054 1847
rect 16088 1813 16122 1847
rect 16156 1813 16190 1847
rect 16224 1813 16258 1847
rect 16292 1813 16326 1847
rect 16360 1813 16394 1847
rect 16428 1813 16462 1847
rect 16496 1813 16530 1847
rect 16564 1813 16598 1847
rect 16632 1813 16666 1847
rect 16700 1813 16734 1847
rect 16768 1813 16802 1847
rect 16836 1813 16870 1847
rect 16904 1813 16938 1847
rect 16972 1813 17006 1847
rect 17040 1813 17074 1847
rect 17108 1813 17142 1847
rect 17176 1813 17210 1847
rect 17244 1813 17278 1847
rect 17312 1813 17346 1847
rect 17380 1813 17414 1847
rect 17448 1813 17482 1847
rect 17516 1813 17550 1847
rect 17584 1813 17618 1847
rect 17652 1813 17686 1847
rect 17720 1813 17754 1847
rect 17788 1813 17822 1847
rect 17856 1813 17890 1847
rect 17924 1813 17958 1847
rect 17992 1813 18026 1847
rect 18060 1813 18094 1847
rect 18128 1813 18162 1847
rect 18196 1813 18230 1847
rect 18264 1813 18298 1847
rect 18332 1813 18366 1847
rect 18400 1813 18434 1847
rect 18468 1813 18502 1847
rect 18536 1813 18570 1847
rect 18604 1813 18638 1847
rect 18672 1813 18706 1847
rect 18740 1813 18774 1847
rect 18808 1813 18842 1847
rect 18876 1813 18910 1847
rect 18944 1813 18978 1847
rect 19012 1813 19046 1847
rect 19080 1813 19114 1847
rect 19148 1813 19182 1847
rect 19216 1813 19250 1847
rect 19284 1813 19318 1847
rect 19352 1813 19386 1847
rect 19420 1813 19454 1847
rect 19488 1813 19522 1847
rect 19556 1813 19590 1847
rect 19624 1813 19658 1847
rect 19692 1813 19726 1847
rect 19760 1813 19794 1847
rect 19828 1813 19862 1847
rect 19896 1813 19930 1847
rect 19964 1813 19998 1847
rect 20032 1813 20066 1847
rect 20100 1813 20134 1847
rect 20168 1813 20202 1847
rect 20236 1813 20270 1847
rect 20304 1813 20338 1847
rect 20372 1813 20406 1847
rect 20440 1813 20474 1847
rect 20508 1813 20542 1847
rect 20576 1813 20610 1847
rect 20644 1813 20678 1847
rect 20712 1813 20746 1847
rect 20780 1813 20814 1847
rect 20848 1813 20882 1847
rect 20916 1813 20950 1847
rect 20984 1813 21018 1847
rect 21052 1813 21086 1847
rect 21120 1813 21154 1847
rect 21188 1813 21222 1847
rect 21256 1813 21290 1847
rect 21324 1813 21358 1847
rect 21392 1813 21426 1847
rect 21460 1813 21494 1847
rect 21528 1813 21562 1847
rect 21596 1813 21630 1847
rect 21664 1813 21698 1847
rect 21732 1813 21766 1847
rect 21800 1813 21834 1847
rect 21868 1813 21902 1847
rect 21936 1813 21970 1847
rect 22004 1813 22038 1847
rect 22072 1813 22106 1847
rect 22140 1813 22174 1847
rect 22208 1813 22242 1847
rect 22276 1813 22310 1847
rect 22344 1813 22378 1847
rect 22412 1813 22446 1847
rect 22480 1813 22514 1847
rect 22548 1813 22582 1847
rect 22616 1813 22650 1847
rect 22684 1813 22718 1847
rect 22752 1813 22786 1847
rect 22820 1813 22854 1847
rect 22888 1813 22922 1847
rect 22956 1813 22990 1847
rect 23024 1813 23058 1847
rect 23092 1813 23126 1847
rect 23160 1813 23194 1847
rect 23228 1813 23262 1847
rect 23296 1813 23330 1847
rect 23364 1813 23398 1847
rect 23432 1813 23466 1847
rect 23500 1813 23534 1847
rect 23568 1813 23602 1847
rect 23636 1813 23670 1847
rect 23704 1813 23738 1847
rect 23772 1813 23806 1847
rect 23840 1813 23874 1847
rect 23908 1813 23942 1847
rect 23976 1813 24010 1847
rect 24044 1813 24078 1847
rect 24112 1813 24146 1847
rect 24180 1813 24214 1847
rect 24248 1813 24282 1847
rect 24316 1813 24350 1847
rect 24384 1813 24418 1847
rect 24452 1813 24486 1847
rect 24520 1813 24554 1847
rect 24588 1813 24622 1847
rect 24656 1813 24690 1847
rect 24724 1813 24758 1847
rect 24792 1813 24826 1847
rect 24860 1813 24894 1847
rect 24928 1813 24962 1847
rect 24996 1813 25030 1847
rect 25064 1813 25098 1847
rect 25132 1813 25166 1847
rect 25200 1813 25234 1847
rect 25268 1813 25302 1847
rect 25336 1813 25370 1847
rect 25404 1813 25438 1847
rect 25472 1813 25506 1847
rect 25540 1813 25574 1847
rect 25608 1813 25642 1847
rect 25676 1813 25710 1847
rect 25744 1813 25778 1847
rect 25812 1813 25846 1847
rect 25880 1813 25914 1847
rect 25948 1813 25982 1847
rect 26016 1813 26050 1847
rect 26084 1813 26118 1847
rect 26152 1813 26186 1847
rect 26220 1813 26254 1847
rect 26288 1813 26322 1847
rect 26356 1813 26390 1847
rect 26424 1813 26458 1847
rect 26492 1813 26526 1847
rect 26560 1813 26594 1847
rect 26628 1813 26662 1847
rect 26696 1813 26730 1847
rect 26764 1813 26798 1847
rect 26832 1813 26866 1847
rect 26900 1813 26934 1847
rect 26968 1813 27002 1847
rect 27036 1813 27070 1847
rect 27104 1813 27138 1847
rect 27172 1813 27206 1847
rect 27240 1813 27274 1847
rect 27308 1813 27342 1847
rect 27376 1813 27410 1847
rect 27444 1813 27478 1847
rect 27512 1783 27546 1817
rect 27580 1784 27614 1818
rect 27648 1784 27682 1818
rect 2009 1739 2043 1773
rect 2078 1739 2112 1773
rect 2147 1739 2181 1773
rect 2216 1739 2250 1773
rect 2284 1739 2318 1773
rect 2352 1739 2386 1773
rect 2420 1739 2454 1773
rect 2488 1739 2522 1773
rect 2556 1739 2590 1773
rect 2624 1739 2658 1773
rect 2692 1739 2726 1773
rect 2760 1739 2794 1773
rect 2828 1739 2862 1773
rect 2896 1739 2930 1773
rect 2964 1739 2998 1773
rect 3032 1739 3066 1773
rect 3100 1739 3134 1773
rect 3168 1739 3202 1773
rect 3236 1739 3270 1773
rect 3304 1739 3338 1773
rect 3372 1739 3406 1773
rect 3440 1739 3474 1773
rect 3508 1739 3542 1773
rect 3576 1739 3610 1773
rect 3644 1739 3678 1773
rect 3712 1739 3746 1773
rect 3780 1739 3814 1773
rect 3848 1739 3882 1773
rect 3916 1739 3950 1773
rect 3984 1739 4018 1773
rect 4052 1739 4086 1773
rect 4120 1739 4154 1773
rect 4188 1739 4222 1773
rect 4256 1739 4290 1773
rect 4324 1739 4358 1773
rect 4392 1739 4426 1773
rect 4460 1739 4494 1773
rect 4528 1739 4562 1773
rect 4596 1739 4630 1773
rect 4664 1739 4698 1773
rect 4732 1739 4766 1773
rect 4800 1739 4834 1773
rect 4868 1739 4902 1773
rect 4936 1739 4970 1773
rect 5004 1739 5038 1773
rect 5072 1739 5106 1773
rect 5140 1739 5174 1773
rect 5208 1739 5242 1773
rect 5276 1739 5310 1773
rect 5344 1739 5378 1773
rect 5412 1739 5446 1773
rect 5480 1739 5514 1773
rect 5548 1739 5582 1773
rect 5616 1739 5650 1773
rect 5684 1739 5718 1773
rect 5752 1739 5786 1773
rect 5820 1739 5854 1773
rect 5888 1739 5922 1773
rect 5956 1739 5990 1773
rect 6024 1739 6058 1773
rect 6092 1739 6126 1773
rect 6160 1739 6194 1773
rect 6228 1739 6262 1773
rect 6296 1739 6330 1773
rect 6364 1739 6398 1773
rect 6432 1739 6466 1773
rect 6500 1739 6534 1773
rect 6568 1739 6602 1773
rect 6636 1739 6670 1773
rect 6704 1739 6738 1773
rect 6772 1739 6806 1773
rect 6840 1739 6874 1773
rect 6908 1739 6942 1773
rect 6976 1739 7010 1773
rect 7044 1739 7078 1773
rect 7112 1739 7146 1773
rect 7180 1739 7214 1773
rect 7248 1739 7282 1773
rect 7316 1739 7350 1773
rect 7384 1739 7418 1773
rect 7452 1739 7486 1773
rect 7520 1739 7554 1773
rect 7588 1739 7622 1773
rect 7656 1739 7690 1773
rect 7724 1739 7758 1773
rect 7792 1739 7826 1773
rect 7860 1739 7894 1773
rect 7928 1739 7962 1773
rect 7996 1739 8030 1773
rect 8064 1739 8098 1773
rect 8132 1739 8166 1773
rect 8200 1739 8234 1773
rect 8268 1739 8302 1773
rect 8336 1739 8370 1773
rect 8404 1739 8438 1773
rect 8472 1739 8506 1773
rect 8540 1739 8574 1773
rect 8608 1739 8642 1773
rect 8676 1739 8710 1773
rect 8744 1739 8778 1773
rect 8812 1739 8846 1773
rect 8880 1739 8914 1773
rect 8948 1739 8982 1773
rect 9016 1739 9050 1773
rect 9084 1739 9118 1773
rect 9152 1739 9186 1773
rect 9220 1739 9254 1773
rect 9288 1739 9322 1773
rect 9356 1739 9390 1773
rect 9424 1739 9458 1773
rect 9492 1739 9526 1773
rect 9560 1739 9594 1773
rect 9628 1739 9662 1773
rect 9696 1739 9730 1773
rect 9764 1739 9798 1773
rect 9832 1739 9866 1773
rect 9900 1739 9934 1773
rect 9968 1739 10002 1773
rect 10036 1739 10070 1773
rect 10104 1739 10138 1773
rect 10172 1739 10206 1773
rect 10240 1739 10274 1773
rect 10308 1739 10342 1773
rect 10376 1739 10410 1773
rect 10444 1739 10478 1773
rect 10512 1739 10546 1773
rect 10580 1739 10614 1773
rect 10648 1739 10682 1773
rect 10716 1739 10750 1773
rect 10784 1739 10818 1773
rect 10852 1739 10886 1773
rect 10920 1739 10954 1773
rect 10988 1739 11022 1773
rect 11056 1739 11090 1773
rect 11124 1739 11158 1773
rect 11192 1739 11226 1773
rect 11260 1739 11294 1773
rect 11328 1739 11362 1773
rect 11396 1739 11430 1773
rect 11464 1739 11498 1773
rect 11532 1739 11566 1773
rect 11600 1739 11634 1773
rect 11668 1739 11702 1773
rect 11736 1739 11770 1773
rect 11804 1739 11838 1773
rect 11872 1739 11906 1773
rect 11940 1739 11974 1773
rect 12008 1739 12042 1773
rect 12076 1739 12110 1773
rect 12144 1739 12178 1773
rect 12212 1739 12246 1773
rect 12280 1739 12314 1773
rect 12348 1739 12382 1773
rect 12416 1739 12450 1773
rect 12484 1739 12518 1773
rect 12552 1739 12586 1773
rect 12620 1739 12654 1773
rect 12688 1739 12722 1773
rect 12756 1739 12790 1773
rect 12824 1739 12858 1773
rect 12892 1739 12926 1773
rect 12960 1739 12994 1773
rect 13028 1739 13062 1773
rect 13096 1739 13130 1773
rect 13164 1739 13198 1773
rect 13232 1739 13266 1773
rect 13300 1739 13334 1773
rect 13368 1739 13402 1773
rect 13436 1739 13470 1773
rect 13504 1739 13538 1773
rect 13572 1739 13606 1773
rect 13640 1739 13674 1773
rect 13708 1739 13742 1773
rect 13776 1739 13810 1773
rect 13844 1739 13878 1773
rect 13912 1739 13946 1773
rect 13980 1739 14014 1773
rect 14048 1739 14082 1773
rect 14116 1739 14150 1773
rect 14184 1739 14218 1773
rect 14252 1739 14286 1773
rect 14320 1739 14354 1773
rect 14388 1739 14422 1773
rect 14456 1739 14490 1773
rect 14524 1739 14558 1773
rect 14592 1739 14626 1773
rect 14660 1739 14694 1773
rect 14728 1739 14762 1773
rect 14796 1739 14830 1773
rect 14864 1739 14898 1773
rect 14932 1739 14966 1773
rect 15000 1739 15034 1773
rect 15068 1739 15102 1773
rect 15136 1739 15170 1773
rect 15204 1739 15238 1773
rect 15272 1739 15306 1773
rect 15340 1739 15374 1773
rect 15408 1739 15442 1773
rect 15476 1739 15510 1773
rect 15544 1739 15578 1773
rect 15612 1739 15646 1773
rect 15680 1739 15714 1773
rect 15748 1739 15782 1773
rect 15816 1739 15850 1773
rect 15884 1739 15918 1773
rect 15952 1739 15986 1773
rect 16020 1739 16054 1773
rect 16088 1739 16122 1773
rect 16156 1739 16190 1773
rect 16224 1739 16258 1773
rect 16292 1739 16326 1773
rect 16360 1739 16394 1773
rect 16428 1739 16462 1773
rect 16496 1739 16530 1773
rect 16564 1739 16598 1773
rect 16632 1739 16666 1773
rect 16700 1739 16734 1773
rect 16768 1739 16802 1773
rect 16836 1739 16870 1773
rect 16904 1739 16938 1773
rect 16972 1739 17006 1773
rect 17040 1739 17074 1773
rect 17108 1739 17142 1773
rect 17176 1739 17210 1773
rect 17244 1739 17278 1773
rect 17312 1739 17346 1773
rect 17380 1739 17414 1773
rect 17448 1739 17482 1773
rect 17516 1739 17550 1773
rect 17584 1739 17618 1773
rect 17652 1739 17686 1773
rect 17720 1739 17754 1773
rect 17788 1739 17822 1773
rect 17856 1739 17890 1773
rect 17924 1739 17958 1773
rect 17992 1739 18026 1773
rect 18060 1739 18094 1773
rect 18128 1739 18162 1773
rect 18196 1739 18230 1773
rect 18264 1739 18298 1773
rect 18332 1739 18366 1773
rect 18400 1739 18434 1773
rect 18468 1739 18502 1773
rect 18536 1739 18570 1773
rect 18604 1739 18638 1773
rect 18672 1739 18706 1773
rect 18740 1739 18774 1773
rect 18808 1739 18842 1773
rect 18876 1739 18910 1773
rect 18944 1739 18978 1773
rect 19012 1739 19046 1773
rect 19080 1739 19114 1773
rect 19148 1739 19182 1773
rect 19216 1739 19250 1773
rect 19284 1739 19318 1773
rect 19352 1739 19386 1773
rect 19420 1739 19454 1773
rect 19488 1739 19522 1773
rect 19556 1739 19590 1773
rect 19624 1739 19658 1773
rect 19692 1739 19726 1773
rect 19760 1739 19794 1773
rect 19828 1739 19862 1773
rect 19896 1739 19930 1773
rect 19964 1739 19998 1773
rect 20032 1739 20066 1773
rect 20100 1739 20134 1773
rect 20168 1739 20202 1773
rect 20236 1739 20270 1773
rect 20304 1739 20338 1773
rect 20372 1739 20406 1773
rect 20440 1739 20474 1773
rect 20508 1739 20542 1773
rect 20576 1739 20610 1773
rect 20644 1739 20678 1773
rect 20712 1739 20746 1773
rect 20780 1739 20814 1773
rect 20848 1739 20882 1773
rect 20916 1739 20950 1773
rect 20984 1739 21018 1773
rect 21052 1739 21086 1773
rect 21120 1739 21154 1773
rect 21188 1739 21222 1773
rect 21256 1739 21290 1773
rect 21324 1739 21358 1773
rect 21392 1739 21426 1773
rect 21460 1739 21494 1773
rect 21528 1739 21562 1773
rect 21596 1739 21630 1773
rect 21664 1739 21698 1773
rect 21732 1739 21766 1773
rect 21800 1739 21834 1773
rect 21868 1739 21902 1773
rect 21936 1739 21970 1773
rect 22004 1739 22038 1773
rect 22072 1739 22106 1773
rect 22140 1739 22174 1773
rect 22208 1739 22242 1773
rect 22276 1739 22310 1773
rect 22344 1739 22378 1773
rect 22412 1739 22446 1773
rect 22480 1739 22514 1773
rect 22548 1739 22582 1773
rect 22616 1739 22650 1773
rect 22684 1739 22718 1773
rect 22752 1739 22786 1773
rect 22820 1739 22854 1773
rect 22888 1739 22922 1773
rect 22956 1739 22990 1773
rect 23024 1739 23058 1773
rect 23092 1739 23126 1773
rect 23160 1739 23194 1773
rect 23228 1739 23262 1773
rect 23296 1739 23330 1773
rect 23364 1739 23398 1773
rect 23432 1739 23466 1773
rect 23500 1739 23534 1773
rect 23568 1739 23602 1773
rect 23636 1739 23670 1773
rect 23704 1739 23738 1773
rect 23772 1739 23806 1773
rect 23840 1739 23874 1773
rect 23908 1739 23942 1773
rect 23976 1739 24010 1773
rect 24044 1739 24078 1773
rect 24112 1739 24146 1773
rect 24180 1739 24214 1773
rect 24248 1739 24282 1773
rect 24316 1739 24350 1773
rect 24384 1739 24418 1773
rect 24452 1739 24486 1773
rect 24520 1739 24554 1773
rect 24588 1739 24622 1773
rect 24656 1739 24690 1773
rect 24724 1739 24758 1773
rect 24792 1739 24826 1773
rect 24860 1739 24894 1773
rect 24928 1739 24962 1773
rect 24996 1739 25030 1773
rect 25064 1739 25098 1773
rect 25132 1739 25166 1773
rect 25200 1739 25234 1773
rect 25268 1739 25302 1773
rect 25336 1739 25370 1773
rect 25404 1739 25438 1773
rect 25472 1739 25506 1773
rect 25540 1739 25574 1773
rect 25608 1739 25642 1773
rect 25676 1739 25710 1773
rect 25744 1739 25778 1773
rect 25812 1739 25846 1773
rect 25880 1739 25914 1773
rect 25948 1739 25982 1773
rect 26016 1739 26050 1773
rect 26084 1739 26118 1773
rect 26152 1739 26186 1773
rect 26220 1739 26254 1773
rect 26288 1739 26322 1773
rect 26356 1739 26390 1773
rect 26424 1739 26458 1773
rect 26492 1739 26526 1773
rect 26560 1739 26594 1773
rect 26628 1739 26662 1773
rect 26696 1739 26730 1773
rect 26764 1739 26798 1773
rect 26832 1739 26866 1773
rect 26900 1739 26934 1773
rect 26968 1739 27002 1773
rect 27036 1739 27070 1773
rect 27104 1739 27138 1773
rect 27172 1739 27206 1773
rect 27240 1739 27274 1773
rect 27308 1739 27342 1773
rect 27376 1739 27410 1773
rect 27444 1739 27478 1773
rect 27512 1714 27546 1748
rect 27580 1715 27614 1749
rect 27648 1715 27682 1749
rect 2009 1665 2043 1699
rect 2078 1665 2112 1699
rect 2147 1665 2181 1699
rect 2216 1665 2250 1699
rect 2284 1665 2318 1699
rect 2352 1665 2386 1699
rect 2420 1665 2454 1699
rect 2488 1665 2522 1699
rect 2556 1665 2590 1699
rect 2624 1665 2658 1699
rect 2692 1665 2726 1699
rect 2760 1665 2794 1699
rect 2828 1665 2862 1699
rect 2896 1665 2930 1699
rect 2964 1665 2998 1699
rect 3032 1665 3066 1699
rect 3100 1665 3134 1699
rect 3168 1665 3202 1699
rect 3236 1665 3270 1699
rect 3304 1665 3338 1699
rect 3372 1665 3406 1699
rect 3440 1665 3474 1699
rect 3508 1665 3542 1699
rect 3576 1665 3610 1699
rect 3644 1665 3678 1699
rect 3712 1665 3746 1699
rect 3780 1665 3814 1699
rect 3848 1665 3882 1699
rect 3916 1665 3950 1699
rect 3984 1665 4018 1699
rect 4052 1665 4086 1699
rect 4120 1665 4154 1699
rect 4188 1665 4222 1699
rect 4256 1665 4290 1699
rect 4324 1665 4358 1699
rect 4392 1665 4426 1699
rect 4460 1665 4494 1699
rect 4528 1665 4562 1699
rect 4596 1665 4630 1699
rect 4664 1665 4698 1699
rect 4732 1665 4766 1699
rect 4800 1665 4834 1699
rect 4868 1665 4902 1699
rect 4936 1665 4970 1699
rect 5004 1665 5038 1699
rect 5072 1665 5106 1699
rect 5140 1665 5174 1699
rect 5208 1665 5242 1699
rect 5276 1665 5310 1699
rect 5344 1665 5378 1699
rect 5412 1665 5446 1699
rect 5480 1665 5514 1699
rect 5548 1665 5582 1699
rect 5616 1665 5650 1699
rect 5684 1665 5718 1699
rect 5752 1665 5786 1699
rect 5820 1665 5854 1699
rect 5888 1665 5922 1699
rect 5956 1665 5990 1699
rect 6024 1665 6058 1699
rect 6092 1665 6126 1699
rect 6160 1665 6194 1699
rect 6228 1665 6262 1699
rect 6296 1665 6330 1699
rect 6364 1665 6398 1699
rect 6432 1665 6466 1699
rect 6500 1665 6534 1699
rect 6568 1665 6602 1699
rect 6636 1665 6670 1699
rect 6704 1665 6738 1699
rect 6772 1665 6806 1699
rect 6840 1665 6874 1699
rect 6908 1665 6942 1699
rect 6976 1665 7010 1699
rect 7044 1665 7078 1699
rect 7112 1665 7146 1699
rect 7180 1665 7214 1699
rect 7248 1665 7282 1699
rect 7316 1665 7350 1699
rect 7384 1665 7418 1699
rect 7452 1665 7486 1699
rect 7520 1665 7554 1699
rect 7588 1665 7622 1699
rect 7656 1665 7690 1699
rect 7724 1665 7758 1699
rect 7792 1665 7826 1699
rect 7860 1665 7894 1699
rect 7928 1665 7962 1699
rect 7996 1665 8030 1699
rect 8064 1665 8098 1699
rect 8132 1665 8166 1699
rect 8200 1665 8234 1699
rect 8268 1665 8302 1699
rect 8336 1665 8370 1699
rect 8404 1665 8438 1699
rect 8472 1665 8506 1699
rect 8540 1665 8574 1699
rect 8608 1665 8642 1699
rect 8676 1665 8710 1699
rect 8744 1665 8778 1699
rect 8812 1665 8846 1699
rect 8880 1665 8914 1699
rect 8948 1665 8982 1699
rect 9016 1665 9050 1699
rect 9084 1665 9118 1699
rect 9152 1665 9186 1699
rect 9220 1665 9254 1699
rect 9288 1665 9322 1699
rect 9356 1665 9390 1699
rect 9424 1665 9458 1699
rect 9492 1665 9526 1699
rect 9560 1665 9594 1699
rect 9628 1665 9662 1699
rect 9696 1665 9730 1699
rect 9764 1665 9798 1699
rect 9832 1665 9866 1699
rect 9900 1665 9934 1699
rect 9968 1665 10002 1699
rect 10036 1665 10070 1699
rect 10104 1665 10138 1699
rect 10172 1665 10206 1699
rect 10240 1665 10274 1699
rect 10308 1665 10342 1699
rect 10376 1665 10410 1699
rect 10444 1665 10478 1699
rect 10512 1665 10546 1699
rect 10580 1665 10614 1699
rect 10648 1665 10682 1699
rect 10716 1665 10750 1699
rect 10784 1665 10818 1699
rect 10852 1665 10886 1699
rect 10920 1665 10954 1699
rect 10988 1665 11022 1699
rect 11056 1665 11090 1699
rect 11124 1665 11158 1699
rect 11192 1665 11226 1699
rect 11260 1665 11294 1699
rect 11328 1665 11362 1699
rect 11396 1665 11430 1699
rect 11464 1665 11498 1699
rect 11532 1665 11566 1699
rect 11600 1665 11634 1699
rect 11668 1665 11702 1699
rect 11736 1665 11770 1699
rect 11804 1665 11838 1699
rect 11872 1665 11906 1699
rect 11940 1665 11974 1699
rect 12008 1665 12042 1699
rect 12076 1665 12110 1699
rect 12144 1665 12178 1699
rect 12212 1665 12246 1699
rect 12280 1665 12314 1699
rect 12348 1665 12382 1699
rect 12416 1665 12450 1699
rect 12484 1665 12518 1699
rect 12552 1665 12586 1699
rect 12620 1665 12654 1699
rect 12688 1665 12722 1699
rect 12756 1665 12790 1699
rect 12824 1665 12858 1699
rect 12892 1665 12926 1699
rect 12960 1665 12994 1699
rect 13028 1665 13062 1699
rect 13096 1665 13130 1699
rect 13164 1665 13198 1699
rect 13232 1665 13266 1699
rect 13300 1665 13334 1699
rect 13368 1665 13402 1699
rect 13436 1665 13470 1699
rect 13504 1665 13538 1699
rect 13572 1665 13606 1699
rect 13640 1665 13674 1699
rect 13708 1665 13742 1699
rect 13776 1665 13810 1699
rect 13844 1665 13878 1699
rect 13912 1665 13946 1699
rect 13980 1665 14014 1699
rect 14048 1665 14082 1699
rect 14116 1665 14150 1699
rect 14184 1665 14218 1699
rect 14252 1665 14286 1699
rect 14320 1665 14354 1699
rect 14388 1665 14422 1699
rect 14456 1665 14490 1699
rect 14524 1665 14558 1699
rect 14592 1665 14626 1699
rect 14660 1665 14694 1699
rect 14728 1665 14762 1699
rect 14796 1665 14830 1699
rect 14864 1665 14898 1699
rect 14932 1665 14966 1699
rect 15000 1665 15034 1699
rect 15068 1665 15102 1699
rect 15136 1665 15170 1699
rect 15204 1665 15238 1699
rect 15272 1665 15306 1699
rect 15340 1665 15374 1699
rect 15408 1665 15442 1699
rect 15476 1665 15510 1699
rect 15544 1665 15578 1699
rect 15612 1665 15646 1699
rect 15680 1665 15714 1699
rect 15748 1665 15782 1699
rect 15816 1665 15850 1699
rect 15884 1665 15918 1699
rect 15952 1665 15986 1699
rect 16020 1665 16054 1699
rect 16088 1665 16122 1699
rect 16156 1665 16190 1699
rect 16224 1665 16258 1699
rect 16292 1665 16326 1699
rect 16360 1665 16394 1699
rect 16428 1665 16462 1699
rect 16496 1665 16530 1699
rect 16564 1665 16598 1699
rect 16632 1665 16666 1699
rect 16700 1665 16734 1699
rect 16768 1665 16802 1699
rect 16836 1665 16870 1699
rect 16904 1665 16938 1699
rect 16972 1665 17006 1699
rect 17040 1665 17074 1699
rect 17108 1665 17142 1699
rect 17176 1665 17210 1699
rect 17244 1665 17278 1699
rect 17312 1665 17346 1699
rect 17380 1665 17414 1699
rect 17448 1665 17482 1699
rect 17516 1665 17550 1699
rect 17584 1665 17618 1699
rect 17652 1665 17686 1699
rect 17720 1665 17754 1699
rect 17788 1665 17822 1699
rect 17856 1665 17890 1699
rect 17924 1665 17958 1699
rect 17992 1665 18026 1699
rect 18060 1665 18094 1699
rect 18128 1665 18162 1699
rect 18196 1665 18230 1699
rect 18264 1665 18298 1699
rect 18332 1665 18366 1699
rect 18400 1665 18434 1699
rect 18468 1665 18502 1699
rect 18536 1665 18570 1699
rect 18604 1665 18638 1699
rect 18672 1665 18706 1699
rect 18740 1665 18774 1699
rect 18808 1665 18842 1699
rect 18876 1665 18910 1699
rect 18944 1665 18978 1699
rect 19012 1665 19046 1699
rect 19080 1665 19114 1699
rect 19148 1665 19182 1699
rect 19216 1665 19250 1699
rect 19284 1665 19318 1699
rect 19352 1665 19386 1699
rect 19420 1665 19454 1699
rect 19488 1665 19522 1699
rect 19556 1665 19590 1699
rect 19624 1665 19658 1699
rect 19692 1665 19726 1699
rect 19760 1665 19794 1699
rect 19828 1665 19862 1699
rect 19896 1665 19930 1699
rect 19964 1665 19998 1699
rect 20032 1665 20066 1699
rect 20100 1665 20134 1699
rect 20168 1665 20202 1699
rect 20236 1665 20270 1699
rect 20304 1665 20338 1699
rect 20372 1665 20406 1699
rect 20440 1665 20474 1699
rect 20508 1665 20542 1699
rect 20576 1665 20610 1699
rect 20644 1665 20678 1699
rect 20712 1665 20746 1699
rect 20780 1665 20814 1699
rect 20848 1665 20882 1699
rect 20916 1665 20950 1699
rect 20984 1665 21018 1699
rect 21052 1665 21086 1699
rect 21120 1665 21154 1699
rect 21188 1665 21222 1699
rect 21256 1665 21290 1699
rect 21324 1665 21358 1699
rect 21392 1665 21426 1699
rect 21460 1665 21494 1699
rect 21528 1665 21562 1699
rect 21596 1665 21630 1699
rect 21664 1665 21698 1699
rect 21732 1665 21766 1699
rect 21800 1665 21834 1699
rect 21868 1665 21902 1699
rect 21936 1665 21970 1699
rect 22004 1665 22038 1699
rect 22072 1665 22106 1699
rect 22140 1665 22174 1699
rect 22208 1665 22242 1699
rect 22276 1665 22310 1699
rect 22344 1665 22378 1699
rect 22412 1665 22446 1699
rect 22480 1665 22514 1699
rect 22548 1665 22582 1699
rect 22616 1665 22650 1699
rect 22684 1665 22718 1699
rect 22752 1665 22786 1699
rect 22820 1665 22854 1699
rect 22888 1665 22922 1699
rect 22956 1665 22990 1699
rect 23024 1665 23058 1699
rect 23092 1665 23126 1699
rect 23160 1665 23194 1699
rect 23228 1665 23262 1699
rect 23296 1665 23330 1699
rect 23364 1665 23398 1699
rect 23432 1665 23466 1699
rect 23500 1665 23534 1699
rect 23568 1665 23602 1699
rect 23636 1665 23670 1699
rect 23704 1665 23738 1699
rect 23772 1665 23806 1699
rect 23840 1665 23874 1699
rect 23908 1665 23942 1699
rect 23976 1665 24010 1699
rect 24044 1665 24078 1699
rect 24112 1665 24146 1699
rect 24180 1665 24214 1699
rect 24248 1665 24282 1699
rect 24316 1665 24350 1699
rect 24384 1665 24418 1699
rect 24452 1665 24486 1699
rect 24520 1665 24554 1699
rect 24588 1665 24622 1699
rect 24656 1665 24690 1699
rect 24724 1665 24758 1699
rect 24792 1665 24826 1699
rect 24860 1665 24894 1699
rect 24928 1665 24962 1699
rect 24996 1665 25030 1699
rect 25064 1665 25098 1699
rect 25132 1665 25166 1699
rect 25200 1665 25234 1699
rect 25268 1665 25302 1699
rect 25336 1665 25370 1699
rect 25404 1665 25438 1699
rect 25472 1665 25506 1699
rect 25540 1665 25574 1699
rect 25608 1665 25642 1699
rect 25676 1665 25710 1699
rect 25744 1665 25778 1699
rect 25812 1665 25846 1699
rect 25880 1665 25914 1699
rect 25948 1665 25982 1699
rect 26016 1665 26050 1699
rect 26084 1665 26118 1699
rect 26152 1665 26186 1699
rect 26220 1665 26254 1699
rect 26288 1665 26322 1699
rect 26356 1665 26390 1699
rect 26424 1665 26458 1699
rect 26492 1665 26526 1699
rect 26560 1665 26594 1699
rect 26628 1665 26662 1699
rect 26696 1665 26730 1699
rect 26764 1665 26798 1699
rect 26832 1665 26866 1699
rect 26900 1665 26934 1699
rect 26968 1665 27002 1699
rect 27036 1665 27070 1699
rect 27104 1665 27138 1699
rect 27172 1665 27206 1699
rect 27240 1665 27274 1699
rect 27308 1665 27342 1699
rect 27376 1665 27410 1699
rect 27444 1665 27478 1699
rect 27512 1645 27546 1679
rect 27580 1646 27614 1680
rect 27648 1646 27682 1680
rect 2009 1591 2043 1625
rect 2078 1591 2112 1625
rect 2147 1591 2181 1625
rect 2216 1591 2250 1625
rect 2284 1591 2318 1625
rect 2352 1591 2386 1625
rect 2420 1591 2454 1625
rect 2488 1591 2522 1625
rect 2556 1591 2590 1625
rect 2624 1591 2658 1625
rect 2692 1591 2726 1625
rect 2760 1591 2794 1625
rect 2828 1591 2862 1625
rect 2896 1591 2930 1625
rect 2964 1591 2998 1625
rect 3032 1591 3066 1625
rect 3100 1591 3134 1625
rect 3168 1591 3202 1625
rect 3236 1591 3270 1625
rect 3304 1591 3338 1625
rect 3372 1591 3406 1625
rect 3440 1591 3474 1625
rect 3508 1591 3542 1625
rect 3576 1591 3610 1625
rect 3644 1591 3678 1625
rect 3712 1591 3746 1625
rect 3780 1591 3814 1625
rect 3848 1591 3882 1625
rect 3916 1591 3950 1625
rect 3984 1591 4018 1625
rect 4052 1591 4086 1625
rect 4120 1591 4154 1625
rect 4188 1591 4222 1625
rect 4256 1591 4290 1625
rect 4324 1591 4358 1625
rect 4392 1591 4426 1625
rect 4460 1591 4494 1625
rect 4528 1591 4562 1625
rect 4596 1591 4630 1625
rect 4664 1591 4698 1625
rect 4732 1591 4766 1625
rect 4800 1591 4834 1625
rect 4868 1591 4902 1625
rect 4936 1591 4970 1625
rect 5004 1591 5038 1625
rect 5072 1591 5106 1625
rect 5140 1591 5174 1625
rect 5208 1591 5242 1625
rect 5276 1591 5310 1625
rect 5344 1591 5378 1625
rect 5412 1591 5446 1625
rect 5480 1591 5514 1625
rect 5548 1591 5582 1625
rect 5616 1591 5650 1625
rect 5684 1591 5718 1625
rect 5752 1591 5786 1625
rect 5820 1591 5854 1625
rect 5888 1591 5922 1625
rect 5956 1591 5990 1625
rect 6024 1591 6058 1625
rect 6092 1591 6126 1625
rect 6160 1591 6194 1625
rect 6228 1591 6262 1625
rect 6296 1591 6330 1625
rect 6364 1591 6398 1625
rect 6432 1591 6466 1625
rect 6500 1591 6534 1625
rect 6568 1591 6602 1625
rect 6636 1591 6670 1625
rect 6704 1591 6738 1625
rect 6772 1591 6806 1625
rect 6840 1591 6874 1625
rect 6908 1591 6942 1625
rect 6976 1591 7010 1625
rect 7044 1591 7078 1625
rect 7112 1591 7146 1625
rect 7180 1591 7214 1625
rect 7248 1591 7282 1625
rect 7316 1591 7350 1625
rect 7384 1591 7418 1625
rect 7452 1591 7486 1625
rect 7520 1591 7554 1625
rect 7588 1591 7622 1625
rect 7656 1591 7690 1625
rect 7724 1591 7758 1625
rect 7792 1591 7826 1625
rect 7860 1591 7894 1625
rect 7928 1591 7962 1625
rect 7996 1591 8030 1625
rect 8064 1591 8098 1625
rect 8132 1591 8166 1625
rect 8200 1591 8234 1625
rect 8268 1591 8302 1625
rect 8336 1591 8370 1625
rect 8404 1591 8438 1625
rect 8472 1591 8506 1625
rect 8540 1591 8574 1625
rect 8608 1591 8642 1625
rect 8676 1591 8710 1625
rect 8744 1591 8778 1625
rect 8812 1591 8846 1625
rect 8880 1591 8914 1625
rect 8948 1591 8982 1625
rect 9016 1591 9050 1625
rect 9084 1591 9118 1625
rect 9152 1591 9186 1625
rect 9220 1591 9254 1625
rect 9288 1591 9322 1625
rect 9356 1591 9390 1625
rect 9424 1591 9458 1625
rect 9492 1591 9526 1625
rect 9560 1591 9594 1625
rect 9628 1591 9662 1625
rect 9696 1591 9730 1625
rect 9764 1591 9798 1625
rect 9832 1591 9866 1625
rect 9900 1591 9934 1625
rect 9968 1591 10002 1625
rect 10036 1591 10070 1625
rect 10104 1591 10138 1625
rect 10172 1591 10206 1625
rect 10240 1591 10274 1625
rect 10308 1591 10342 1625
rect 10376 1591 10410 1625
rect 10444 1591 10478 1625
rect 10512 1591 10546 1625
rect 10580 1591 10614 1625
rect 10648 1591 10682 1625
rect 10716 1591 10750 1625
rect 10784 1591 10818 1625
rect 10852 1591 10886 1625
rect 10920 1591 10954 1625
rect 10988 1591 11022 1625
rect 11056 1591 11090 1625
rect 11124 1591 11158 1625
rect 11192 1591 11226 1625
rect 11260 1591 11294 1625
rect 11328 1591 11362 1625
rect 11396 1591 11430 1625
rect 11464 1591 11498 1625
rect 11532 1591 11566 1625
rect 11600 1591 11634 1625
rect 11668 1591 11702 1625
rect 11736 1591 11770 1625
rect 11804 1591 11838 1625
rect 11872 1591 11906 1625
rect 11940 1591 11974 1625
rect 12008 1591 12042 1625
rect 12076 1591 12110 1625
rect 12144 1591 12178 1625
rect 12212 1591 12246 1625
rect 12280 1591 12314 1625
rect 12348 1591 12382 1625
rect 12416 1591 12450 1625
rect 12484 1591 12518 1625
rect 12552 1591 12586 1625
rect 12620 1591 12654 1625
rect 12688 1591 12722 1625
rect 12756 1591 12790 1625
rect 12824 1591 12858 1625
rect 12892 1591 12926 1625
rect 12960 1591 12994 1625
rect 13028 1591 13062 1625
rect 13096 1591 13130 1625
rect 13164 1591 13198 1625
rect 13232 1591 13266 1625
rect 13300 1591 13334 1625
rect 13368 1591 13402 1625
rect 13436 1591 13470 1625
rect 13504 1591 13538 1625
rect 13572 1591 13606 1625
rect 13640 1591 13674 1625
rect 13708 1591 13742 1625
rect 13776 1591 13810 1625
rect 13844 1591 13878 1625
rect 13912 1591 13946 1625
rect 13980 1591 14014 1625
rect 14048 1591 14082 1625
rect 14116 1591 14150 1625
rect 14184 1591 14218 1625
rect 14252 1591 14286 1625
rect 14320 1591 14354 1625
rect 14388 1591 14422 1625
rect 14456 1591 14490 1625
rect 14524 1591 14558 1625
rect 14592 1591 14626 1625
rect 14660 1591 14694 1625
rect 14728 1591 14762 1625
rect 14796 1591 14830 1625
rect 14864 1591 14898 1625
rect 14932 1591 14966 1625
rect 15000 1591 15034 1625
rect 15068 1591 15102 1625
rect 15136 1591 15170 1625
rect 15204 1591 15238 1625
rect 15272 1591 15306 1625
rect 15340 1591 15374 1625
rect 15408 1591 15442 1625
rect 15476 1591 15510 1625
rect 15544 1591 15578 1625
rect 15612 1591 15646 1625
rect 15680 1591 15714 1625
rect 15748 1591 15782 1625
rect 15816 1591 15850 1625
rect 15884 1591 15918 1625
rect 15952 1591 15986 1625
rect 16020 1591 16054 1625
rect 16088 1591 16122 1625
rect 16156 1591 16190 1625
rect 16224 1591 16258 1625
rect 16292 1591 16326 1625
rect 16360 1591 16394 1625
rect 16428 1591 16462 1625
rect 16496 1591 16530 1625
rect 16564 1591 16598 1625
rect 16632 1591 16666 1625
rect 16700 1591 16734 1625
rect 16768 1591 16802 1625
rect 16836 1591 16870 1625
rect 16904 1591 16938 1625
rect 16972 1591 17006 1625
rect 17040 1591 17074 1625
rect 17108 1591 17142 1625
rect 17176 1591 17210 1625
rect 17244 1591 17278 1625
rect 17312 1591 17346 1625
rect 17380 1591 17414 1625
rect 17448 1591 17482 1625
rect 17516 1591 17550 1625
rect 17584 1591 17618 1625
rect 17652 1591 17686 1625
rect 17720 1591 17754 1625
rect 17788 1591 17822 1625
rect 17856 1591 17890 1625
rect 17924 1591 17958 1625
rect 17992 1591 18026 1625
rect 18060 1591 18094 1625
rect 18128 1591 18162 1625
rect 18196 1591 18230 1625
rect 18264 1591 18298 1625
rect 18332 1591 18366 1625
rect 18400 1591 18434 1625
rect 18468 1591 18502 1625
rect 18536 1591 18570 1625
rect 18604 1591 18638 1625
rect 18672 1591 18706 1625
rect 18740 1591 18774 1625
rect 18808 1591 18842 1625
rect 18876 1591 18910 1625
rect 18944 1591 18978 1625
rect 19012 1591 19046 1625
rect 19080 1591 19114 1625
rect 19148 1591 19182 1625
rect 19216 1591 19250 1625
rect 19284 1591 19318 1625
rect 19352 1591 19386 1625
rect 19420 1591 19454 1625
rect 19488 1591 19522 1625
rect 19556 1591 19590 1625
rect 19624 1591 19658 1625
rect 19692 1591 19726 1625
rect 19760 1591 19794 1625
rect 19828 1591 19862 1625
rect 19896 1591 19930 1625
rect 19964 1591 19998 1625
rect 20032 1591 20066 1625
rect 20100 1591 20134 1625
rect 20168 1591 20202 1625
rect 20236 1591 20270 1625
rect 20304 1591 20338 1625
rect 20372 1591 20406 1625
rect 20440 1591 20474 1625
rect 20508 1591 20542 1625
rect 20576 1591 20610 1625
rect 20644 1591 20678 1625
rect 20712 1591 20746 1625
rect 20780 1591 20814 1625
rect 20848 1591 20882 1625
rect 20916 1591 20950 1625
rect 20984 1591 21018 1625
rect 21052 1591 21086 1625
rect 21120 1591 21154 1625
rect 21188 1591 21222 1625
rect 21256 1591 21290 1625
rect 21324 1591 21358 1625
rect 21392 1591 21426 1625
rect 21460 1591 21494 1625
rect 21528 1591 21562 1625
rect 21596 1591 21630 1625
rect 21664 1591 21698 1625
rect 21732 1591 21766 1625
rect 21800 1591 21834 1625
rect 21868 1591 21902 1625
rect 21936 1591 21970 1625
rect 22004 1591 22038 1625
rect 22072 1591 22106 1625
rect 22140 1591 22174 1625
rect 22208 1591 22242 1625
rect 22276 1591 22310 1625
rect 22344 1591 22378 1625
rect 22412 1591 22446 1625
rect 22480 1591 22514 1625
rect 22548 1591 22582 1625
rect 22616 1591 22650 1625
rect 22684 1591 22718 1625
rect 22752 1591 22786 1625
rect 22820 1591 22854 1625
rect 22888 1591 22922 1625
rect 22956 1591 22990 1625
rect 23024 1591 23058 1625
rect 23092 1591 23126 1625
rect 23160 1591 23194 1625
rect 23228 1591 23262 1625
rect 23296 1591 23330 1625
rect 23364 1591 23398 1625
rect 23432 1591 23466 1625
rect 23500 1591 23534 1625
rect 23568 1591 23602 1625
rect 23636 1591 23670 1625
rect 23704 1591 23738 1625
rect 23772 1591 23806 1625
rect 23840 1591 23874 1625
rect 23908 1591 23942 1625
rect 23976 1591 24010 1625
rect 24044 1591 24078 1625
rect 24112 1591 24146 1625
rect 24180 1591 24214 1625
rect 24248 1591 24282 1625
rect 24316 1591 24350 1625
rect 24384 1591 24418 1625
rect 24452 1591 24486 1625
rect 24520 1591 24554 1625
rect 24588 1591 24622 1625
rect 24656 1591 24690 1625
rect 24724 1591 24758 1625
rect 24792 1591 24826 1625
rect 24860 1591 24894 1625
rect 24928 1591 24962 1625
rect 24996 1591 25030 1625
rect 25064 1591 25098 1625
rect 25132 1591 25166 1625
rect 25200 1591 25234 1625
rect 25268 1591 25302 1625
rect 25336 1591 25370 1625
rect 25404 1591 25438 1625
rect 25472 1591 25506 1625
rect 25540 1591 25574 1625
rect 25608 1591 25642 1625
rect 25676 1591 25710 1625
rect 25744 1591 25778 1625
rect 25812 1591 25846 1625
rect 25880 1591 25914 1625
rect 25948 1591 25982 1625
rect 26016 1591 26050 1625
rect 26084 1591 26118 1625
rect 26152 1591 26186 1625
rect 26220 1591 26254 1625
rect 26288 1591 26322 1625
rect 26356 1591 26390 1625
rect 26424 1591 26458 1625
rect 26492 1591 26526 1625
rect 26560 1591 26594 1625
rect 26628 1591 26662 1625
rect 26696 1591 26730 1625
rect 26764 1591 26798 1625
rect 26832 1591 26866 1625
rect 26900 1591 26934 1625
rect 26968 1591 27002 1625
rect 27036 1591 27070 1625
rect 27104 1591 27138 1625
rect 27172 1591 27206 1625
rect 27240 1591 27274 1625
rect 27308 1591 27342 1625
rect 27376 1591 27410 1625
rect 27444 1591 27478 1625
rect 27512 1576 27546 1610
rect 27580 1577 27614 1611
rect 27648 1577 27682 1611
rect 2009 1517 2043 1551
rect 2078 1517 2112 1551
rect 2147 1517 2181 1551
rect 2216 1517 2250 1551
rect 2284 1517 2318 1551
rect 2352 1517 2386 1551
rect 2420 1517 2454 1551
rect 2488 1517 2522 1551
rect 2556 1517 2590 1551
rect 2624 1517 2658 1551
rect 2692 1517 2726 1551
rect 2760 1517 2794 1551
rect 2828 1517 2862 1551
rect 2896 1517 2930 1551
rect 2964 1517 2998 1551
rect 3032 1517 3066 1551
rect 3100 1517 3134 1551
rect 3168 1517 3202 1551
rect 3236 1517 3270 1551
rect 3304 1517 3338 1551
rect 3372 1517 3406 1551
rect 3440 1517 3474 1551
rect 3508 1517 3542 1551
rect 3576 1517 3610 1551
rect 3644 1517 3678 1551
rect 3712 1517 3746 1551
rect 3780 1517 3814 1551
rect 3848 1517 3882 1551
rect 3916 1517 3950 1551
rect 3984 1517 4018 1551
rect 4052 1517 4086 1551
rect 4120 1517 4154 1551
rect 4188 1517 4222 1551
rect 4256 1517 4290 1551
rect 4324 1517 4358 1551
rect 4392 1517 4426 1551
rect 4460 1517 4494 1551
rect 4528 1517 4562 1551
rect 4596 1517 4630 1551
rect 4664 1517 4698 1551
rect 4732 1517 4766 1551
rect 4800 1517 4834 1551
rect 4868 1517 4902 1551
rect 4936 1517 4970 1551
rect 5004 1517 5038 1551
rect 5072 1517 5106 1551
rect 5140 1517 5174 1551
rect 5208 1517 5242 1551
rect 5276 1517 5310 1551
rect 5344 1517 5378 1551
rect 5412 1517 5446 1551
rect 5480 1517 5514 1551
rect 5548 1517 5582 1551
rect 5616 1517 5650 1551
rect 5684 1517 5718 1551
rect 5752 1517 5786 1551
rect 5820 1517 5854 1551
rect 5888 1517 5922 1551
rect 5956 1517 5990 1551
rect 6024 1517 6058 1551
rect 6092 1517 6126 1551
rect 6160 1517 6194 1551
rect 6228 1517 6262 1551
rect 6296 1517 6330 1551
rect 6364 1517 6398 1551
rect 6432 1517 6466 1551
rect 6500 1517 6534 1551
rect 6568 1517 6602 1551
rect 6636 1517 6670 1551
rect 6704 1517 6738 1551
rect 6772 1517 6806 1551
rect 6840 1517 6874 1551
rect 6908 1517 6942 1551
rect 6976 1517 7010 1551
rect 7044 1517 7078 1551
rect 7112 1517 7146 1551
rect 7180 1517 7214 1551
rect 7248 1517 7282 1551
rect 7316 1517 7350 1551
rect 7384 1517 7418 1551
rect 7452 1517 7486 1551
rect 7520 1517 7554 1551
rect 7588 1517 7622 1551
rect 7656 1517 7690 1551
rect 7724 1517 7758 1551
rect 7792 1517 7826 1551
rect 7860 1517 7894 1551
rect 7928 1517 7962 1551
rect 7996 1517 8030 1551
rect 8064 1517 8098 1551
rect 8132 1517 8166 1551
rect 8200 1517 8234 1551
rect 8268 1517 8302 1551
rect 8336 1517 8370 1551
rect 8404 1517 8438 1551
rect 8472 1517 8506 1551
rect 8540 1517 8574 1551
rect 8608 1517 8642 1551
rect 8676 1517 8710 1551
rect 8744 1517 8778 1551
rect 8812 1517 8846 1551
rect 8880 1517 8914 1551
rect 8948 1517 8982 1551
rect 9016 1517 9050 1551
rect 9084 1517 9118 1551
rect 9152 1517 9186 1551
rect 9220 1517 9254 1551
rect 9288 1517 9322 1551
rect 9356 1517 9390 1551
rect 9424 1517 9458 1551
rect 9492 1517 9526 1551
rect 9560 1517 9594 1551
rect 9628 1517 9662 1551
rect 9696 1517 9730 1551
rect 9764 1517 9798 1551
rect 9832 1517 9866 1551
rect 9900 1517 9934 1551
rect 9968 1517 10002 1551
rect 10036 1517 10070 1551
rect 10104 1517 10138 1551
rect 10172 1517 10206 1551
rect 10240 1517 10274 1551
rect 10308 1517 10342 1551
rect 10376 1517 10410 1551
rect 10444 1517 10478 1551
rect 10512 1517 10546 1551
rect 10580 1517 10614 1551
rect 10648 1517 10682 1551
rect 10716 1517 10750 1551
rect 10784 1517 10818 1551
rect 10852 1517 10886 1551
rect 10920 1517 10954 1551
rect 10988 1517 11022 1551
rect 11056 1517 11090 1551
rect 11124 1517 11158 1551
rect 11192 1517 11226 1551
rect 11260 1517 11294 1551
rect 11328 1517 11362 1551
rect 11396 1517 11430 1551
rect 11464 1517 11498 1551
rect 11532 1517 11566 1551
rect 11600 1517 11634 1551
rect 11668 1517 11702 1551
rect 11736 1517 11770 1551
rect 11804 1517 11838 1551
rect 11872 1517 11906 1551
rect 11940 1517 11974 1551
rect 12008 1517 12042 1551
rect 12076 1517 12110 1551
rect 12144 1517 12178 1551
rect 12212 1517 12246 1551
rect 12280 1517 12314 1551
rect 12348 1517 12382 1551
rect 12416 1517 12450 1551
rect 12484 1517 12518 1551
rect 12552 1517 12586 1551
rect 12620 1517 12654 1551
rect 12688 1517 12722 1551
rect 12756 1517 12790 1551
rect 12824 1517 12858 1551
rect 12892 1517 12926 1551
rect 12960 1517 12994 1551
rect 13028 1517 13062 1551
rect 13096 1517 13130 1551
rect 13164 1517 13198 1551
rect 13232 1517 13266 1551
rect 13300 1517 13334 1551
rect 13368 1517 13402 1551
rect 13436 1517 13470 1551
rect 13504 1517 13538 1551
rect 13572 1517 13606 1551
rect 13640 1517 13674 1551
rect 13708 1517 13742 1551
rect 13776 1517 13810 1551
rect 13844 1517 13878 1551
rect 13912 1517 13946 1551
rect 13980 1517 14014 1551
rect 14048 1517 14082 1551
rect 14116 1517 14150 1551
rect 14184 1517 14218 1551
rect 14252 1517 14286 1551
rect 14320 1517 14354 1551
rect 14388 1517 14422 1551
rect 14456 1517 14490 1551
rect 14524 1517 14558 1551
rect 14592 1517 14626 1551
rect 14660 1517 14694 1551
rect 14728 1517 14762 1551
rect 14796 1517 14830 1551
rect 14864 1517 14898 1551
rect 14932 1517 14966 1551
rect 15000 1517 15034 1551
rect 15068 1517 15102 1551
rect 15136 1517 15170 1551
rect 15204 1517 15238 1551
rect 15272 1517 15306 1551
rect 15340 1517 15374 1551
rect 15408 1517 15442 1551
rect 15476 1517 15510 1551
rect 15544 1517 15578 1551
rect 15612 1517 15646 1551
rect 15680 1517 15714 1551
rect 15748 1517 15782 1551
rect 15816 1517 15850 1551
rect 15884 1517 15918 1551
rect 15952 1517 15986 1551
rect 16020 1517 16054 1551
rect 16088 1517 16122 1551
rect 16156 1517 16190 1551
rect 16224 1517 16258 1551
rect 16292 1517 16326 1551
rect 16360 1517 16394 1551
rect 16428 1517 16462 1551
rect 16496 1517 16530 1551
rect 16564 1517 16598 1551
rect 16632 1517 16666 1551
rect 16700 1517 16734 1551
rect 16768 1517 16802 1551
rect 16836 1517 16870 1551
rect 16904 1517 16938 1551
rect 16972 1517 17006 1551
rect 17040 1517 17074 1551
rect 17108 1517 17142 1551
rect 17176 1517 17210 1551
rect 17244 1517 17278 1551
rect 17312 1517 17346 1551
rect 17380 1517 17414 1551
rect 17448 1517 17482 1551
rect 17516 1517 17550 1551
rect 17584 1517 17618 1551
rect 17652 1517 17686 1551
rect 17720 1517 17754 1551
rect 17788 1517 17822 1551
rect 17856 1517 17890 1551
rect 17924 1517 17958 1551
rect 17992 1517 18026 1551
rect 18060 1517 18094 1551
rect 18128 1517 18162 1551
rect 18196 1517 18230 1551
rect 18264 1517 18298 1551
rect 18332 1517 18366 1551
rect 18400 1517 18434 1551
rect 18468 1517 18502 1551
rect 18536 1517 18570 1551
rect 18604 1517 18638 1551
rect 18672 1517 18706 1551
rect 18740 1517 18774 1551
rect 18808 1517 18842 1551
rect 18876 1517 18910 1551
rect 18944 1517 18978 1551
rect 19012 1517 19046 1551
rect 19080 1517 19114 1551
rect 19148 1517 19182 1551
rect 19216 1517 19250 1551
rect 19284 1517 19318 1551
rect 19352 1517 19386 1551
rect 19420 1517 19454 1551
rect 19488 1517 19522 1551
rect 19556 1517 19590 1551
rect 19624 1517 19658 1551
rect 19692 1517 19726 1551
rect 19760 1517 19794 1551
rect 19828 1517 19862 1551
rect 19896 1517 19930 1551
rect 19964 1517 19998 1551
rect 20032 1517 20066 1551
rect 20100 1517 20134 1551
rect 20168 1517 20202 1551
rect 20236 1517 20270 1551
rect 20304 1517 20338 1551
rect 20372 1517 20406 1551
rect 20440 1517 20474 1551
rect 20508 1517 20542 1551
rect 20576 1517 20610 1551
rect 20644 1517 20678 1551
rect 20712 1517 20746 1551
rect 20780 1517 20814 1551
rect 20848 1517 20882 1551
rect 20916 1517 20950 1551
rect 20984 1517 21018 1551
rect 21052 1517 21086 1551
rect 21120 1517 21154 1551
rect 21188 1517 21222 1551
rect 21256 1517 21290 1551
rect 21324 1517 21358 1551
rect 21392 1517 21426 1551
rect 21460 1517 21494 1551
rect 21528 1517 21562 1551
rect 21596 1517 21630 1551
rect 21664 1517 21698 1551
rect 21732 1517 21766 1551
rect 21800 1517 21834 1551
rect 21868 1517 21902 1551
rect 21936 1517 21970 1551
rect 22004 1517 22038 1551
rect 22072 1517 22106 1551
rect 22140 1517 22174 1551
rect 22208 1517 22242 1551
rect 22276 1517 22310 1551
rect 22344 1517 22378 1551
rect 22412 1517 22446 1551
rect 22480 1517 22514 1551
rect 22548 1517 22582 1551
rect 22616 1517 22650 1551
rect 22684 1517 22718 1551
rect 22752 1517 22786 1551
rect 22820 1517 22854 1551
rect 22888 1517 22922 1551
rect 22956 1517 22990 1551
rect 23024 1517 23058 1551
rect 23092 1517 23126 1551
rect 23160 1517 23194 1551
rect 23228 1517 23262 1551
rect 23296 1517 23330 1551
rect 23364 1517 23398 1551
rect 23432 1517 23466 1551
rect 23500 1517 23534 1551
rect 23568 1517 23602 1551
rect 23636 1517 23670 1551
rect 23704 1517 23738 1551
rect 23772 1517 23806 1551
rect 23840 1517 23874 1551
rect 23908 1517 23942 1551
rect 23976 1517 24010 1551
rect 24044 1517 24078 1551
rect 24112 1517 24146 1551
rect 24180 1517 24214 1551
rect 24248 1517 24282 1551
rect 24316 1517 24350 1551
rect 24384 1517 24418 1551
rect 24452 1517 24486 1551
rect 24520 1517 24554 1551
rect 24588 1517 24622 1551
rect 24656 1517 24690 1551
rect 24724 1517 24758 1551
rect 24792 1517 24826 1551
rect 24860 1517 24894 1551
rect 24928 1517 24962 1551
rect 24996 1517 25030 1551
rect 25064 1517 25098 1551
rect 25132 1517 25166 1551
rect 25200 1517 25234 1551
rect 25268 1517 25302 1551
rect 25336 1517 25370 1551
rect 25404 1517 25438 1551
rect 25472 1517 25506 1551
rect 25540 1517 25574 1551
rect 25608 1517 25642 1551
rect 25676 1517 25710 1551
rect 25744 1517 25778 1551
rect 25812 1517 25846 1551
rect 25880 1517 25914 1551
rect 25948 1517 25982 1551
rect 26016 1517 26050 1551
rect 26084 1517 26118 1551
rect 26152 1517 26186 1551
rect 26220 1517 26254 1551
rect 26288 1517 26322 1551
rect 26356 1517 26390 1551
rect 26424 1517 26458 1551
rect 26492 1517 26526 1551
rect 26560 1517 26594 1551
rect 26628 1517 26662 1551
rect 26696 1517 26730 1551
rect 26764 1517 26798 1551
rect 26832 1517 26866 1551
rect 26900 1517 26934 1551
rect 26968 1517 27002 1551
rect 27036 1517 27070 1551
rect 27104 1517 27138 1551
rect 27172 1517 27206 1551
rect 27240 1517 27274 1551
rect 27308 1517 27342 1551
rect 27376 1517 27410 1551
rect 27444 1517 27478 1551
rect 27512 1507 27546 1541
rect 27580 1508 27614 1542
rect 27648 1508 27682 1542
rect 2010 1438 2044 1472
rect 2079 1438 2113 1472
rect 1805 1370 1907 1438
rect 2148 1404 27546 1472
rect 27580 1439 27614 1473
rect 27648 1439 27682 1473
rect 1942 1370 1976 1404
rect 2011 1370 2045 1404
rect 1873 1302 1907 1336
rect 1942 1302 1976 1336
rect 2011 1302 2045 1336
rect 2080 1302 27614 1404
rect 27648 1370 27682 1404
<< mvnsubdiffcont >>
rect 1480 9246 1514 9280
rect 1357 9144 1459 9212
rect 1548 9178 27966 9280
rect 1357 978 1527 9144
rect 1616 9110 27966 9178
rect 2273 8424 2307 8458
rect 2191 8322 2293 8390
rect 2341 8356 27195 8458
rect 2191 2916 2361 8322
rect 2409 8288 27127 8356
rect 27229 8323 27263 8357
rect 2191 2484 2361 2790
rect 2191 2416 2293 2484
rect 27161 8221 27263 8289
rect 2191 2348 2225 2382
rect 2327 2373 27045 2441
rect 27093 2407 27263 8221
rect 2259 2271 27113 2373
rect 27161 2339 27263 2407
rect 27147 2271 27181 2305
rect 27915 978 28085 9036
rect 1357 882 1595 978
rect 1630 944 1664 978
rect 1699 944 1733 978
rect 1768 944 1802 978
rect 1837 944 1871 978
rect 1906 944 1940 978
rect 1975 944 2009 978
rect 2044 944 2078 978
rect 2113 944 2147 978
rect 2182 944 2216 978
rect 2251 944 2285 978
rect 2320 944 2354 978
rect 2389 944 2423 978
rect 2458 944 2492 978
rect 2527 944 2561 978
rect 2596 944 2630 978
rect 2665 944 2699 978
rect 2734 944 2768 978
rect 2803 944 2837 978
rect 2872 944 2906 978
rect 2941 944 2975 978
rect 3010 944 3044 978
rect 3079 944 3113 978
rect 3148 944 3182 978
rect 3217 944 3251 978
rect 3286 944 3320 978
rect 3355 944 3389 978
rect 3424 944 3458 978
rect 3493 944 3527 978
rect 3562 944 3596 978
rect 3631 944 3665 978
rect 3700 944 3734 978
rect 3769 944 3803 978
rect 3838 944 3872 978
rect 3907 944 3941 978
rect 3976 944 4010 978
rect 4045 944 4079 978
rect 4114 944 4148 978
rect 1561 876 1595 882
rect 1630 876 1664 910
rect 1699 876 1733 910
rect 1768 876 1802 910
rect 1837 876 1871 910
rect 1906 876 1940 910
rect 1975 876 2009 910
rect 2044 876 2078 910
rect 2113 876 2147 910
rect 2182 876 2216 910
rect 2251 876 2285 910
rect 2320 876 2354 910
rect 2389 876 2423 910
rect 2458 876 2492 910
rect 2527 876 2561 910
rect 2596 876 2630 910
rect 2665 876 2699 910
rect 2734 876 2768 910
rect 2803 876 2837 910
rect 2872 876 2906 910
rect 2941 876 2975 910
rect 3010 876 3044 910
rect 3079 876 3113 910
rect 3148 876 3182 910
rect 3217 876 3251 910
rect 3286 876 3320 910
rect 3355 876 3389 910
rect 3424 876 3458 910
rect 3493 876 3527 910
rect 3562 876 3596 910
rect 3631 876 3665 910
rect 3700 876 3734 910
rect 3769 876 3803 910
rect 3838 876 3872 910
rect 3907 876 3941 910
rect 3976 876 4010 910
rect 4045 876 4079 910
rect 4114 876 4148 910
rect 4183 842 28085 978
rect 1561 808 1595 842
rect 1630 808 1664 842
rect 1699 808 1733 842
rect 1768 808 1802 842
rect 1837 808 1871 842
rect 1906 808 1940 842
rect 1975 808 2009 842
rect 2044 808 2078 842
rect 2113 808 2147 842
rect 2182 808 2216 842
rect 2251 808 2285 842
rect 2320 808 2354 842
rect 2389 808 2423 842
rect 2458 808 2492 842
rect 2527 808 2561 842
rect 2596 808 2630 842
rect 2665 808 2699 842
rect 2734 808 2768 842
rect 2803 808 2837 842
rect 2872 808 2906 842
rect 2941 808 2975 842
rect 3010 808 3044 842
rect 3079 808 3113 842
rect 3148 808 3182 842
rect 3217 808 3251 842
rect 3286 808 3320 842
rect 3355 808 3389 842
rect 3424 808 3458 842
rect 3493 808 3527 842
rect 3562 808 3596 842
rect 3631 808 3665 842
rect 3700 808 3734 842
rect 3769 808 3803 842
rect 3838 808 3872 842
rect 3907 808 3941 842
rect 3976 808 4010 842
rect 4045 808 4079 842
rect 4114 808 4148 842
rect 4183 808 27881 842
<< locali >>
rect 1357 9246 1480 9280
rect 1514 9246 1548 9280
rect 1357 9232 1548 9246
rect 1347 9226 1548 9232
rect 1347 9212 1425 9226
rect 1347 9154 1357 9212
rect 1459 9192 1498 9226
rect 1532 9192 1548 9226
rect 1459 9178 1548 9192
rect 1459 9154 1616 9178
rect 1347 1992 1353 9154
rect 1459 9144 1498 9154
rect 1532 9120 1571 9154
rect 1605 9120 1616 9154
rect 27966 9194 28095 9280
rect 27966 9160 27983 9194
rect 28017 9160 28055 9194
rect 28089 9160 28095 9194
rect 1527 9110 1616 9120
rect 27966 9114 28095 9160
rect 27966 9110 27983 9114
rect 1527 9082 5585 9110
rect 1531 9048 1570 9082
rect 1604 9048 1643 9082
rect 1677 9048 1716 9082
rect 1750 9048 1789 9082
rect 1823 9048 1862 9082
rect 1896 9048 1935 9082
rect 1969 9048 2008 9082
rect 2042 9048 2081 9082
rect 2115 9048 2154 9082
rect 2188 9048 2227 9082
rect 2261 9048 2300 9082
rect 2334 9048 2373 9082
rect 2407 9048 2446 9082
rect 2480 9048 2519 9082
rect 2553 9048 2592 9082
rect 2626 9048 2665 9082
rect 2699 9048 2738 9082
rect 2772 9048 2811 9082
rect 2845 9048 2884 9082
rect 2918 9048 2957 9082
rect 2991 9048 3030 9082
rect 3064 9048 3103 9082
rect 3137 9048 3176 9082
rect 3210 9048 3249 9082
rect 3283 9048 3322 9082
rect 3356 9048 3395 9082
rect 3429 9048 3468 9082
rect 3502 9048 3541 9082
rect 3575 9048 3614 9082
rect 3648 9048 3687 9082
rect 3721 9048 3760 9082
rect 3794 9048 3833 9082
rect 3867 9048 3906 9082
rect 3940 9048 3979 9082
rect 4013 9048 4052 9082
rect 4086 9048 4125 9082
rect 4159 9048 4198 9082
rect 4232 9048 4271 9082
rect 4305 9048 4344 9082
rect 4378 9048 4417 9082
rect 4451 9048 4490 9082
rect 4524 9048 4563 9082
rect 4597 9048 4636 9082
rect 4670 9048 4709 9082
rect 4743 9048 4782 9082
rect 4816 9048 4855 9082
rect 4889 9048 4928 9082
rect 4962 9048 5001 9082
rect 5035 9048 5074 9082
rect 5108 9048 5147 9082
rect 5181 9048 5220 9082
rect 5254 9048 5293 9082
rect 5327 9048 5366 9082
rect 5400 9048 5439 9082
rect 5473 9048 5512 9082
rect 5546 9048 5585 9082
rect 27867 9080 27911 9110
rect 27945 9080 27983 9110
rect 28017 9080 28055 9114
rect 28089 9080 28095 9114
rect 27867 9048 28095 9080
rect 1531 9042 28095 9048
rect 1531 2064 1537 9042
rect 27905 9036 28095 9042
rect 27905 9034 27915 9036
rect 28085 9034 28095 9036
rect 27905 9000 27911 9034
rect 28089 9000 28095 9034
rect 27905 8954 27915 9000
rect 28085 8954 28095 9000
rect 27905 8920 27911 8954
rect 28089 8920 28095 8954
rect 27905 8875 27915 8920
rect 28085 8875 28095 8920
rect 1527 2025 1537 2064
rect 1347 1953 1357 1992
rect 1531 1991 1537 2025
rect 1347 1919 1353 1953
rect 1527 1952 1537 1991
rect 1347 1880 1357 1919
rect 1531 1918 1537 1952
rect 1347 1846 1353 1880
rect 1527 1879 1537 1918
rect 1347 1807 1357 1846
rect 1531 1845 1537 1879
rect 1347 1773 1353 1807
rect 1527 1806 1537 1845
rect 1347 1734 1357 1773
rect 1531 1772 1537 1806
rect 1347 1700 1353 1734
rect 1527 1733 1537 1772
rect 1347 1661 1357 1700
rect 1531 1699 1537 1733
rect 1347 1627 1353 1661
rect 1527 1660 1537 1699
rect 1347 1588 1357 1627
rect 1531 1626 1537 1660
rect 1347 1554 1353 1588
rect 1527 1587 1537 1626
rect 1347 1515 1357 1554
rect 1531 1553 1537 1587
rect 1347 1481 1353 1515
rect 1527 1514 1537 1553
rect 1347 1442 1357 1481
rect 1531 1480 1537 1514
rect 1347 1408 1353 1442
rect 1527 1441 1537 1480
rect 1347 1369 1357 1408
rect 1531 1407 1537 1441
rect 1347 1335 1353 1369
rect 1527 1368 1537 1407
rect 1347 1296 1357 1335
rect 1531 1334 1537 1368
rect 1347 1262 1353 1296
rect 1527 1295 1537 1334
rect 1347 1223 1357 1262
rect 1531 1261 1537 1295
rect 1795 8847 27692 8853
rect 1795 8775 1873 8847
rect 1907 8843 1946 8847
rect 1980 8843 2019 8847
rect 2053 8843 2092 8847
rect 1795 5357 1801 8775
rect 27614 8775 27692 8847
rect 27686 8741 27692 8775
rect 1907 8703 1941 8741
rect 27542 8707 27580 8741
rect 1979 8669 2018 8673
rect 2052 8669 2091 8673
rect 2125 8669 2164 8673
rect 27682 8701 27692 8741
rect 1979 8663 27512 8669
rect 27686 8667 27692 8701
rect 1979 5429 1985 8663
rect 27502 8629 27512 8663
rect 27502 8595 27508 8629
rect 27682 8627 27692 8667
rect 27502 8555 27512 8595
rect 27686 8593 27692 8627
rect 27502 8521 27508 8555
rect 27682 8553 27692 8593
rect 27502 8481 27512 8521
rect 27686 8519 27692 8553
rect 1907 5390 1985 5429
rect 1907 5369 1945 5390
rect 1795 5335 1805 5357
rect 1839 5335 1873 5357
rect 1907 5335 1941 5369
rect 1979 5356 1985 5390
rect 1975 5335 1985 5356
rect 1795 5318 1985 5335
rect 1795 5284 1801 5318
rect 1835 5300 1873 5318
rect 1907 5317 1985 5318
rect 1907 5300 1945 5317
rect 1795 5266 1805 5284
rect 1839 5266 1873 5300
rect 1907 5266 1941 5300
rect 1979 5283 1985 5317
rect 1975 5266 1985 5283
rect 1795 5245 1985 5266
rect 1795 5211 1801 5245
rect 1835 5231 1873 5245
rect 1907 5244 1985 5245
rect 1907 5231 1945 5244
rect 1795 5197 1805 5211
rect 1839 5197 1873 5231
rect 1907 5197 1941 5231
rect 1979 5210 1985 5244
rect 1975 5197 1985 5210
rect 1795 5172 1985 5197
rect 1795 5138 1801 5172
rect 1835 5162 1873 5172
rect 1907 5171 1985 5172
rect 1907 5162 1945 5171
rect 1795 5128 1805 5138
rect 1839 5128 1873 5162
rect 1907 5128 1941 5162
rect 1979 5137 1985 5171
rect 1975 5128 1985 5137
rect 1795 5099 1985 5128
rect 1795 5065 1801 5099
rect 1835 5093 1873 5099
rect 1907 5098 1985 5099
rect 1907 5093 1945 5098
rect 1795 5059 1805 5065
rect 1839 5059 1873 5093
rect 1907 5059 1941 5093
rect 1979 5064 1985 5098
rect 1975 5059 1985 5064
rect 1795 5026 1985 5059
rect 1795 4992 1801 5026
rect 1835 5024 1873 5026
rect 1907 5025 1985 5026
rect 1907 5024 1945 5025
rect 1795 4990 1805 4992
rect 1839 4990 1873 5024
rect 1907 4990 1941 5024
rect 1979 4991 1985 5025
rect 1975 4990 1985 4991
rect 1795 4955 1985 4990
rect 1795 4953 1805 4955
rect 1795 4919 1801 4953
rect 1839 4921 1873 4955
rect 1907 4921 1941 4955
rect 1975 4952 1985 4955
rect 1835 4919 1873 4921
rect 1907 4919 1945 4921
rect 1795 4918 1945 4919
rect 1979 4918 1985 4952
rect 1795 4886 1985 4918
rect 1795 4880 1805 4886
rect 1795 4846 1801 4880
rect 1839 4852 1873 4886
rect 1907 4852 1941 4886
rect 1975 4879 1985 4886
rect 1835 4846 1873 4852
rect 1907 4846 1945 4852
rect 1795 4845 1945 4846
rect 1979 4845 1985 4879
rect 1795 4817 1985 4845
rect 1795 4807 1805 4817
rect 1795 4773 1801 4807
rect 1839 4783 1873 4817
rect 1907 4783 1941 4817
rect 1975 4806 1985 4817
rect 1835 4773 1873 4783
rect 1907 4773 1945 4783
rect 1795 4772 1945 4773
rect 1979 4772 1985 4806
rect 1795 4748 1985 4772
rect 1795 4734 1805 4748
rect 1795 4700 1801 4734
rect 1839 4714 1873 4748
rect 1907 4714 1941 4748
rect 1975 4733 1985 4748
rect 1835 4700 1873 4714
rect 1907 4700 1945 4714
rect 1795 4699 1945 4700
rect 1979 4699 1985 4733
rect 1795 4679 1985 4699
rect 1795 4661 1805 4679
rect 1795 4627 1801 4661
rect 1839 4645 1873 4679
rect 1907 4645 1941 4679
rect 1975 4660 1985 4679
rect 1835 4627 1873 4645
rect 1907 4627 1945 4645
rect 1795 4626 1945 4627
rect 1979 4626 1985 4660
rect 1795 4610 1985 4626
rect 1795 4588 1805 4610
rect 1795 4554 1801 4588
rect 1839 4576 1873 4610
rect 1907 4576 1941 4610
rect 1975 4587 1985 4610
rect 1835 4554 1873 4576
rect 1907 4554 1945 4576
rect 1795 4553 1945 4554
rect 1979 4553 1985 4587
rect 1795 4541 1985 4553
rect 1795 4515 1805 4541
rect 1795 4481 1801 4515
rect 1839 4507 1873 4541
rect 1907 4507 1941 4541
rect 1975 4514 1985 4541
rect 1835 4481 1873 4507
rect 1907 4481 1945 4507
rect 1795 4480 1945 4481
rect 1979 4480 1985 4514
rect 1795 4472 1985 4480
rect 1795 4442 1805 4472
rect 1795 4408 1801 4442
rect 1839 4438 1873 4472
rect 1907 4438 1941 4472
rect 1975 4441 1985 4472
rect 1835 4408 1873 4438
rect 1907 4408 1945 4438
rect 1795 4407 1945 4408
rect 1979 4407 1985 4441
rect 1795 4403 1985 4407
rect 1795 4369 1805 4403
rect 1839 4369 1873 4403
rect 1907 4369 1941 4403
rect 1975 4369 1985 4403
rect 1795 4335 1801 4369
rect 1835 4335 1873 4369
rect 1907 4368 1985 4369
rect 1907 4335 1945 4368
rect 1795 4334 1945 4335
rect 1979 4334 1985 4368
rect 1795 4300 1805 4334
rect 1839 4300 1873 4334
rect 1907 4300 1941 4334
rect 1975 4300 1985 4334
rect 1795 4296 1985 4300
rect 1795 4262 1801 4296
rect 1835 4265 1873 4296
rect 1907 4295 1985 4296
rect 1907 4265 1945 4295
rect 1795 4231 1805 4262
rect 1839 4231 1873 4265
rect 1907 4231 1941 4265
rect 1979 4261 1985 4295
rect 1975 4231 1985 4261
rect 1795 4223 1985 4231
rect 1795 4189 1801 4223
rect 1835 4196 1873 4223
rect 1907 4222 1985 4223
rect 1907 4196 1945 4222
rect 1795 4162 1805 4189
rect 1839 4162 1873 4196
rect 1907 4162 1941 4196
rect 1979 4188 1985 4222
rect 1975 4162 1985 4188
rect 1795 4150 1985 4162
rect 1795 4116 1801 4150
rect 1835 4127 1873 4150
rect 1907 4149 1985 4150
rect 1907 4127 1945 4149
rect 1795 4093 1805 4116
rect 1839 4093 1873 4127
rect 1907 4093 1941 4127
rect 1979 4115 1985 4149
rect 1975 4093 1985 4115
rect 1795 4077 1985 4093
rect 1795 4043 1801 4077
rect 1835 4058 1873 4077
rect 1907 4076 1985 4077
rect 1907 4058 1945 4076
rect 1795 4024 1805 4043
rect 1839 4024 1873 4058
rect 1907 4024 1941 4058
rect 1979 4042 1985 4076
rect 1975 4024 1985 4042
rect 1795 4004 1985 4024
rect 1795 3970 1801 4004
rect 1835 3989 1873 4004
rect 1907 4003 1985 4004
rect 1907 3989 1945 4003
rect 1795 3955 1805 3970
rect 1839 3955 1873 3989
rect 1907 3955 1941 3989
rect 1979 3969 1985 4003
rect 1975 3955 1985 3969
rect 1795 3931 1985 3955
rect 1795 3897 1801 3931
rect 1835 3920 1873 3931
rect 1907 3930 1985 3931
rect 1907 3920 1945 3930
rect 1795 3858 1805 3897
rect 1979 3896 1985 3930
rect 1795 3824 1801 3858
rect 1975 3857 1985 3896
rect 1795 3785 1805 3824
rect 1979 3823 1985 3857
rect 1795 3751 1801 3785
rect 1975 3784 1985 3823
rect 1795 3712 1805 3751
rect 1979 3750 1985 3784
rect 1795 3678 1801 3712
rect 1975 3711 1985 3750
rect 1795 3639 1805 3678
rect 1979 3677 1985 3711
rect 1795 3605 1801 3639
rect 1975 3638 1985 3677
rect 1795 3566 1805 3605
rect 1979 3604 1985 3638
rect 1795 3532 1801 3566
rect 1975 3565 1985 3604
rect 1795 3493 1805 3532
rect 1979 3531 1985 3565
rect 1795 3459 1801 3493
rect 1975 3492 1985 3531
rect 1795 3420 1805 3459
rect 1979 3458 1985 3492
rect 1795 3386 1801 3420
rect 1975 3419 1985 3458
rect 1795 3347 1805 3386
rect 1979 3385 1985 3419
rect 1795 3313 1801 3347
rect 1975 3346 1985 3385
rect 1795 3274 1805 3313
rect 1979 3312 1985 3346
rect 1795 3240 1801 3274
rect 1975 3273 1985 3312
rect 1795 3201 1805 3240
rect 1979 3239 1985 3273
rect 1795 3167 1801 3201
rect 1975 3200 1985 3239
rect 1795 3128 1805 3167
rect 1979 3166 1985 3200
rect 1795 3094 1801 3128
rect 1975 3127 1985 3166
rect 1795 3055 1805 3094
rect 1979 3093 1985 3127
rect 1795 3021 1801 3055
rect 1975 3054 1985 3093
rect 1795 2982 1805 3021
rect 1979 3020 1985 3054
rect 1795 2948 1801 2982
rect 1975 2981 1985 3020
rect 1795 2909 1805 2948
rect 1979 2947 1985 2981
rect 1795 2875 1801 2909
rect 1975 2908 1985 2947
rect 1795 2836 1805 2875
rect 1979 2874 1985 2908
rect 1795 2802 1801 2836
rect 1975 2835 1985 2874
rect 1795 2763 1805 2802
rect 1979 2801 1985 2835
rect 1795 2729 1801 2763
rect 1975 2762 1985 2801
rect 1795 2690 1805 2729
rect 1979 2728 1985 2762
rect 1795 2656 1801 2690
rect 1975 2689 1985 2728
rect 1795 2617 1805 2656
rect 1979 2655 1985 2689
rect 1795 2583 1801 2617
rect 1975 2616 1985 2655
rect 1795 2544 1805 2583
rect 1979 2582 1985 2616
rect 1795 2510 1801 2544
rect 1975 2543 1985 2582
rect 1795 2471 1805 2510
rect 1979 2509 1985 2543
rect 1795 2437 1801 2471
rect 1975 2470 1985 2509
rect 1795 2398 1805 2437
rect 1979 2436 1985 2470
rect 1795 2364 1801 2398
rect 1975 2397 1985 2436
rect 1795 2325 1805 2364
rect 1979 2363 1985 2397
rect 1795 2291 1801 2325
rect 1975 2324 1985 2363
rect 1795 2252 1805 2291
rect 1979 2290 1985 2324
rect 1795 2218 1801 2252
rect 1975 2251 1985 2290
rect 2181 8461 27294 8467
rect 2181 8427 2259 8461
rect 2293 8458 2332 8461
rect 2366 8458 2405 8461
rect 2439 8458 2478 8461
rect 2512 8458 2551 8461
rect 2585 8458 2624 8461
rect 2658 8458 2697 8461
rect 2731 8458 2770 8461
rect 2804 8458 2843 8461
rect 2877 8458 2916 8461
rect 2950 8458 2989 8461
rect 3023 8458 3062 8461
rect 2307 8427 2332 8458
rect 2181 8424 2273 8427
rect 2307 8424 2341 8427
rect 2181 8390 2341 8424
rect 2181 8389 2191 8390
rect 2293 8389 2341 8390
rect 2181 5259 2187 8389
rect 2293 8355 2332 8389
rect 2366 8355 2405 8356
rect 27216 8389 27294 8461
rect 27216 8357 27254 8389
rect 27216 8355 27229 8357
rect 27288 8355 27294 8389
rect 2293 8322 2409 8355
rect 2361 8317 2409 8322
rect 2365 8283 2404 8317
rect 27144 8323 27229 8355
rect 27263 8323 27294 8355
rect 27144 8315 27294 8323
rect 27144 8289 27182 8315
rect 27216 8289 27254 8315
rect 2438 8283 2477 8288
rect 2511 8283 2550 8288
rect 2584 8283 2623 8288
rect 2657 8283 2696 8288
rect 2730 8283 2769 8288
rect 2803 8283 2842 8288
rect 2876 8283 2915 8288
rect 2949 8283 2988 8288
rect 3022 8283 3061 8288
rect 3095 8283 3134 8288
rect 27144 8283 27161 8289
rect 2365 8277 27161 8283
rect 27288 8281 27294 8315
rect 2365 5331 2371 8277
rect 2361 5292 2371 5331
rect 2181 5220 2191 5259
rect 2365 5258 2371 5292
rect 2181 5186 2187 5220
rect 2361 5219 2371 5258
rect 2181 5147 2191 5186
rect 2365 5185 2371 5219
rect 2181 5113 2187 5147
rect 2361 5146 2371 5185
rect 2181 5074 2191 5113
rect 2365 5112 2371 5146
rect 2181 5040 2187 5074
rect 2361 5073 2371 5112
rect 2181 5001 2191 5040
rect 2365 5039 2371 5073
rect 2181 4967 2187 5001
rect 2361 5000 2371 5039
rect 2181 4928 2191 4967
rect 2365 4966 2371 5000
rect 2181 4894 2187 4928
rect 2361 4927 2371 4966
rect 2181 4855 2191 4894
rect 2365 4893 2371 4927
rect 2181 4821 2187 4855
rect 2361 4854 2371 4893
rect 2181 4782 2191 4821
rect 2365 4820 2371 4854
rect 2181 4748 2187 4782
rect 2361 4781 2371 4820
rect 2181 4709 2191 4748
rect 2365 4747 2371 4781
rect 2181 4675 2187 4709
rect 2361 4708 2371 4747
rect 2181 4636 2191 4675
rect 2365 4674 2371 4708
rect 2181 4602 2187 4636
rect 2361 4635 2371 4674
rect 2181 4563 2191 4602
rect 2365 4601 2371 4635
rect 2181 4529 2187 4563
rect 2361 4562 2371 4601
rect 2181 4490 2191 4529
rect 2365 4528 2371 4562
rect 2181 4456 2187 4490
rect 2361 4489 2371 4528
rect 2181 4417 2191 4456
rect 2365 4455 2371 4489
rect 2181 4383 2187 4417
rect 2361 4416 2371 4455
rect 2181 4344 2191 4383
rect 2365 4382 2371 4416
rect 2181 4310 2187 4344
rect 2361 4343 2371 4382
rect 2181 4271 2191 4310
rect 2365 4309 2371 4343
rect 2181 4237 2187 4271
rect 2361 4270 2371 4309
rect 2181 4198 2191 4237
rect 2365 4236 2371 4270
rect 2181 4164 2187 4198
rect 2361 4197 2371 4236
rect 2181 4125 2191 4164
rect 2365 4163 2371 4197
rect 2181 4091 2187 4125
rect 2361 4124 2371 4163
rect 2181 4052 2191 4091
rect 2365 4090 2371 4124
rect 2181 4018 2187 4052
rect 2361 4051 2371 4090
rect 2181 3979 2191 4018
rect 2365 4017 2371 4051
rect 2181 3945 2187 3979
rect 2361 3978 2371 4017
rect 2181 3906 2191 3945
rect 2365 3944 2371 3978
rect 2181 3872 2187 3906
rect 2361 3905 2371 3944
rect 2181 3833 2191 3872
rect 2365 3871 2371 3905
rect 2181 3799 2187 3833
rect 2361 3832 2371 3871
rect 2181 3760 2191 3799
rect 2365 3798 2371 3832
rect 2181 3726 2187 3760
rect 2361 3759 2371 3798
rect 2181 3687 2191 3726
rect 2365 3725 2371 3759
rect 2181 3653 2187 3687
rect 2361 3686 2371 3725
rect 2181 3614 2191 3653
rect 2365 3652 2371 3686
rect 2181 3580 2187 3614
rect 2361 3613 2371 3652
rect 2181 3541 2191 3580
rect 2365 3579 2371 3613
rect 2181 3507 2187 3541
rect 2361 3540 2371 3579
rect 2181 3468 2191 3507
rect 2365 3506 2371 3540
rect 2181 3434 2187 3468
rect 2361 3467 2371 3506
rect 2181 3395 2191 3434
rect 2365 3433 2371 3467
rect 2181 3361 2187 3395
rect 2361 3394 2371 3433
rect 2181 3322 2191 3361
rect 2365 3360 2371 3394
rect 2181 3288 2187 3322
rect 2361 3321 2371 3360
rect 2181 3249 2191 3288
rect 2365 3287 2371 3321
rect 2181 3215 2187 3249
rect 2361 3248 2371 3287
rect 2181 3176 2191 3215
rect 2365 3214 2371 3248
rect 2181 3142 2187 3176
rect 2361 3175 2371 3214
rect 2181 3103 2191 3142
rect 2365 3141 2371 3175
rect 2181 3069 2187 3103
rect 2361 3102 2371 3141
rect 2181 3030 2191 3069
rect 2365 3068 2371 3102
rect 2181 2996 2187 3030
rect 2361 3029 2371 3068
rect 2181 2957 2191 2996
rect 2365 2995 2371 3029
rect 2181 2923 2187 2957
rect 2361 2956 2371 2995
rect 2181 2916 2191 2923
rect 2365 2922 2371 2956
rect 2361 2916 2371 2922
rect 2181 2884 2371 2916
rect 2181 2850 2187 2884
rect 2221 2850 2259 2884
rect 2293 2883 2371 2884
rect 2293 2850 2331 2883
rect 2181 2849 2331 2850
rect 2365 2849 2371 2883
rect 2181 2811 2371 2849
rect 2181 2777 2187 2811
rect 2221 2790 2259 2811
rect 2293 2810 2371 2811
rect 2293 2790 2331 2810
rect 2181 2738 2191 2777
rect 2365 2776 2371 2810
rect 2181 2704 2187 2738
rect 2361 2737 2371 2776
rect 2181 2665 2191 2704
rect 2365 2703 2371 2737
rect 2181 2631 2187 2665
rect 2361 2664 2371 2703
rect 2181 2592 2191 2631
rect 2365 2630 2371 2664
rect 2181 2558 2187 2592
rect 2361 2591 2371 2630
rect 2181 2519 2191 2558
rect 2365 2557 2371 2591
rect 2181 2485 2187 2519
rect 2361 2518 2371 2557
rect 2181 2446 2191 2485
rect 2365 2484 2371 2518
rect 2293 2451 2371 2484
rect 27093 8243 27161 8277
rect 27093 8221 27110 8243
rect 27144 8221 27161 8243
rect 27263 8241 27294 8281
rect 27288 8207 27294 8241
rect 27263 8167 27294 8207
rect 27288 8133 27294 8167
rect 27263 8093 27294 8133
rect 27288 8059 27294 8093
rect 27263 8019 27294 8059
rect 27288 7985 27294 8019
rect 27263 7946 27294 7985
rect 27288 7912 27294 7946
rect 27263 7873 27294 7912
rect 27288 7839 27294 7873
rect 27263 7763 27294 7839
rect 27288 7729 27294 7763
rect 27263 7690 27294 7729
rect 27288 7656 27294 7690
rect 27263 7617 27294 7656
rect 27288 7583 27294 7617
rect 27263 7544 27294 7583
rect 27288 7510 27294 7544
rect 27263 7471 27294 7510
rect 27288 7437 27294 7471
rect 27263 7398 27294 7437
rect 27288 7364 27294 7398
rect 27263 7325 27294 7364
rect 27288 7291 27294 7325
rect 27263 7252 27294 7291
rect 27288 7218 27294 7252
rect 27263 7179 27294 7218
rect 27288 7145 27294 7179
rect 27263 7106 27294 7145
rect 27288 7072 27294 7106
rect 27263 7033 27294 7072
rect 27288 6999 27294 7033
rect 27263 6960 27294 6999
rect 27288 6926 27294 6960
rect 27263 6887 27294 6926
rect 27288 6853 27294 6887
rect 27263 6814 27294 6853
rect 27288 6780 27294 6814
rect 27263 6741 27294 6780
rect 27288 6707 27294 6741
rect 27263 6668 27294 6707
rect 27288 6634 27294 6668
rect 27263 6595 27294 6634
rect 27288 6561 27294 6595
rect 27263 6522 27294 6561
rect 27288 6488 27294 6522
rect 27263 6449 27294 6488
rect 27288 6415 27294 6449
rect 27263 6376 27294 6415
rect 27288 6342 27294 6376
rect 27263 6303 27294 6342
rect 27288 6269 27294 6303
rect 27263 6230 27294 6269
rect 27288 6196 27294 6230
rect 27263 6157 27294 6196
rect 27288 6123 27294 6157
rect 27263 6084 27294 6123
rect 27288 6050 27294 6084
rect 27263 6011 27294 6050
rect 27288 5977 27294 6011
rect 27263 5938 27294 5977
rect 27288 5904 27294 5938
rect 27263 5865 27294 5904
rect 27288 5831 27294 5865
rect 27263 5792 27294 5831
rect 27288 5758 27294 5792
rect 27263 5719 27294 5758
rect 27288 5685 27294 5719
rect 27263 5646 27294 5685
rect 27288 5612 27294 5646
rect 27263 5573 27294 5612
rect 27288 5539 27294 5573
rect 27263 5500 27294 5539
rect 27288 5466 27294 5500
rect 27263 5427 27294 5466
rect 27288 5393 27294 5427
rect 27263 5354 27294 5393
rect 27288 5320 27294 5354
rect 27263 5281 27294 5320
rect 27288 5247 27294 5281
rect 27263 5208 27294 5247
rect 27288 5174 27294 5208
rect 27263 5135 27294 5174
rect 27288 5101 27294 5135
rect 27263 5062 27294 5101
rect 27288 5028 27294 5062
rect 27263 4989 27294 5028
rect 27288 4955 27294 4989
rect 27263 4916 27294 4955
rect 27288 4882 27294 4916
rect 27263 4843 27294 4882
rect 27288 4809 27294 4843
rect 27263 4770 27294 4809
rect 27288 4736 27294 4770
rect 27263 4697 27294 4736
rect 27288 4663 27294 4697
rect 27263 4624 27294 4663
rect 27288 4590 27294 4624
rect 27263 4551 27294 4590
rect 27288 4517 27294 4551
rect 27263 4478 27294 4517
rect 27288 4444 27294 4478
rect 27263 4405 27294 4444
rect 27288 4371 27294 4405
rect 27263 4332 27294 4371
rect 27288 4298 27294 4332
rect 27263 4259 27294 4298
rect 27288 4225 27294 4259
rect 27263 4186 27294 4225
rect 27288 4152 27294 4186
rect 27263 4113 27294 4152
rect 27288 4079 27294 4113
rect 27263 4040 27294 4079
rect 27288 4006 27294 4040
rect 27263 3967 27294 4006
rect 27288 3933 27294 3967
rect 27263 3894 27294 3933
rect 27288 3860 27294 3894
rect 27263 3821 27294 3860
rect 27288 3787 27294 3821
rect 27263 3748 27294 3787
rect 27288 3714 27294 3748
rect 27263 3675 27294 3714
rect 27288 3641 27294 3675
rect 27263 3602 27294 3641
rect 27288 3568 27294 3602
rect 27263 3529 27294 3568
rect 27288 3495 27294 3529
rect 27263 3456 27294 3495
rect 27288 3422 27294 3456
rect 27263 3383 27294 3422
rect 27288 3349 27294 3383
rect 27263 3310 27294 3349
rect 27288 3276 27294 3310
rect 27263 3237 27294 3276
rect 2181 2412 2187 2446
rect 2293 2445 27093 2451
rect 2293 2441 2331 2445
rect 26341 2441 26380 2445
rect 26414 2441 26453 2445
rect 26487 2441 26526 2445
rect 26560 2441 26599 2445
rect 26633 2441 26672 2445
rect 26706 2441 26745 2445
rect 26779 2441 26818 2445
rect 26852 2441 26891 2445
rect 26925 2441 26964 2445
rect 26998 2441 27037 2445
rect 2221 2412 2259 2416
rect 2293 2412 2327 2441
rect 2181 2382 2327 2412
rect 2181 2373 2191 2382
rect 2225 2373 2327 2382
rect 27071 2411 27093 2445
rect 27045 2407 27093 2411
rect 27045 2373 27161 2407
rect 2181 2339 2187 2373
rect 2225 2348 2259 2373
rect 2221 2339 2259 2348
rect 2181 2267 2259 2339
rect 27143 2339 27161 2373
rect 27288 2339 27294 3237
rect 27113 2305 27294 2339
rect 27113 2301 27147 2305
rect 27143 2271 27147 2301
rect 27181 2301 27294 2305
rect 27181 2271 27182 2301
rect 26413 2267 26452 2271
rect 26486 2267 26525 2271
rect 26559 2267 26598 2271
rect 26632 2267 26671 2271
rect 26705 2267 26744 2271
rect 26778 2267 26817 2271
rect 26851 2267 26890 2271
rect 26924 2267 26963 2271
rect 26997 2267 27036 2271
rect 27070 2267 27109 2271
rect 27143 2267 27182 2271
rect 27216 2267 27294 2301
rect 2181 2261 27294 2267
rect 27502 8447 27508 8481
rect 27682 8479 27692 8519
rect 27502 8407 27512 8447
rect 27686 8445 27692 8479
rect 27502 8373 27508 8407
rect 27682 8405 27692 8445
rect 27502 8333 27512 8373
rect 27686 8371 27692 8405
rect 27502 8299 27508 8333
rect 27682 8332 27692 8371
rect 27502 8259 27512 8299
rect 27686 8298 27692 8332
rect 27682 8259 27692 8298
rect 27502 8225 27508 8259
rect 27686 8225 27692 8259
rect 27502 8149 27512 8225
rect 27682 8149 27692 8225
rect 27502 8115 27508 8149
rect 27686 8115 27692 8149
rect 27502 8076 27512 8115
rect 27682 8076 27692 8115
rect 27502 8042 27508 8076
rect 27686 8042 27692 8076
rect 27502 8003 27512 8042
rect 27682 8003 27692 8042
rect 27502 7969 27508 8003
rect 27686 7969 27692 8003
rect 27502 7930 27512 7969
rect 27682 7930 27692 7969
rect 27502 7896 27508 7930
rect 27686 7896 27692 7930
rect 27502 7857 27512 7896
rect 27682 7857 27692 7896
rect 27502 7823 27508 7857
rect 27686 7823 27692 7857
rect 27502 7784 27512 7823
rect 27682 7784 27692 7823
rect 1795 2179 1805 2218
rect 1979 2217 1985 2251
rect 1795 2145 1801 2179
rect 1975 2178 1985 2217
rect 1795 2106 1805 2145
rect 1979 2144 1985 2178
rect 1795 2072 1801 2106
rect 1975 2105 1985 2144
rect 1795 2033 1805 2072
rect 1979 2071 1985 2105
rect 1795 1999 1801 2033
rect 1975 2032 1985 2071
rect 1795 1960 1805 1999
rect 1979 1998 1985 2032
rect 1975 1996 1985 1998
rect 27502 1996 27508 7784
rect 1975 1995 27508 1996
rect 1975 1961 2009 1995
rect 2043 1961 2078 1995
rect 2112 1961 2147 1995
rect 2181 1961 2216 1995
rect 2250 1961 2284 1995
rect 2318 1961 2352 1995
rect 2386 1961 2420 1995
rect 2454 1961 2488 1995
rect 2522 1961 2556 1995
rect 2590 1961 2624 1995
rect 2658 1961 2692 1995
rect 2726 1961 2760 1995
rect 2794 1961 2828 1995
rect 2862 1961 2896 1995
rect 2930 1961 2964 1995
rect 2998 1961 3032 1995
rect 3066 1961 3100 1995
rect 3134 1961 3168 1995
rect 3202 1961 3236 1995
rect 3270 1961 3304 1995
rect 3338 1961 3372 1995
rect 3406 1961 3440 1995
rect 3474 1961 3508 1995
rect 3542 1961 3576 1995
rect 3610 1961 3644 1995
rect 3678 1961 3712 1995
rect 3746 1961 3780 1995
rect 3814 1961 3848 1995
rect 3882 1961 3916 1995
rect 3950 1961 3984 1995
rect 4018 1961 4052 1995
rect 4086 1961 4120 1995
rect 4154 1961 4188 1995
rect 4222 1961 4256 1995
rect 4290 1961 4324 1995
rect 4358 1961 4392 1995
rect 4426 1961 4460 1995
rect 4494 1961 4528 1995
rect 4562 1961 4596 1995
rect 4630 1961 4664 1995
rect 4698 1961 4732 1995
rect 4766 1961 4800 1995
rect 4834 1961 4868 1995
rect 4902 1961 4936 1995
rect 4970 1961 5004 1995
rect 5038 1961 5072 1995
rect 5106 1961 5140 1995
rect 5174 1961 5208 1995
rect 5242 1961 5276 1995
rect 5310 1961 5344 1995
rect 5378 1961 5412 1995
rect 5446 1961 5480 1995
rect 5514 1961 5548 1995
rect 5582 1961 5616 1995
rect 5650 1961 5684 1995
rect 5718 1961 5752 1995
rect 5786 1961 5820 1995
rect 5854 1961 5888 1995
rect 5922 1961 5956 1995
rect 5990 1961 6024 1995
rect 6058 1961 6092 1995
rect 6126 1961 6160 1995
rect 6194 1961 6228 1995
rect 6262 1961 6296 1995
rect 6330 1961 6364 1995
rect 6398 1961 6432 1995
rect 6466 1961 6500 1995
rect 6534 1961 6568 1995
rect 6602 1961 6636 1995
rect 6670 1961 6704 1995
rect 6738 1961 6772 1995
rect 6806 1961 6840 1995
rect 6874 1961 6908 1995
rect 6942 1961 6976 1995
rect 7010 1961 7044 1995
rect 7078 1961 7112 1995
rect 7146 1961 7180 1995
rect 7214 1961 7248 1995
rect 7282 1961 7316 1995
rect 7350 1961 7384 1995
rect 7418 1961 7452 1995
rect 7486 1961 7520 1995
rect 7554 1961 7588 1995
rect 7622 1961 7656 1995
rect 7690 1961 7724 1995
rect 7758 1961 7792 1995
rect 7826 1961 7860 1995
rect 7894 1961 7928 1995
rect 7962 1961 7996 1995
rect 8030 1961 8064 1995
rect 8098 1961 8132 1995
rect 8166 1961 8200 1995
rect 8234 1961 8268 1995
rect 8302 1961 8336 1995
rect 8370 1961 8404 1995
rect 8438 1961 8472 1995
rect 8506 1961 8540 1995
rect 8574 1961 8608 1995
rect 8642 1961 8676 1995
rect 8710 1961 8744 1995
rect 8778 1961 8812 1995
rect 8846 1961 8880 1995
rect 8914 1961 8948 1995
rect 8982 1961 9016 1995
rect 9050 1961 9084 1995
rect 9118 1961 9152 1995
rect 9186 1961 9220 1995
rect 9254 1961 9288 1995
rect 9322 1961 9356 1995
rect 9390 1961 9424 1995
rect 9458 1961 9492 1995
rect 9526 1961 9560 1995
rect 9594 1961 9628 1995
rect 9662 1961 9696 1995
rect 9730 1961 9764 1995
rect 9798 1961 9832 1995
rect 9866 1961 9900 1995
rect 9934 1961 9968 1995
rect 10002 1961 10036 1995
rect 10070 1961 10104 1995
rect 10138 1961 10172 1995
rect 10206 1961 10240 1995
rect 10274 1961 10308 1995
rect 10342 1961 10376 1995
rect 10410 1961 10444 1995
rect 10478 1961 10512 1995
rect 10546 1961 10580 1995
rect 10614 1961 10648 1995
rect 10682 1961 10716 1995
rect 10750 1961 10784 1995
rect 10818 1961 10852 1995
rect 10886 1961 10920 1995
rect 10954 1961 10988 1995
rect 11022 1961 11056 1995
rect 11090 1961 11124 1995
rect 11158 1961 11192 1995
rect 11226 1961 11260 1995
rect 11294 1961 11328 1995
rect 11362 1961 11396 1995
rect 11430 1961 11464 1995
rect 11498 1961 11532 1995
rect 11566 1961 11600 1995
rect 11634 1961 11668 1995
rect 11702 1961 11736 1995
rect 11770 1961 11804 1995
rect 11838 1961 11872 1995
rect 11906 1961 11940 1995
rect 11974 1961 12008 1995
rect 12042 1961 12076 1995
rect 12110 1961 12144 1995
rect 12178 1961 12212 1995
rect 12246 1961 12280 1995
rect 12314 1961 12348 1995
rect 12382 1961 12416 1995
rect 12450 1961 12484 1995
rect 12518 1961 12552 1995
rect 12586 1961 12620 1995
rect 12654 1961 12688 1995
rect 12722 1961 12756 1995
rect 12790 1961 12824 1995
rect 12858 1961 12892 1995
rect 12926 1961 12960 1995
rect 12994 1961 13028 1995
rect 13062 1961 13096 1995
rect 13130 1961 13164 1995
rect 13198 1961 13232 1995
rect 13266 1961 13300 1995
rect 13334 1961 13368 1995
rect 13402 1961 13436 1995
rect 13470 1961 13504 1995
rect 13538 1961 13572 1995
rect 13606 1961 13640 1995
rect 13674 1961 13708 1995
rect 13742 1961 13776 1995
rect 13810 1961 13844 1995
rect 13878 1961 13912 1995
rect 13946 1961 13980 1995
rect 14014 1961 14048 1995
rect 14082 1961 14116 1995
rect 14150 1961 14184 1995
rect 14218 1961 14252 1995
rect 14286 1961 14320 1995
rect 14354 1961 14388 1995
rect 14422 1961 14456 1995
rect 14490 1961 14524 1995
rect 14558 1961 14592 1995
rect 14626 1961 14660 1995
rect 14694 1961 14728 1995
rect 14762 1961 14796 1995
rect 14830 1961 14864 1995
rect 14898 1961 14932 1995
rect 14966 1961 15000 1995
rect 15034 1961 15068 1995
rect 15102 1961 15136 1995
rect 15170 1961 15204 1995
rect 15238 1961 15272 1995
rect 15306 1961 15340 1995
rect 15374 1961 15408 1995
rect 15442 1961 15476 1995
rect 15510 1961 15544 1995
rect 15578 1961 15612 1995
rect 15646 1961 15680 1995
rect 15714 1961 15748 1995
rect 15782 1961 15816 1995
rect 15850 1961 15884 1995
rect 15918 1961 15952 1995
rect 15986 1961 16020 1995
rect 16054 1961 16088 1995
rect 16122 1961 16156 1995
rect 16190 1961 16224 1995
rect 16258 1961 16292 1995
rect 16326 1961 16360 1995
rect 16394 1961 16428 1995
rect 16462 1961 16496 1995
rect 16530 1961 16564 1995
rect 16598 1961 16632 1995
rect 16666 1961 16700 1995
rect 16734 1961 16768 1995
rect 16802 1961 16836 1995
rect 16870 1961 16904 1995
rect 16938 1961 16972 1995
rect 17006 1961 17040 1995
rect 17074 1961 17108 1995
rect 17142 1961 17176 1995
rect 17210 1961 17244 1995
rect 17278 1961 17312 1995
rect 17346 1961 17380 1995
rect 17414 1961 17448 1995
rect 17482 1961 17516 1995
rect 17550 1961 17584 1995
rect 17618 1961 17652 1995
rect 17686 1961 17720 1995
rect 17754 1961 17788 1995
rect 17822 1961 17856 1995
rect 17890 1961 17924 1995
rect 17958 1961 17992 1995
rect 18026 1961 18060 1995
rect 18094 1961 18128 1995
rect 18162 1961 18196 1995
rect 18230 1961 18264 1995
rect 18298 1961 18332 1995
rect 18366 1961 18400 1995
rect 18434 1961 18468 1995
rect 18502 1961 18536 1995
rect 18570 1961 18604 1995
rect 18638 1961 18672 1995
rect 18706 1961 18740 1995
rect 18774 1961 18808 1995
rect 18842 1961 18876 1995
rect 18910 1961 18944 1995
rect 18978 1961 19012 1995
rect 19046 1961 19080 1995
rect 19114 1961 19148 1995
rect 19182 1961 19216 1995
rect 19250 1961 19284 1995
rect 19318 1961 19352 1995
rect 19386 1961 19420 1995
rect 19454 1961 19488 1995
rect 19522 1961 19556 1995
rect 19590 1961 19624 1995
rect 19658 1961 19692 1995
rect 19726 1961 19760 1995
rect 19794 1961 19828 1995
rect 19862 1961 19896 1995
rect 19930 1961 19964 1995
rect 19998 1961 20032 1995
rect 20066 1961 20100 1995
rect 20134 1961 20168 1995
rect 20202 1961 20236 1995
rect 20270 1961 20304 1995
rect 20338 1961 20372 1995
rect 20406 1961 20440 1995
rect 20474 1961 20508 1995
rect 20542 1961 20576 1995
rect 20610 1961 20644 1995
rect 20678 1961 20712 1995
rect 20746 1961 20780 1995
rect 20814 1961 20848 1995
rect 20882 1961 20916 1995
rect 20950 1961 20984 1995
rect 21018 1961 21052 1995
rect 21086 1961 21120 1995
rect 21154 1961 21188 1995
rect 21222 1961 21256 1995
rect 21290 1961 21324 1995
rect 21358 1961 21392 1995
rect 21426 1961 21460 1995
rect 21494 1961 21528 1995
rect 21562 1961 21596 1995
rect 21630 1961 21664 1995
rect 21698 1961 21732 1995
rect 21766 1961 21800 1995
rect 21834 1961 21868 1995
rect 21902 1961 21936 1995
rect 21970 1961 22004 1995
rect 22038 1961 22072 1995
rect 22106 1961 22140 1995
rect 22174 1961 22208 1995
rect 22242 1961 22276 1995
rect 22310 1961 22344 1995
rect 22378 1961 22412 1995
rect 22446 1961 22480 1995
rect 22514 1961 22548 1995
rect 22582 1961 22616 1995
rect 22650 1961 22684 1995
rect 22718 1961 22752 1995
rect 22786 1961 22820 1995
rect 22854 1961 22888 1995
rect 22922 1961 22956 1995
rect 22990 1961 23024 1995
rect 23058 1961 23092 1995
rect 23126 1961 23160 1995
rect 23194 1961 23228 1995
rect 23262 1961 23296 1995
rect 23330 1961 23364 1995
rect 23398 1961 23432 1995
rect 23466 1961 23500 1995
rect 23534 1961 23568 1995
rect 23602 1961 23636 1995
rect 23670 1961 23704 1995
rect 23738 1961 23772 1995
rect 23806 1961 23840 1995
rect 23874 1961 23908 1995
rect 23942 1961 23976 1995
rect 24010 1961 24044 1995
rect 24078 1961 24112 1995
rect 24146 1961 24180 1995
rect 24214 1961 24248 1995
rect 24282 1961 24316 1995
rect 24350 1961 24384 1995
rect 24418 1961 24452 1995
rect 24486 1961 24520 1995
rect 24554 1961 24588 1995
rect 24622 1961 24656 1995
rect 24690 1961 24724 1995
rect 24758 1961 24792 1995
rect 24826 1961 24860 1995
rect 24894 1961 24928 1995
rect 24962 1961 24996 1995
rect 25030 1961 25064 1995
rect 25098 1961 25132 1995
rect 25166 1961 25200 1995
rect 25234 1961 25268 1995
rect 25302 1961 25336 1995
rect 25370 1961 25404 1995
rect 25438 1961 25472 1995
rect 25506 1961 25540 1995
rect 25574 1961 25608 1995
rect 25642 1961 25676 1995
rect 25710 1961 25744 1995
rect 25778 1961 25812 1995
rect 25846 1961 25880 1995
rect 25914 1961 25948 1995
rect 25982 1961 26016 1995
rect 26050 1961 26084 1995
rect 26118 1961 26152 1995
rect 26186 1961 26220 1995
rect 26254 1961 26288 1995
rect 26322 1961 26356 1995
rect 26390 1961 26424 1995
rect 26458 1961 26492 1995
rect 26526 1961 26560 1995
rect 26594 1961 26628 1995
rect 26662 1961 26696 1995
rect 26730 1961 26764 1995
rect 26798 1961 26832 1995
rect 26866 1961 26900 1995
rect 26934 1961 26968 1995
rect 27002 1961 27036 1995
rect 27070 1961 27104 1995
rect 27138 1961 27172 1995
rect 27206 1961 27240 1995
rect 27274 1961 27308 1995
rect 27342 1961 27376 1995
rect 27410 1961 27444 1995
rect 27478 1961 27508 1995
rect 1795 1926 1801 1960
rect 1975 1959 27508 1961
rect 1795 1887 1805 1926
rect 1979 1925 27508 1959
rect 1975 1921 27508 1925
rect 1975 1887 2009 1921
rect 2043 1887 2078 1921
rect 2112 1887 2147 1921
rect 2181 1887 2216 1921
rect 2250 1887 2284 1921
rect 2318 1887 2352 1921
rect 2386 1887 2420 1921
rect 2454 1887 2488 1921
rect 2522 1887 2556 1921
rect 2590 1887 2624 1921
rect 2658 1887 2692 1921
rect 2726 1887 2760 1921
rect 2794 1887 2828 1921
rect 2862 1887 2896 1921
rect 2930 1887 2964 1921
rect 2998 1887 3032 1921
rect 3066 1887 3100 1921
rect 3134 1887 3168 1921
rect 3202 1887 3236 1921
rect 3270 1887 3304 1921
rect 3338 1887 3372 1921
rect 3406 1887 3440 1921
rect 3474 1887 3508 1921
rect 3542 1887 3576 1921
rect 3610 1887 3644 1921
rect 3678 1887 3712 1921
rect 3746 1887 3780 1921
rect 3814 1887 3848 1921
rect 3882 1887 3916 1921
rect 3950 1887 3984 1921
rect 4018 1887 4052 1921
rect 4086 1887 4120 1921
rect 4154 1887 4188 1921
rect 4222 1887 4256 1921
rect 4290 1887 4324 1921
rect 4358 1887 4392 1921
rect 4426 1887 4460 1921
rect 4494 1887 4528 1921
rect 4562 1887 4596 1921
rect 4630 1887 4664 1921
rect 4698 1887 4732 1921
rect 4766 1887 4800 1921
rect 4834 1887 4868 1921
rect 4902 1887 4936 1921
rect 4970 1887 5004 1921
rect 5038 1887 5072 1921
rect 5106 1887 5140 1921
rect 5174 1887 5208 1921
rect 5242 1887 5276 1921
rect 5310 1887 5344 1921
rect 5378 1887 5412 1921
rect 5446 1887 5480 1921
rect 5514 1887 5548 1921
rect 5582 1887 5616 1921
rect 5650 1887 5684 1921
rect 5718 1887 5752 1921
rect 5786 1887 5820 1921
rect 5854 1887 5888 1921
rect 5922 1887 5956 1921
rect 5990 1887 6024 1921
rect 6058 1887 6092 1921
rect 6126 1887 6160 1921
rect 6194 1887 6228 1921
rect 6262 1887 6296 1921
rect 6330 1887 6364 1921
rect 6398 1887 6432 1921
rect 6466 1887 6500 1921
rect 6534 1887 6568 1921
rect 6602 1887 6636 1921
rect 6670 1887 6704 1921
rect 6738 1887 6772 1921
rect 6806 1887 6840 1921
rect 6874 1887 6908 1921
rect 6942 1887 6976 1921
rect 7010 1887 7044 1921
rect 7078 1887 7112 1921
rect 7146 1887 7180 1921
rect 7214 1887 7248 1921
rect 7282 1887 7316 1921
rect 7350 1887 7384 1921
rect 7418 1887 7452 1921
rect 7486 1887 7520 1921
rect 7554 1887 7588 1921
rect 7622 1887 7656 1921
rect 7690 1887 7724 1921
rect 7758 1887 7792 1921
rect 7826 1887 7860 1921
rect 7894 1887 7928 1921
rect 7962 1887 7996 1921
rect 8030 1887 8064 1921
rect 8098 1887 8132 1921
rect 8166 1887 8200 1921
rect 8234 1887 8268 1921
rect 8302 1887 8336 1921
rect 8370 1887 8404 1921
rect 8438 1887 8472 1921
rect 8506 1887 8540 1921
rect 8574 1887 8608 1921
rect 8642 1887 8676 1921
rect 8710 1887 8744 1921
rect 8778 1887 8812 1921
rect 8846 1887 8880 1921
rect 8914 1887 8948 1921
rect 8982 1887 9016 1921
rect 9050 1887 9084 1921
rect 9118 1887 9152 1921
rect 9186 1887 9220 1921
rect 9254 1887 9288 1921
rect 9322 1887 9356 1921
rect 9390 1887 9424 1921
rect 9458 1887 9492 1921
rect 9526 1887 9560 1921
rect 9594 1887 9628 1921
rect 9662 1887 9696 1921
rect 9730 1887 9764 1921
rect 9798 1887 9832 1921
rect 9866 1887 9900 1921
rect 9934 1887 9968 1921
rect 10002 1887 10036 1921
rect 10070 1887 10104 1921
rect 10138 1887 10172 1921
rect 10206 1887 10240 1921
rect 10274 1887 10308 1921
rect 10342 1887 10376 1921
rect 10410 1887 10444 1921
rect 10478 1887 10512 1921
rect 10546 1887 10580 1921
rect 10614 1887 10648 1921
rect 10682 1887 10716 1921
rect 10750 1887 10784 1921
rect 10818 1887 10852 1921
rect 10886 1887 10920 1921
rect 10954 1887 10988 1921
rect 11022 1887 11056 1921
rect 11090 1887 11124 1921
rect 11158 1887 11192 1921
rect 11226 1887 11260 1921
rect 11294 1887 11328 1921
rect 11362 1887 11396 1921
rect 11430 1887 11464 1921
rect 11498 1887 11532 1921
rect 11566 1887 11600 1921
rect 11634 1887 11668 1921
rect 11702 1887 11736 1921
rect 11770 1887 11804 1921
rect 11838 1887 11872 1921
rect 11906 1887 11940 1921
rect 11974 1887 12008 1921
rect 12042 1887 12076 1921
rect 12110 1887 12144 1921
rect 12178 1887 12212 1921
rect 12246 1887 12280 1921
rect 12314 1887 12348 1921
rect 12382 1887 12416 1921
rect 12450 1887 12484 1921
rect 12518 1887 12552 1921
rect 12586 1887 12620 1921
rect 12654 1887 12688 1921
rect 12722 1887 12756 1921
rect 12790 1887 12824 1921
rect 12858 1887 12892 1921
rect 12926 1887 12960 1921
rect 12994 1887 13028 1921
rect 13062 1887 13096 1921
rect 13130 1887 13164 1921
rect 13198 1887 13232 1921
rect 13266 1887 13300 1921
rect 13334 1887 13368 1921
rect 13402 1887 13436 1921
rect 13470 1887 13504 1921
rect 13538 1887 13572 1921
rect 13606 1887 13640 1921
rect 13674 1887 13708 1921
rect 13742 1887 13776 1921
rect 13810 1887 13844 1921
rect 13878 1887 13912 1921
rect 13946 1887 13980 1921
rect 14014 1887 14048 1921
rect 14082 1887 14116 1921
rect 14150 1887 14184 1921
rect 14218 1887 14252 1921
rect 14286 1887 14320 1921
rect 14354 1887 14388 1921
rect 14422 1887 14456 1921
rect 14490 1887 14524 1921
rect 14558 1887 14592 1921
rect 14626 1887 14660 1921
rect 14694 1887 14728 1921
rect 14762 1887 14796 1921
rect 14830 1887 14864 1921
rect 14898 1887 14932 1921
rect 14966 1887 15000 1921
rect 15034 1887 15068 1921
rect 15102 1887 15136 1921
rect 15170 1887 15204 1921
rect 15238 1887 15272 1921
rect 15306 1887 15340 1921
rect 15374 1887 15408 1921
rect 15442 1887 15476 1921
rect 15510 1887 15544 1921
rect 15578 1887 15612 1921
rect 15646 1887 15680 1921
rect 15714 1887 15748 1921
rect 15782 1887 15816 1921
rect 15850 1887 15884 1921
rect 15918 1887 15952 1921
rect 15986 1887 16020 1921
rect 16054 1887 16088 1921
rect 16122 1887 16156 1921
rect 16190 1887 16224 1921
rect 16258 1887 16292 1921
rect 16326 1887 16360 1921
rect 16394 1887 16428 1921
rect 16462 1887 16496 1921
rect 16530 1887 16564 1921
rect 16598 1887 16632 1921
rect 16666 1887 16700 1921
rect 16734 1887 16768 1921
rect 16802 1887 16836 1921
rect 16870 1887 16904 1921
rect 16938 1887 16972 1921
rect 17006 1887 17040 1921
rect 17074 1887 17108 1921
rect 17142 1887 17176 1921
rect 17210 1887 17244 1921
rect 17278 1887 17312 1921
rect 17346 1887 17380 1921
rect 17414 1887 17448 1921
rect 17482 1887 17516 1921
rect 17550 1887 17584 1921
rect 17618 1887 17652 1921
rect 17686 1887 17720 1921
rect 17754 1887 17788 1921
rect 17822 1887 17856 1921
rect 17890 1887 17924 1921
rect 17958 1887 17992 1921
rect 18026 1887 18060 1921
rect 18094 1887 18128 1921
rect 18162 1887 18196 1921
rect 18230 1887 18264 1921
rect 18298 1887 18332 1921
rect 18366 1887 18400 1921
rect 18434 1887 18468 1921
rect 18502 1887 18536 1921
rect 18570 1887 18604 1921
rect 18638 1887 18672 1921
rect 18706 1887 18740 1921
rect 18774 1887 18808 1921
rect 18842 1887 18876 1921
rect 18910 1887 18944 1921
rect 18978 1887 19012 1921
rect 19046 1887 19080 1921
rect 19114 1887 19148 1921
rect 19182 1887 19216 1921
rect 19250 1887 19284 1921
rect 19318 1887 19352 1921
rect 19386 1887 19420 1921
rect 19454 1887 19488 1921
rect 19522 1887 19556 1921
rect 19590 1887 19624 1921
rect 19658 1887 19692 1921
rect 19726 1887 19760 1921
rect 19794 1887 19828 1921
rect 19862 1887 19896 1921
rect 19930 1887 19964 1921
rect 19998 1887 20032 1921
rect 20066 1887 20100 1921
rect 20134 1887 20168 1921
rect 20202 1887 20236 1921
rect 20270 1887 20304 1921
rect 20338 1887 20372 1921
rect 20406 1887 20440 1921
rect 20474 1887 20508 1921
rect 20542 1887 20576 1921
rect 20610 1887 20644 1921
rect 20678 1887 20712 1921
rect 20746 1887 20780 1921
rect 20814 1887 20848 1921
rect 20882 1887 20916 1921
rect 20950 1887 20984 1921
rect 21018 1887 21052 1921
rect 21086 1887 21120 1921
rect 21154 1887 21188 1921
rect 21222 1887 21256 1921
rect 21290 1887 21324 1921
rect 21358 1887 21392 1921
rect 21426 1887 21460 1921
rect 21494 1887 21528 1921
rect 21562 1887 21596 1921
rect 21630 1887 21664 1921
rect 21698 1887 21732 1921
rect 21766 1887 21800 1921
rect 21834 1887 21868 1921
rect 21902 1887 21936 1921
rect 21970 1887 22004 1921
rect 22038 1887 22072 1921
rect 22106 1887 22140 1921
rect 22174 1887 22208 1921
rect 22242 1887 22276 1921
rect 22310 1887 22344 1921
rect 22378 1887 22412 1921
rect 22446 1887 22480 1921
rect 22514 1887 22548 1921
rect 22582 1887 22616 1921
rect 22650 1887 22684 1921
rect 22718 1887 22752 1921
rect 22786 1887 22820 1921
rect 22854 1887 22888 1921
rect 22922 1887 22956 1921
rect 22990 1887 23024 1921
rect 23058 1887 23092 1921
rect 23126 1887 23160 1921
rect 23194 1887 23228 1921
rect 23262 1887 23296 1921
rect 23330 1887 23364 1921
rect 23398 1887 23432 1921
rect 23466 1887 23500 1921
rect 23534 1887 23568 1921
rect 23602 1887 23636 1921
rect 23670 1887 23704 1921
rect 23738 1887 23772 1921
rect 23806 1887 23840 1921
rect 23874 1887 23908 1921
rect 23942 1887 23976 1921
rect 24010 1887 24044 1921
rect 24078 1887 24112 1921
rect 24146 1887 24180 1921
rect 24214 1887 24248 1921
rect 24282 1887 24316 1921
rect 24350 1887 24384 1921
rect 24418 1887 24452 1921
rect 24486 1887 24520 1921
rect 24554 1887 24588 1921
rect 24622 1887 24656 1921
rect 24690 1887 24724 1921
rect 24758 1887 24792 1921
rect 24826 1887 24860 1921
rect 24894 1887 24928 1921
rect 24962 1887 24996 1921
rect 25030 1887 25064 1921
rect 25098 1887 25132 1921
rect 25166 1887 25200 1921
rect 25234 1887 25268 1921
rect 25302 1887 25336 1921
rect 25370 1887 25404 1921
rect 25438 1887 25472 1921
rect 25506 1887 25540 1921
rect 25574 1887 25608 1921
rect 25642 1887 25676 1921
rect 25710 1887 25744 1921
rect 25778 1887 25812 1921
rect 25846 1887 25880 1921
rect 25914 1887 25948 1921
rect 25982 1887 26016 1921
rect 26050 1887 26084 1921
rect 26118 1887 26152 1921
rect 26186 1887 26220 1921
rect 26254 1887 26288 1921
rect 26322 1887 26356 1921
rect 26390 1887 26424 1921
rect 26458 1887 26492 1921
rect 26526 1887 26560 1921
rect 26594 1887 26628 1921
rect 26662 1887 26696 1921
rect 26730 1887 26764 1921
rect 26798 1887 26832 1921
rect 26866 1887 26900 1921
rect 26934 1887 26968 1921
rect 27002 1887 27036 1921
rect 27070 1887 27104 1921
rect 27138 1887 27172 1921
rect 27206 1887 27240 1921
rect 27274 1887 27308 1921
rect 27342 1887 27376 1921
rect 27410 1887 27444 1921
rect 27478 1887 27508 1921
rect 1795 1853 1801 1887
rect 1975 1886 27508 1887
rect 1795 1814 1805 1853
rect 1979 1852 27508 1886
rect 1975 1847 27508 1852
rect 1795 1780 1801 1814
rect 1975 1813 2009 1847
rect 2043 1813 2078 1847
rect 2112 1813 2147 1847
rect 2181 1813 2216 1847
rect 2250 1813 2284 1847
rect 2318 1813 2352 1847
rect 2386 1813 2420 1847
rect 2454 1813 2488 1847
rect 2522 1813 2556 1847
rect 2590 1813 2624 1847
rect 2658 1813 2692 1847
rect 2726 1813 2760 1847
rect 2794 1813 2828 1847
rect 2862 1813 2896 1847
rect 2930 1813 2964 1847
rect 2998 1813 3032 1847
rect 3066 1813 3100 1847
rect 3134 1813 3168 1847
rect 3202 1813 3236 1847
rect 3270 1813 3304 1847
rect 3338 1813 3372 1847
rect 3406 1813 3440 1847
rect 3474 1813 3508 1847
rect 3542 1813 3576 1847
rect 3610 1813 3644 1847
rect 3678 1813 3712 1847
rect 3746 1813 3780 1847
rect 3814 1813 3848 1847
rect 3882 1813 3916 1847
rect 3950 1813 3984 1847
rect 4018 1813 4052 1847
rect 4086 1813 4120 1847
rect 4154 1813 4188 1847
rect 4222 1813 4256 1847
rect 4290 1813 4324 1847
rect 4358 1813 4392 1847
rect 4426 1813 4460 1847
rect 4494 1813 4528 1847
rect 4562 1813 4596 1847
rect 4630 1813 4664 1847
rect 4698 1813 4732 1847
rect 4766 1813 4800 1847
rect 4834 1813 4868 1847
rect 4902 1813 4936 1847
rect 4970 1813 5004 1847
rect 5038 1813 5072 1847
rect 5106 1813 5140 1847
rect 5174 1813 5208 1847
rect 5242 1813 5276 1847
rect 5310 1813 5344 1847
rect 5378 1813 5412 1847
rect 5446 1813 5480 1847
rect 5514 1813 5548 1847
rect 5582 1813 5616 1847
rect 5650 1813 5684 1847
rect 5718 1813 5752 1847
rect 5786 1813 5820 1847
rect 5854 1813 5888 1847
rect 5922 1813 5956 1847
rect 5990 1813 6024 1847
rect 6058 1813 6092 1847
rect 6126 1813 6160 1847
rect 6194 1813 6228 1847
rect 6262 1813 6296 1847
rect 6330 1813 6364 1847
rect 6398 1813 6432 1847
rect 6466 1813 6500 1847
rect 6534 1813 6568 1847
rect 6602 1813 6636 1847
rect 6670 1813 6704 1847
rect 6738 1813 6772 1847
rect 6806 1813 6840 1847
rect 6874 1813 6908 1847
rect 6942 1813 6976 1847
rect 7010 1813 7044 1847
rect 7078 1813 7112 1847
rect 7146 1813 7180 1847
rect 7214 1813 7248 1847
rect 7282 1813 7316 1847
rect 7350 1813 7384 1847
rect 7418 1813 7452 1847
rect 7486 1813 7520 1847
rect 7554 1813 7588 1847
rect 7622 1813 7656 1847
rect 7690 1813 7724 1847
rect 7758 1813 7792 1847
rect 7826 1813 7860 1847
rect 7894 1813 7928 1847
rect 7962 1813 7996 1847
rect 8030 1813 8064 1847
rect 8098 1813 8132 1847
rect 8166 1813 8200 1847
rect 8234 1813 8268 1847
rect 8302 1813 8336 1847
rect 8370 1813 8404 1847
rect 8438 1813 8472 1847
rect 8506 1813 8540 1847
rect 8574 1813 8608 1847
rect 8642 1813 8676 1847
rect 8710 1813 8744 1847
rect 8778 1813 8812 1847
rect 8846 1813 8880 1847
rect 8914 1813 8948 1847
rect 8982 1813 9016 1847
rect 9050 1813 9084 1847
rect 9118 1813 9152 1847
rect 9186 1813 9220 1847
rect 9254 1813 9288 1847
rect 9322 1813 9356 1847
rect 9390 1813 9424 1847
rect 9458 1813 9492 1847
rect 9526 1813 9560 1847
rect 9594 1813 9628 1847
rect 9662 1813 9696 1847
rect 9730 1813 9764 1847
rect 9798 1813 9832 1847
rect 9866 1813 9900 1847
rect 9934 1813 9968 1847
rect 10002 1813 10036 1847
rect 10070 1813 10104 1847
rect 10138 1813 10172 1847
rect 10206 1813 10240 1847
rect 10274 1813 10308 1847
rect 10342 1813 10376 1847
rect 10410 1813 10444 1847
rect 10478 1813 10512 1847
rect 10546 1813 10580 1847
rect 10614 1813 10648 1847
rect 10682 1813 10716 1847
rect 10750 1813 10784 1847
rect 10818 1813 10852 1847
rect 10886 1813 10920 1847
rect 10954 1813 10988 1847
rect 11022 1813 11056 1847
rect 11090 1813 11124 1847
rect 11158 1813 11192 1847
rect 11226 1813 11260 1847
rect 11294 1813 11328 1847
rect 11362 1813 11396 1847
rect 11430 1813 11464 1847
rect 11498 1813 11532 1847
rect 11566 1813 11600 1847
rect 11634 1813 11668 1847
rect 11702 1813 11736 1847
rect 11770 1813 11804 1847
rect 11838 1813 11872 1847
rect 11906 1813 11940 1847
rect 11974 1813 12008 1847
rect 12042 1813 12076 1847
rect 12110 1813 12144 1847
rect 12178 1813 12212 1847
rect 12246 1813 12280 1847
rect 12314 1813 12348 1847
rect 12382 1813 12416 1847
rect 12450 1813 12484 1847
rect 12518 1813 12552 1847
rect 12586 1813 12620 1847
rect 12654 1813 12688 1847
rect 12722 1813 12756 1847
rect 12790 1813 12824 1847
rect 12858 1813 12892 1847
rect 12926 1813 12960 1847
rect 12994 1813 13028 1847
rect 13062 1813 13096 1847
rect 13130 1813 13164 1847
rect 13198 1813 13232 1847
rect 13266 1813 13300 1847
rect 13334 1813 13368 1847
rect 13402 1813 13436 1847
rect 13470 1813 13504 1847
rect 13538 1813 13572 1847
rect 13606 1813 13640 1847
rect 13674 1813 13708 1847
rect 13742 1813 13776 1847
rect 13810 1813 13844 1847
rect 13878 1813 13912 1847
rect 13946 1813 13980 1847
rect 14014 1813 14048 1847
rect 14082 1813 14116 1847
rect 14150 1813 14184 1847
rect 14218 1813 14252 1847
rect 14286 1813 14320 1847
rect 14354 1813 14388 1847
rect 14422 1813 14456 1847
rect 14490 1813 14524 1847
rect 14558 1813 14592 1847
rect 14626 1813 14660 1847
rect 14694 1813 14728 1847
rect 14762 1813 14796 1847
rect 14830 1813 14864 1847
rect 14898 1813 14932 1847
rect 14966 1813 15000 1847
rect 15034 1813 15068 1847
rect 15102 1813 15136 1847
rect 15170 1813 15204 1847
rect 15238 1813 15272 1847
rect 15306 1813 15340 1847
rect 15374 1813 15408 1847
rect 15442 1813 15476 1847
rect 15510 1813 15544 1847
rect 15578 1813 15612 1847
rect 15646 1813 15680 1847
rect 15714 1813 15748 1847
rect 15782 1813 15816 1847
rect 15850 1813 15884 1847
rect 15918 1813 15952 1847
rect 15986 1813 16020 1847
rect 16054 1813 16088 1847
rect 16122 1813 16156 1847
rect 16190 1813 16224 1847
rect 16258 1813 16292 1847
rect 16326 1813 16360 1847
rect 16394 1813 16428 1847
rect 16462 1813 16496 1847
rect 16530 1813 16564 1847
rect 16598 1813 16632 1847
rect 16666 1813 16700 1847
rect 16734 1813 16768 1847
rect 16802 1813 16836 1847
rect 16870 1813 16904 1847
rect 16938 1813 16972 1847
rect 17006 1813 17040 1847
rect 17074 1813 17108 1847
rect 17142 1813 17176 1847
rect 17210 1813 17244 1847
rect 17278 1813 17312 1847
rect 17346 1813 17380 1847
rect 17414 1813 17448 1847
rect 17482 1813 17516 1847
rect 17550 1813 17584 1847
rect 17618 1813 17652 1847
rect 17686 1813 17720 1847
rect 17754 1813 17788 1847
rect 17822 1813 17856 1847
rect 17890 1813 17924 1847
rect 17958 1813 17992 1847
rect 18026 1813 18060 1847
rect 18094 1813 18128 1847
rect 18162 1813 18196 1847
rect 18230 1813 18264 1847
rect 18298 1813 18332 1847
rect 18366 1813 18400 1847
rect 18434 1813 18468 1847
rect 18502 1813 18536 1847
rect 18570 1813 18604 1847
rect 18638 1813 18672 1847
rect 18706 1813 18740 1847
rect 18774 1813 18808 1847
rect 18842 1813 18876 1847
rect 18910 1813 18944 1847
rect 18978 1813 19012 1847
rect 19046 1813 19080 1847
rect 19114 1813 19148 1847
rect 19182 1813 19216 1847
rect 19250 1813 19284 1847
rect 19318 1813 19352 1847
rect 19386 1813 19420 1847
rect 19454 1813 19488 1847
rect 19522 1813 19556 1847
rect 19590 1813 19624 1847
rect 19658 1813 19692 1847
rect 19726 1813 19760 1847
rect 19794 1813 19828 1847
rect 19862 1813 19896 1847
rect 19930 1813 19964 1847
rect 19998 1813 20032 1847
rect 20066 1813 20100 1847
rect 20134 1813 20168 1847
rect 20202 1813 20236 1847
rect 20270 1813 20304 1847
rect 20338 1813 20372 1847
rect 20406 1813 20440 1847
rect 20474 1813 20508 1847
rect 20542 1813 20576 1847
rect 20610 1813 20644 1847
rect 20678 1813 20712 1847
rect 20746 1813 20780 1847
rect 20814 1813 20848 1847
rect 20882 1813 20916 1847
rect 20950 1813 20984 1847
rect 21018 1813 21052 1847
rect 21086 1813 21120 1847
rect 21154 1813 21188 1847
rect 21222 1813 21256 1847
rect 21290 1813 21324 1847
rect 21358 1813 21392 1847
rect 21426 1813 21460 1847
rect 21494 1813 21528 1847
rect 21562 1813 21596 1847
rect 21630 1813 21664 1847
rect 21698 1813 21732 1847
rect 21766 1813 21800 1847
rect 21834 1813 21868 1847
rect 21902 1813 21936 1847
rect 21970 1813 22004 1847
rect 22038 1813 22072 1847
rect 22106 1813 22140 1847
rect 22174 1813 22208 1847
rect 22242 1813 22276 1847
rect 22310 1813 22344 1847
rect 22378 1813 22412 1847
rect 22446 1813 22480 1847
rect 22514 1813 22548 1847
rect 22582 1813 22616 1847
rect 22650 1813 22684 1847
rect 22718 1813 22752 1847
rect 22786 1813 22820 1847
rect 22854 1813 22888 1847
rect 22922 1813 22956 1847
rect 22990 1813 23024 1847
rect 23058 1813 23092 1847
rect 23126 1813 23160 1847
rect 23194 1813 23228 1847
rect 23262 1813 23296 1847
rect 23330 1813 23364 1847
rect 23398 1813 23432 1847
rect 23466 1813 23500 1847
rect 23534 1813 23568 1847
rect 23602 1813 23636 1847
rect 23670 1813 23704 1847
rect 23738 1813 23772 1847
rect 23806 1813 23840 1847
rect 23874 1813 23908 1847
rect 23942 1813 23976 1847
rect 24010 1813 24044 1847
rect 24078 1813 24112 1847
rect 24146 1813 24180 1847
rect 24214 1813 24248 1847
rect 24282 1813 24316 1847
rect 24350 1813 24384 1847
rect 24418 1813 24452 1847
rect 24486 1813 24520 1847
rect 24554 1813 24588 1847
rect 24622 1813 24656 1847
rect 24690 1813 24724 1847
rect 24758 1813 24792 1847
rect 24826 1813 24860 1847
rect 24894 1813 24928 1847
rect 24962 1813 24996 1847
rect 25030 1813 25064 1847
rect 25098 1813 25132 1847
rect 25166 1813 25200 1847
rect 25234 1813 25268 1847
rect 25302 1813 25336 1847
rect 25370 1813 25404 1847
rect 25438 1813 25472 1847
rect 25506 1813 25540 1847
rect 25574 1813 25608 1847
rect 25642 1813 25676 1847
rect 25710 1813 25744 1847
rect 25778 1813 25812 1847
rect 25846 1813 25880 1847
rect 25914 1813 25948 1847
rect 25982 1813 26016 1847
rect 26050 1813 26084 1847
rect 26118 1813 26152 1847
rect 26186 1813 26220 1847
rect 26254 1813 26288 1847
rect 26322 1813 26356 1847
rect 26390 1813 26424 1847
rect 26458 1813 26492 1847
rect 26526 1813 26560 1847
rect 26594 1813 26628 1847
rect 26662 1813 26696 1847
rect 26730 1813 26764 1847
rect 26798 1813 26832 1847
rect 26866 1813 26900 1847
rect 26934 1813 26968 1847
rect 27002 1813 27036 1847
rect 27070 1813 27104 1847
rect 27138 1813 27172 1847
rect 27206 1813 27240 1847
rect 27274 1813 27308 1847
rect 27342 1813 27376 1847
rect 27410 1813 27444 1847
rect 27478 1813 27508 1847
rect 1795 1741 1805 1780
rect 1979 1779 27508 1813
rect 1975 1773 27508 1779
rect 1795 1707 1801 1741
rect 1975 1740 2009 1773
rect 1795 1668 1805 1707
rect 1979 1739 2009 1740
rect 2043 1739 2078 1773
rect 2112 1739 2147 1773
rect 2181 1739 2216 1773
rect 2250 1739 2284 1773
rect 2318 1739 2352 1773
rect 2386 1739 2420 1773
rect 2454 1739 2488 1773
rect 2522 1739 2556 1773
rect 2590 1739 2624 1773
rect 2658 1739 2692 1773
rect 2726 1739 2760 1773
rect 2794 1739 2828 1773
rect 2862 1739 2896 1773
rect 2930 1739 2964 1773
rect 2998 1739 3032 1773
rect 3066 1739 3100 1773
rect 3134 1739 3168 1773
rect 3202 1739 3236 1773
rect 3270 1739 3304 1773
rect 3338 1739 3372 1773
rect 3406 1739 3440 1773
rect 3474 1739 3508 1773
rect 3542 1739 3576 1773
rect 3610 1739 3644 1773
rect 3678 1739 3712 1773
rect 3746 1739 3780 1773
rect 3814 1739 3848 1773
rect 3882 1739 3916 1773
rect 3950 1739 3984 1773
rect 4018 1739 4052 1773
rect 4086 1739 4120 1773
rect 4154 1739 4188 1773
rect 4222 1739 4256 1773
rect 4290 1739 4324 1773
rect 4358 1739 4392 1773
rect 4426 1739 4460 1773
rect 4494 1739 4528 1773
rect 4562 1739 4596 1773
rect 4630 1739 4664 1773
rect 4698 1739 4732 1773
rect 4766 1739 4800 1773
rect 4834 1739 4868 1773
rect 4902 1739 4936 1773
rect 4970 1739 5004 1773
rect 5038 1739 5072 1773
rect 5106 1739 5140 1773
rect 5174 1739 5208 1773
rect 5242 1739 5276 1773
rect 5310 1739 5344 1773
rect 5378 1739 5412 1773
rect 5446 1739 5480 1773
rect 5514 1739 5548 1773
rect 5582 1739 5616 1773
rect 5650 1739 5684 1773
rect 5718 1739 5752 1773
rect 5786 1739 5820 1773
rect 5854 1739 5888 1773
rect 5922 1739 5956 1773
rect 5990 1739 6024 1773
rect 6058 1739 6092 1773
rect 6126 1739 6160 1773
rect 6194 1739 6228 1773
rect 6262 1739 6296 1773
rect 6330 1739 6364 1773
rect 6398 1739 6432 1773
rect 6466 1739 6500 1773
rect 6534 1739 6568 1773
rect 6602 1739 6636 1773
rect 6670 1739 6704 1773
rect 6738 1739 6772 1773
rect 6806 1739 6840 1773
rect 6874 1739 6908 1773
rect 6942 1739 6976 1773
rect 7010 1739 7044 1773
rect 7078 1739 7112 1773
rect 7146 1739 7180 1773
rect 7214 1739 7248 1773
rect 7282 1739 7316 1773
rect 7350 1739 7384 1773
rect 7418 1739 7452 1773
rect 7486 1739 7520 1773
rect 7554 1739 7588 1773
rect 7622 1739 7656 1773
rect 7690 1739 7724 1773
rect 7758 1739 7792 1773
rect 7826 1739 7860 1773
rect 7894 1739 7928 1773
rect 7962 1739 7996 1773
rect 8030 1739 8064 1773
rect 8098 1739 8132 1773
rect 8166 1739 8200 1773
rect 8234 1739 8268 1773
rect 8302 1739 8336 1773
rect 8370 1739 8404 1773
rect 8438 1739 8472 1773
rect 8506 1739 8540 1773
rect 8574 1739 8608 1773
rect 8642 1739 8676 1773
rect 8710 1739 8744 1773
rect 8778 1739 8812 1773
rect 8846 1739 8880 1773
rect 8914 1739 8948 1773
rect 8982 1739 9016 1773
rect 9050 1739 9084 1773
rect 9118 1739 9152 1773
rect 9186 1739 9220 1773
rect 9254 1739 9288 1773
rect 9322 1739 9356 1773
rect 9390 1739 9424 1773
rect 9458 1739 9492 1773
rect 9526 1739 9560 1773
rect 9594 1739 9628 1773
rect 9662 1739 9696 1773
rect 9730 1739 9764 1773
rect 9798 1739 9832 1773
rect 9866 1739 9900 1773
rect 9934 1739 9968 1773
rect 10002 1739 10036 1773
rect 10070 1739 10104 1773
rect 10138 1739 10172 1773
rect 10206 1739 10240 1773
rect 10274 1739 10308 1773
rect 10342 1739 10376 1773
rect 10410 1739 10444 1773
rect 10478 1739 10512 1773
rect 10546 1739 10580 1773
rect 10614 1739 10648 1773
rect 10682 1739 10716 1773
rect 10750 1739 10784 1773
rect 10818 1739 10852 1773
rect 10886 1739 10920 1773
rect 10954 1739 10988 1773
rect 11022 1739 11056 1773
rect 11090 1739 11124 1773
rect 11158 1739 11192 1773
rect 11226 1739 11260 1773
rect 11294 1739 11328 1773
rect 11362 1739 11396 1773
rect 11430 1739 11464 1773
rect 11498 1739 11532 1773
rect 11566 1739 11600 1773
rect 11634 1739 11668 1773
rect 11702 1739 11736 1773
rect 11770 1739 11804 1773
rect 11838 1739 11872 1773
rect 11906 1739 11940 1773
rect 11974 1739 12008 1773
rect 12042 1739 12076 1773
rect 12110 1739 12144 1773
rect 12178 1739 12212 1773
rect 12246 1739 12280 1773
rect 12314 1739 12348 1773
rect 12382 1739 12416 1773
rect 12450 1739 12484 1773
rect 12518 1739 12552 1773
rect 12586 1739 12620 1773
rect 12654 1739 12688 1773
rect 12722 1739 12756 1773
rect 12790 1739 12824 1773
rect 12858 1739 12892 1773
rect 12926 1739 12960 1773
rect 12994 1739 13028 1773
rect 13062 1739 13096 1773
rect 13130 1739 13164 1773
rect 13198 1739 13232 1773
rect 13266 1739 13300 1773
rect 13334 1739 13368 1773
rect 13402 1739 13436 1773
rect 13470 1739 13504 1773
rect 13538 1739 13572 1773
rect 13606 1739 13640 1773
rect 13674 1739 13708 1773
rect 13742 1739 13776 1773
rect 13810 1739 13844 1773
rect 13878 1739 13912 1773
rect 13946 1739 13980 1773
rect 14014 1739 14048 1773
rect 14082 1739 14116 1773
rect 14150 1739 14184 1773
rect 14218 1739 14252 1773
rect 14286 1739 14320 1773
rect 14354 1739 14388 1773
rect 14422 1739 14456 1773
rect 14490 1739 14524 1773
rect 14558 1739 14592 1773
rect 14626 1739 14660 1773
rect 14694 1739 14728 1773
rect 14762 1739 14796 1773
rect 14830 1739 14864 1773
rect 14898 1739 14932 1773
rect 14966 1739 15000 1773
rect 15034 1739 15068 1773
rect 15102 1739 15136 1773
rect 15170 1739 15204 1773
rect 15238 1739 15272 1773
rect 15306 1739 15340 1773
rect 15374 1739 15408 1773
rect 15442 1739 15476 1773
rect 15510 1739 15544 1773
rect 15578 1739 15612 1773
rect 15646 1739 15680 1773
rect 15714 1739 15748 1773
rect 15782 1739 15816 1773
rect 15850 1739 15884 1773
rect 15918 1739 15952 1773
rect 15986 1739 16020 1773
rect 16054 1739 16088 1773
rect 16122 1739 16156 1773
rect 16190 1739 16224 1773
rect 16258 1739 16292 1773
rect 16326 1739 16360 1773
rect 16394 1739 16428 1773
rect 16462 1739 16496 1773
rect 16530 1739 16564 1773
rect 16598 1739 16632 1773
rect 16666 1739 16700 1773
rect 16734 1739 16768 1773
rect 16802 1739 16836 1773
rect 16870 1739 16904 1773
rect 16938 1739 16972 1773
rect 17006 1739 17040 1773
rect 17074 1739 17108 1773
rect 17142 1739 17176 1773
rect 17210 1739 17244 1773
rect 17278 1739 17312 1773
rect 17346 1739 17380 1773
rect 17414 1739 17448 1773
rect 17482 1739 17516 1773
rect 17550 1739 17584 1773
rect 17618 1739 17652 1773
rect 17686 1739 17720 1773
rect 17754 1739 17788 1773
rect 17822 1739 17856 1773
rect 17890 1739 17924 1773
rect 17958 1739 17992 1773
rect 18026 1739 18060 1773
rect 18094 1739 18128 1773
rect 18162 1739 18196 1773
rect 18230 1739 18264 1773
rect 18298 1739 18332 1773
rect 18366 1739 18400 1773
rect 18434 1739 18468 1773
rect 18502 1739 18536 1773
rect 18570 1739 18604 1773
rect 18638 1739 18672 1773
rect 18706 1739 18740 1773
rect 18774 1739 18808 1773
rect 18842 1739 18876 1773
rect 18910 1739 18944 1773
rect 18978 1739 19012 1773
rect 19046 1739 19080 1773
rect 19114 1739 19148 1773
rect 19182 1739 19216 1773
rect 19250 1739 19284 1773
rect 19318 1739 19352 1773
rect 19386 1739 19420 1773
rect 19454 1739 19488 1773
rect 19522 1739 19556 1773
rect 19590 1739 19624 1773
rect 19658 1739 19692 1773
rect 19726 1739 19760 1773
rect 19794 1739 19828 1773
rect 19862 1739 19896 1773
rect 19930 1739 19964 1773
rect 19998 1739 20032 1773
rect 20066 1739 20100 1773
rect 20134 1739 20168 1773
rect 20202 1739 20236 1773
rect 20270 1739 20304 1773
rect 20338 1739 20372 1773
rect 20406 1739 20440 1773
rect 20474 1739 20508 1773
rect 20542 1739 20576 1773
rect 20610 1739 20644 1773
rect 20678 1739 20712 1773
rect 20746 1739 20780 1773
rect 20814 1739 20848 1773
rect 20882 1739 20916 1773
rect 20950 1739 20984 1773
rect 21018 1739 21052 1773
rect 21086 1739 21120 1773
rect 21154 1739 21188 1773
rect 21222 1739 21256 1773
rect 21290 1739 21324 1773
rect 21358 1739 21392 1773
rect 21426 1739 21460 1773
rect 21494 1739 21528 1773
rect 21562 1739 21596 1773
rect 21630 1739 21664 1773
rect 21698 1739 21732 1773
rect 21766 1739 21800 1773
rect 21834 1739 21868 1773
rect 21902 1739 21936 1773
rect 21970 1739 22004 1773
rect 22038 1739 22072 1773
rect 22106 1739 22140 1773
rect 22174 1739 22208 1773
rect 22242 1739 22276 1773
rect 22310 1739 22344 1773
rect 22378 1739 22412 1773
rect 22446 1739 22480 1773
rect 22514 1739 22548 1773
rect 22582 1739 22616 1773
rect 22650 1739 22684 1773
rect 22718 1739 22752 1773
rect 22786 1739 22820 1773
rect 22854 1739 22888 1773
rect 22922 1739 22956 1773
rect 22990 1739 23024 1773
rect 23058 1739 23092 1773
rect 23126 1739 23160 1773
rect 23194 1739 23228 1773
rect 23262 1739 23296 1773
rect 23330 1739 23364 1773
rect 23398 1739 23432 1773
rect 23466 1739 23500 1773
rect 23534 1739 23568 1773
rect 23602 1739 23636 1773
rect 23670 1739 23704 1773
rect 23738 1739 23772 1773
rect 23806 1739 23840 1773
rect 23874 1739 23908 1773
rect 23942 1739 23976 1773
rect 24010 1739 24044 1773
rect 24078 1739 24112 1773
rect 24146 1739 24180 1773
rect 24214 1739 24248 1773
rect 24282 1739 24316 1773
rect 24350 1739 24384 1773
rect 24418 1739 24452 1773
rect 24486 1739 24520 1773
rect 24554 1739 24588 1773
rect 24622 1739 24656 1773
rect 24690 1739 24724 1773
rect 24758 1739 24792 1773
rect 24826 1739 24860 1773
rect 24894 1739 24928 1773
rect 24962 1739 24996 1773
rect 25030 1739 25064 1773
rect 25098 1739 25132 1773
rect 25166 1739 25200 1773
rect 25234 1739 25268 1773
rect 25302 1739 25336 1773
rect 25370 1739 25404 1773
rect 25438 1739 25472 1773
rect 25506 1739 25540 1773
rect 25574 1739 25608 1773
rect 25642 1739 25676 1773
rect 25710 1739 25744 1773
rect 25778 1739 25812 1773
rect 25846 1739 25880 1773
rect 25914 1739 25948 1773
rect 25982 1739 26016 1773
rect 26050 1739 26084 1773
rect 26118 1739 26152 1773
rect 26186 1739 26220 1773
rect 26254 1739 26288 1773
rect 26322 1739 26356 1773
rect 26390 1739 26424 1773
rect 26458 1739 26492 1773
rect 26526 1739 26560 1773
rect 26594 1739 26628 1773
rect 26662 1739 26696 1773
rect 26730 1739 26764 1773
rect 26798 1739 26832 1773
rect 26866 1739 26900 1773
rect 26934 1739 26968 1773
rect 27002 1739 27036 1773
rect 27070 1739 27104 1773
rect 27138 1739 27172 1773
rect 27206 1739 27240 1773
rect 27274 1739 27308 1773
rect 27342 1739 27376 1773
rect 27410 1739 27444 1773
rect 27478 1739 27508 1773
rect 1979 1706 27508 1739
rect 1975 1699 27508 1706
rect 1795 1634 1801 1668
rect 1975 1667 2009 1699
rect 1795 1595 1805 1634
rect 1979 1665 2009 1667
rect 2043 1665 2078 1699
rect 2112 1665 2147 1699
rect 2181 1665 2216 1699
rect 2250 1665 2284 1699
rect 2318 1665 2352 1699
rect 2386 1665 2420 1699
rect 2454 1665 2488 1699
rect 2522 1665 2556 1699
rect 2590 1665 2624 1699
rect 2658 1665 2692 1699
rect 2726 1665 2760 1699
rect 2794 1665 2828 1699
rect 2862 1665 2896 1699
rect 2930 1665 2964 1699
rect 2998 1665 3032 1699
rect 3066 1665 3100 1699
rect 3134 1665 3168 1699
rect 3202 1665 3236 1699
rect 3270 1665 3304 1699
rect 3338 1665 3372 1699
rect 3406 1665 3440 1699
rect 3474 1665 3508 1699
rect 3542 1665 3576 1699
rect 3610 1665 3644 1699
rect 3678 1665 3712 1699
rect 3746 1665 3780 1699
rect 3814 1665 3848 1699
rect 3882 1665 3916 1699
rect 3950 1665 3984 1699
rect 4018 1665 4052 1699
rect 4086 1665 4120 1699
rect 4154 1665 4188 1699
rect 4222 1665 4256 1699
rect 4290 1665 4324 1699
rect 4358 1665 4392 1699
rect 4426 1665 4460 1699
rect 4494 1665 4528 1699
rect 4562 1665 4596 1699
rect 4630 1665 4664 1699
rect 4698 1665 4732 1699
rect 4766 1665 4800 1699
rect 4834 1665 4868 1699
rect 4902 1665 4936 1699
rect 4970 1665 5004 1699
rect 5038 1665 5072 1699
rect 5106 1665 5140 1699
rect 5174 1665 5208 1699
rect 5242 1665 5276 1699
rect 5310 1665 5344 1699
rect 5378 1665 5412 1699
rect 5446 1665 5480 1699
rect 5514 1665 5548 1699
rect 5582 1665 5616 1699
rect 5650 1665 5684 1699
rect 5718 1665 5752 1699
rect 5786 1665 5820 1699
rect 5854 1665 5888 1699
rect 5922 1665 5956 1699
rect 5990 1665 6024 1699
rect 6058 1665 6092 1699
rect 6126 1665 6160 1699
rect 6194 1665 6228 1699
rect 6262 1665 6296 1699
rect 6330 1665 6364 1699
rect 6398 1665 6432 1699
rect 6466 1665 6500 1699
rect 6534 1665 6568 1699
rect 6602 1665 6636 1699
rect 6670 1665 6704 1699
rect 6738 1665 6772 1699
rect 6806 1665 6840 1699
rect 6874 1665 6908 1699
rect 6942 1665 6976 1699
rect 7010 1665 7044 1699
rect 7078 1665 7112 1699
rect 7146 1665 7180 1699
rect 7214 1665 7248 1699
rect 7282 1665 7316 1699
rect 7350 1665 7384 1699
rect 7418 1665 7452 1699
rect 7486 1665 7520 1699
rect 7554 1665 7588 1699
rect 7622 1665 7656 1699
rect 7690 1665 7724 1699
rect 7758 1665 7792 1699
rect 7826 1665 7860 1699
rect 7894 1665 7928 1699
rect 7962 1665 7996 1699
rect 8030 1665 8064 1699
rect 8098 1665 8132 1699
rect 8166 1665 8200 1699
rect 8234 1665 8268 1699
rect 8302 1665 8336 1699
rect 8370 1665 8404 1699
rect 8438 1665 8472 1699
rect 8506 1665 8540 1699
rect 8574 1665 8608 1699
rect 8642 1665 8676 1699
rect 8710 1665 8744 1699
rect 8778 1665 8812 1699
rect 8846 1665 8880 1699
rect 8914 1665 8948 1699
rect 8982 1665 9016 1699
rect 9050 1665 9084 1699
rect 9118 1665 9152 1699
rect 9186 1665 9220 1699
rect 9254 1665 9288 1699
rect 9322 1665 9356 1699
rect 9390 1665 9424 1699
rect 9458 1665 9492 1699
rect 9526 1665 9560 1699
rect 9594 1665 9628 1699
rect 9662 1665 9696 1699
rect 9730 1665 9764 1699
rect 9798 1665 9832 1699
rect 9866 1665 9900 1699
rect 9934 1665 9968 1699
rect 10002 1665 10036 1699
rect 10070 1665 10104 1699
rect 10138 1665 10172 1699
rect 10206 1665 10240 1699
rect 10274 1665 10308 1699
rect 10342 1665 10376 1699
rect 10410 1665 10444 1699
rect 10478 1665 10512 1699
rect 10546 1665 10580 1699
rect 10614 1665 10648 1699
rect 10682 1665 10716 1699
rect 10750 1665 10784 1699
rect 10818 1665 10852 1699
rect 10886 1665 10920 1699
rect 10954 1665 10988 1699
rect 11022 1665 11056 1699
rect 11090 1665 11124 1699
rect 11158 1665 11192 1699
rect 11226 1665 11260 1699
rect 11294 1665 11328 1699
rect 11362 1665 11396 1699
rect 11430 1665 11464 1699
rect 11498 1665 11532 1699
rect 11566 1665 11600 1699
rect 11634 1665 11668 1699
rect 11702 1665 11736 1699
rect 11770 1665 11804 1699
rect 11838 1665 11872 1699
rect 11906 1665 11940 1699
rect 11974 1665 12008 1699
rect 12042 1665 12076 1699
rect 12110 1665 12144 1699
rect 12178 1665 12212 1699
rect 12246 1665 12280 1699
rect 12314 1665 12348 1699
rect 12382 1665 12416 1699
rect 12450 1665 12484 1699
rect 12518 1665 12552 1699
rect 12586 1665 12620 1699
rect 12654 1665 12688 1699
rect 12722 1665 12756 1699
rect 12790 1665 12824 1699
rect 12858 1665 12892 1699
rect 12926 1665 12960 1699
rect 12994 1665 13028 1699
rect 13062 1665 13096 1699
rect 13130 1665 13164 1699
rect 13198 1665 13232 1699
rect 13266 1665 13300 1699
rect 13334 1665 13368 1699
rect 13402 1665 13436 1699
rect 13470 1665 13504 1699
rect 13538 1665 13572 1699
rect 13606 1665 13640 1699
rect 13674 1665 13708 1699
rect 13742 1665 13776 1699
rect 13810 1665 13844 1699
rect 13878 1665 13912 1699
rect 13946 1665 13980 1699
rect 14014 1665 14048 1699
rect 14082 1665 14116 1699
rect 14150 1665 14184 1699
rect 14218 1665 14252 1699
rect 14286 1665 14320 1699
rect 14354 1665 14388 1699
rect 14422 1665 14456 1699
rect 14490 1665 14524 1699
rect 14558 1665 14592 1699
rect 14626 1665 14660 1699
rect 14694 1665 14728 1699
rect 14762 1665 14796 1699
rect 14830 1665 14864 1699
rect 14898 1665 14932 1699
rect 14966 1665 15000 1699
rect 15034 1665 15068 1699
rect 15102 1665 15136 1699
rect 15170 1665 15204 1699
rect 15238 1665 15272 1699
rect 15306 1665 15340 1699
rect 15374 1665 15408 1699
rect 15442 1665 15476 1699
rect 15510 1665 15544 1699
rect 15578 1665 15612 1699
rect 15646 1665 15680 1699
rect 15714 1665 15748 1699
rect 15782 1665 15816 1699
rect 15850 1665 15884 1699
rect 15918 1665 15952 1699
rect 15986 1665 16020 1699
rect 16054 1665 16088 1699
rect 16122 1665 16156 1699
rect 16190 1665 16224 1699
rect 16258 1665 16292 1699
rect 16326 1665 16360 1699
rect 16394 1665 16428 1699
rect 16462 1665 16496 1699
rect 16530 1665 16564 1699
rect 16598 1665 16632 1699
rect 16666 1665 16700 1699
rect 16734 1665 16768 1699
rect 16802 1665 16836 1699
rect 16870 1665 16904 1699
rect 16938 1665 16972 1699
rect 17006 1665 17040 1699
rect 17074 1665 17108 1699
rect 17142 1665 17176 1699
rect 17210 1665 17244 1699
rect 17278 1665 17312 1699
rect 17346 1665 17380 1699
rect 17414 1665 17448 1699
rect 17482 1665 17516 1699
rect 17550 1665 17584 1699
rect 17618 1665 17652 1699
rect 17686 1665 17720 1699
rect 17754 1665 17788 1699
rect 17822 1665 17856 1699
rect 17890 1665 17924 1699
rect 17958 1665 17992 1699
rect 18026 1665 18060 1699
rect 18094 1665 18128 1699
rect 18162 1665 18196 1699
rect 18230 1665 18264 1699
rect 18298 1665 18332 1699
rect 18366 1665 18400 1699
rect 18434 1665 18468 1699
rect 18502 1665 18536 1699
rect 18570 1665 18604 1699
rect 18638 1665 18672 1699
rect 18706 1665 18740 1699
rect 18774 1665 18808 1699
rect 18842 1665 18876 1699
rect 18910 1665 18944 1699
rect 18978 1665 19012 1699
rect 19046 1665 19080 1699
rect 19114 1665 19148 1699
rect 19182 1665 19216 1699
rect 19250 1665 19284 1699
rect 19318 1665 19352 1699
rect 19386 1665 19420 1699
rect 19454 1665 19488 1699
rect 19522 1665 19556 1699
rect 19590 1665 19624 1699
rect 19658 1665 19692 1699
rect 19726 1665 19760 1699
rect 19794 1665 19828 1699
rect 19862 1665 19896 1699
rect 19930 1665 19964 1699
rect 19998 1665 20032 1699
rect 20066 1665 20100 1699
rect 20134 1665 20168 1699
rect 20202 1665 20236 1699
rect 20270 1665 20304 1699
rect 20338 1665 20372 1699
rect 20406 1665 20440 1699
rect 20474 1665 20508 1699
rect 20542 1665 20576 1699
rect 20610 1665 20644 1699
rect 20678 1665 20712 1699
rect 20746 1665 20780 1699
rect 20814 1665 20848 1699
rect 20882 1665 20916 1699
rect 20950 1665 20984 1699
rect 21018 1665 21052 1699
rect 21086 1665 21120 1699
rect 21154 1665 21188 1699
rect 21222 1665 21256 1699
rect 21290 1665 21324 1699
rect 21358 1665 21392 1699
rect 21426 1665 21460 1699
rect 21494 1665 21528 1699
rect 21562 1665 21596 1699
rect 21630 1665 21664 1699
rect 21698 1665 21732 1699
rect 21766 1665 21800 1699
rect 21834 1665 21868 1699
rect 21902 1665 21936 1699
rect 21970 1665 22004 1699
rect 22038 1665 22072 1699
rect 22106 1665 22140 1699
rect 22174 1665 22208 1699
rect 22242 1665 22276 1699
rect 22310 1665 22344 1699
rect 22378 1665 22412 1699
rect 22446 1665 22480 1699
rect 22514 1665 22548 1699
rect 22582 1665 22616 1699
rect 22650 1665 22684 1699
rect 22718 1665 22752 1699
rect 22786 1665 22820 1699
rect 22854 1665 22888 1699
rect 22922 1665 22956 1699
rect 22990 1665 23024 1699
rect 23058 1665 23092 1699
rect 23126 1665 23160 1699
rect 23194 1665 23228 1699
rect 23262 1665 23296 1699
rect 23330 1665 23364 1699
rect 23398 1665 23432 1699
rect 23466 1665 23500 1699
rect 23534 1665 23568 1699
rect 23602 1665 23636 1699
rect 23670 1665 23704 1699
rect 23738 1665 23772 1699
rect 23806 1665 23840 1699
rect 23874 1665 23908 1699
rect 23942 1665 23976 1699
rect 24010 1665 24044 1699
rect 24078 1665 24112 1699
rect 24146 1665 24180 1699
rect 24214 1665 24248 1699
rect 24282 1665 24316 1699
rect 24350 1665 24384 1699
rect 24418 1665 24452 1699
rect 24486 1665 24520 1699
rect 24554 1665 24588 1699
rect 24622 1665 24656 1699
rect 24690 1665 24724 1699
rect 24758 1665 24792 1699
rect 24826 1665 24860 1699
rect 24894 1665 24928 1699
rect 24962 1665 24996 1699
rect 25030 1665 25064 1699
rect 25098 1665 25132 1699
rect 25166 1665 25200 1699
rect 25234 1665 25268 1699
rect 25302 1665 25336 1699
rect 25370 1665 25404 1699
rect 25438 1665 25472 1699
rect 25506 1665 25540 1699
rect 25574 1665 25608 1699
rect 25642 1665 25676 1699
rect 25710 1665 25744 1699
rect 25778 1665 25812 1699
rect 25846 1665 25880 1699
rect 25914 1665 25948 1699
rect 25982 1665 26016 1699
rect 26050 1665 26084 1699
rect 26118 1665 26152 1699
rect 26186 1665 26220 1699
rect 26254 1665 26288 1699
rect 26322 1665 26356 1699
rect 26390 1665 26424 1699
rect 26458 1665 26492 1699
rect 26526 1665 26560 1699
rect 26594 1665 26628 1699
rect 26662 1665 26696 1699
rect 26730 1665 26764 1699
rect 26798 1665 26832 1699
rect 26866 1665 26900 1699
rect 26934 1665 26968 1699
rect 27002 1665 27036 1699
rect 27070 1665 27104 1699
rect 27138 1665 27172 1699
rect 27206 1665 27240 1699
rect 27274 1665 27308 1699
rect 27342 1665 27376 1699
rect 27410 1665 27444 1699
rect 27478 1665 27508 1699
rect 1979 1633 27508 1665
rect 1975 1625 27508 1633
rect 1795 1561 1801 1595
rect 1975 1594 2009 1625
rect 1795 1522 1805 1561
rect 1979 1591 2009 1594
rect 2043 1591 2078 1625
rect 2112 1591 2147 1625
rect 2181 1591 2216 1625
rect 2250 1591 2284 1625
rect 2318 1591 2352 1625
rect 2386 1591 2420 1625
rect 2454 1591 2488 1625
rect 2522 1591 2556 1625
rect 2590 1591 2624 1625
rect 2658 1591 2692 1625
rect 2726 1591 2760 1625
rect 2794 1591 2828 1625
rect 2862 1591 2896 1625
rect 2930 1591 2964 1625
rect 2998 1591 3032 1625
rect 3066 1591 3100 1625
rect 3134 1591 3168 1625
rect 3202 1591 3236 1625
rect 3270 1591 3304 1625
rect 3338 1591 3372 1625
rect 3406 1591 3440 1625
rect 3474 1591 3508 1625
rect 3542 1591 3576 1625
rect 3610 1591 3644 1625
rect 3678 1591 3712 1625
rect 3746 1591 3780 1625
rect 3814 1591 3848 1625
rect 3882 1591 3916 1625
rect 3950 1591 3984 1625
rect 4018 1591 4052 1625
rect 4086 1591 4120 1625
rect 4154 1591 4188 1625
rect 4222 1591 4256 1625
rect 4290 1591 4324 1625
rect 4358 1591 4392 1625
rect 4426 1591 4460 1625
rect 4494 1591 4528 1625
rect 4562 1591 4596 1625
rect 4630 1591 4664 1625
rect 4698 1591 4732 1625
rect 4766 1591 4800 1625
rect 4834 1591 4868 1625
rect 4902 1591 4936 1625
rect 4970 1591 5004 1625
rect 5038 1591 5072 1625
rect 5106 1591 5140 1625
rect 5174 1591 5208 1625
rect 5242 1591 5276 1625
rect 5310 1591 5344 1625
rect 5378 1591 5412 1625
rect 5446 1591 5480 1625
rect 5514 1591 5548 1625
rect 5582 1591 5616 1625
rect 5650 1591 5684 1625
rect 5718 1591 5752 1625
rect 5786 1591 5820 1625
rect 5854 1591 5888 1625
rect 5922 1591 5956 1625
rect 5990 1591 6024 1625
rect 6058 1591 6092 1625
rect 6126 1591 6160 1625
rect 6194 1591 6228 1625
rect 6262 1591 6296 1625
rect 6330 1591 6364 1625
rect 6398 1591 6432 1625
rect 6466 1591 6500 1625
rect 6534 1591 6568 1625
rect 6602 1591 6636 1625
rect 6670 1591 6704 1625
rect 6738 1591 6772 1625
rect 6806 1591 6840 1625
rect 6874 1591 6908 1625
rect 6942 1591 6976 1625
rect 7010 1591 7044 1625
rect 7078 1591 7112 1625
rect 7146 1591 7180 1625
rect 7214 1591 7248 1625
rect 7282 1591 7316 1625
rect 7350 1591 7384 1625
rect 7418 1591 7452 1625
rect 7486 1591 7520 1625
rect 7554 1591 7588 1625
rect 7622 1591 7656 1625
rect 7690 1591 7724 1625
rect 7758 1591 7792 1625
rect 7826 1591 7860 1625
rect 7894 1591 7928 1625
rect 7962 1591 7996 1625
rect 8030 1591 8064 1625
rect 8098 1591 8132 1625
rect 8166 1591 8200 1625
rect 8234 1591 8268 1625
rect 8302 1591 8336 1625
rect 8370 1591 8404 1625
rect 8438 1591 8472 1625
rect 8506 1591 8540 1625
rect 8574 1591 8608 1625
rect 8642 1591 8676 1625
rect 8710 1591 8744 1625
rect 8778 1591 8812 1625
rect 8846 1591 8880 1625
rect 8914 1591 8948 1625
rect 8982 1591 9016 1625
rect 9050 1591 9084 1625
rect 9118 1591 9152 1625
rect 9186 1591 9220 1625
rect 9254 1591 9288 1625
rect 9322 1591 9356 1625
rect 9390 1591 9424 1625
rect 9458 1591 9492 1625
rect 9526 1591 9560 1625
rect 9594 1591 9628 1625
rect 9662 1591 9696 1625
rect 9730 1591 9764 1625
rect 9798 1591 9832 1625
rect 9866 1591 9900 1625
rect 9934 1591 9968 1625
rect 10002 1591 10036 1625
rect 10070 1591 10104 1625
rect 10138 1591 10172 1625
rect 10206 1591 10240 1625
rect 10274 1591 10308 1625
rect 10342 1591 10376 1625
rect 10410 1591 10444 1625
rect 10478 1591 10512 1625
rect 10546 1591 10580 1625
rect 10614 1591 10648 1625
rect 10682 1591 10716 1625
rect 10750 1591 10784 1625
rect 10818 1591 10852 1625
rect 10886 1591 10920 1625
rect 10954 1591 10988 1625
rect 11022 1591 11056 1625
rect 11090 1591 11124 1625
rect 11158 1591 11192 1625
rect 11226 1591 11260 1625
rect 11294 1591 11328 1625
rect 11362 1591 11396 1625
rect 11430 1591 11464 1625
rect 11498 1591 11532 1625
rect 11566 1591 11600 1625
rect 11634 1591 11668 1625
rect 11702 1591 11736 1625
rect 11770 1591 11804 1625
rect 11838 1591 11872 1625
rect 11906 1591 11940 1625
rect 11974 1591 12008 1625
rect 12042 1591 12076 1625
rect 12110 1591 12144 1625
rect 12178 1591 12212 1625
rect 12246 1591 12280 1625
rect 12314 1591 12348 1625
rect 12382 1591 12416 1625
rect 12450 1591 12484 1625
rect 12518 1591 12552 1625
rect 12586 1591 12620 1625
rect 12654 1591 12688 1625
rect 12722 1591 12756 1625
rect 12790 1591 12824 1625
rect 12858 1591 12892 1625
rect 12926 1591 12960 1625
rect 12994 1591 13028 1625
rect 13062 1591 13096 1625
rect 13130 1591 13164 1625
rect 13198 1591 13232 1625
rect 13266 1591 13300 1625
rect 13334 1591 13368 1625
rect 13402 1591 13436 1625
rect 13470 1591 13504 1625
rect 13538 1591 13572 1625
rect 13606 1591 13640 1625
rect 13674 1591 13708 1625
rect 13742 1591 13776 1625
rect 13810 1591 13844 1625
rect 13878 1591 13912 1625
rect 13946 1591 13980 1625
rect 14014 1591 14048 1625
rect 14082 1591 14116 1625
rect 14150 1591 14184 1625
rect 14218 1591 14252 1625
rect 14286 1591 14320 1625
rect 14354 1591 14388 1625
rect 14422 1591 14456 1625
rect 14490 1591 14524 1625
rect 14558 1591 14592 1625
rect 14626 1591 14660 1625
rect 14694 1591 14728 1625
rect 14762 1591 14796 1625
rect 14830 1591 14864 1625
rect 14898 1591 14932 1625
rect 14966 1591 15000 1625
rect 15034 1591 15068 1625
rect 15102 1591 15136 1625
rect 15170 1591 15204 1625
rect 15238 1591 15272 1625
rect 15306 1591 15340 1625
rect 15374 1591 15408 1625
rect 15442 1591 15476 1625
rect 15510 1591 15544 1625
rect 15578 1591 15612 1625
rect 15646 1591 15680 1625
rect 15714 1591 15748 1625
rect 15782 1591 15816 1625
rect 15850 1591 15884 1625
rect 15918 1591 15952 1625
rect 15986 1591 16020 1625
rect 16054 1591 16088 1625
rect 16122 1591 16156 1625
rect 16190 1591 16224 1625
rect 16258 1591 16292 1625
rect 16326 1591 16360 1625
rect 16394 1591 16428 1625
rect 16462 1591 16496 1625
rect 16530 1591 16564 1625
rect 16598 1591 16632 1625
rect 16666 1591 16700 1625
rect 16734 1591 16768 1625
rect 16802 1591 16836 1625
rect 16870 1591 16904 1625
rect 16938 1591 16972 1625
rect 17006 1591 17040 1625
rect 17074 1591 17108 1625
rect 17142 1591 17176 1625
rect 17210 1591 17244 1625
rect 17278 1591 17312 1625
rect 17346 1591 17380 1625
rect 17414 1591 17448 1625
rect 17482 1591 17516 1625
rect 17550 1591 17584 1625
rect 17618 1591 17652 1625
rect 17686 1591 17720 1625
rect 17754 1591 17788 1625
rect 17822 1591 17856 1625
rect 17890 1591 17924 1625
rect 17958 1591 17992 1625
rect 18026 1591 18060 1625
rect 18094 1591 18128 1625
rect 18162 1591 18196 1625
rect 18230 1591 18264 1625
rect 18298 1591 18332 1625
rect 18366 1591 18400 1625
rect 18434 1591 18468 1625
rect 18502 1591 18536 1625
rect 18570 1591 18604 1625
rect 18638 1591 18672 1625
rect 18706 1591 18740 1625
rect 18774 1591 18808 1625
rect 18842 1591 18876 1625
rect 18910 1591 18944 1625
rect 18978 1591 19012 1625
rect 19046 1591 19080 1625
rect 19114 1591 19148 1625
rect 19182 1591 19216 1625
rect 19250 1591 19284 1625
rect 19318 1591 19352 1625
rect 19386 1591 19420 1625
rect 19454 1591 19488 1625
rect 19522 1591 19556 1625
rect 19590 1591 19624 1625
rect 19658 1591 19692 1625
rect 19726 1591 19760 1625
rect 19794 1591 19828 1625
rect 19862 1591 19896 1625
rect 19930 1591 19964 1625
rect 19998 1591 20032 1625
rect 20066 1591 20100 1625
rect 20134 1591 20168 1625
rect 20202 1591 20236 1625
rect 20270 1591 20304 1625
rect 20338 1591 20372 1625
rect 20406 1591 20440 1625
rect 20474 1591 20508 1625
rect 20542 1591 20576 1625
rect 20610 1591 20644 1625
rect 20678 1591 20712 1625
rect 20746 1591 20780 1625
rect 20814 1591 20848 1625
rect 20882 1591 20916 1625
rect 20950 1591 20984 1625
rect 21018 1591 21052 1625
rect 21086 1591 21120 1625
rect 21154 1591 21188 1625
rect 21222 1591 21256 1625
rect 21290 1591 21324 1625
rect 21358 1591 21392 1625
rect 21426 1591 21460 1625
rect 21494 1591 21528 1625
rect 21562 1591 21596 1625
rect 21630 1591 21664 1625
rect 21698 1591 21732 1625
rect 21766 1591 21800 1625
rect 21834 1591 21868 1625
rect 21902 1591 21936 1625
rect 21970 1591 22004 1625
rect 22038 1591 22072 1625
rect 22106 1591 22140 1625
rect 22174 1591 22208 1625
rect 22242 1591 22276 1625
rect 22310 1591 22344 1625
rect 22378 1591 22412 1625
rect 22446 1591 22480 1625
rect 22514 1591 22548 1625
rect 22582 1591 22616 1625
rect 22650 1591 22684 1625
rect 22718 1591 22752 1625
rect 22786 1591 22820 1625
rect 22854 1591 22888 1625
rect 22922 1591 22956 1625
rect 22990 1591 23024 1625
rect 23058 1591 23092 1625
rect 23126 1591 23160 1625
rect 23194 1591 23228 1625
rect 23262 1591 23296 1625
rect 23330 1591 23364 1625
rect 23398 1591 23432 1625
rect 23466 1591 23500 1625
rect 23534 1591 23568 1625
rect 23602 1591 23636 1625
rect 23670 1591 23704 1625
rect 23738 1591 23772 1625
rect 23806 1591 23840 1625
rect 23874 1591 23908 1625
rect 23942 1591 23976 1625
rect 24010 1591 24044 1625
rect 24078 1591 24112 1625
rect 24146 1591 24180 1625
rect 24214 1591 24248 1625
rect 24282 1591 24316 1625
rect 24350 1591 24384 1625
rect 24418 1591 24452 1625
rect 24486 1591 24520 1625
rect 24554 1591 24588 1625
rect 24622 1591 24656 1625
rect 24690 1591 24724 1625
rect 24758 1591 24792 1625
rect 24826 1591 24860 1625
rect 24894 1591 24928 1625
rect 24962 1591 24996 1625
rect 25030 1591 25064 1625
rect 25098 1591 25132 1625
rect 25166 1591 25200 1625
rect 25234 1591 25268 1625
rect 25302 1591 25336 1625
rect 25370 1591 25404 1625
rect 25438 1591 25472 1625
rect 25506 1591 25540 1625
rect 25574 1591 25608 1625
rect 25642 1591 25676 1625
rect 25710 1591 25744 1625
rect 25778 1591 25812 1625
rect 25846 1591 25880 1625
rect 25914 1591 25948 1625
rect 25982 1591 26016 1625
rect 26050 1591 26084 1625
rect 26118 1591 26152 1625
rect 26186 1591 26220 1625
rect 26254 1591 26288 1625
rect 26322 1591 26356 1625
rect 26390 1591 26424 1625
rect 26458 1591 26492 1625
rect 26526 1591 26560 1625
rect 26594 1591 26628 1625
rect 26662 1591 26696 1625
rect 26730 1591 26764 1625
rect 26798 1591 26832 1625
rect 26866 1591 26900 1625
rect 26934 1591 26968 1625
rect 27002 1591 27036 1625
rect 27070 1591 27104 1625
rect 27138 1591 27172 1625
rect 27206 1591 27240 1625
rect 27274 1591 27308 1625
rect 27342 1591 27376 1625
rect 27410 1591 27444 1625
rect 27478 1591 27508 1625
rect 1979 1560 27508 1591
rect 1975 1551 27508 1560
rect 1795 1488 1801 1522
rect 1975 1521 2009 1551
rect 1795 1449 1805 1488
rect 1979 1517 2009 1521
rect 2043 1517 2078 1551
rect 2112 1517 2147 1551
rect 2181 1517 2216 1551
rect 2250 1517 2284 1551
rect 2318 1517 2352 1551
rect 2386 1517 2420 1551
rect 2454 1517 2488 1551
rect 2522 1517 2556 1551
rect 2590 1517 2624 1551
rect 2658 1517 2692 1551
rect 2726 1517 2760 1551
rect 2794 1517 2828 1551
rect 2862 1517 2896 1551
rect 2930 1517 2964 1551
rect 2998 1517 3032 1551
rect 3066 1517 3100 1551
rect 3134 1517 3168 1551
rect 3202 1517 3236 1551
rect 3270 1517 3304 1551
rect 3338 1517 3372 1551
rect 3406 1517 3440 1551
rect 3474 1517 3508 1551
rect 3542 1517 3576 1551
rect 3610 1517 3644 1551
rect 3678 1517 3712 1551
rect 3746 1517 3780 1551
rect 3814 1517 3848 1551
rect 3882 1517 3916 1551
rect 3950 1517 3984 1551
rect 4018 1517 4052 1551
rect 4086 1517 4120 1551
rect 4154 1517 4188 1551
rect 4222 1517 4256 1551
rect 4290 1517 4324 1551
rect 4358 1517 4392 1551
rect 4426 1517 4460 1551
rect 4494 1517 4528 1551
rect 4562 1517 4596 1551
rect 4630 1517 4664 1551
rect 4698 1517 4732 1551
rect 4766 1517 4800 1551
rect 4834 1517 4868 1551
rect 4902 1517 4936 1551
rect 4970 1517 5004 1551
rect 5038 1517 5072 1551
rect 5106 1517 5140 1551
rect 5174 1517 5208 1551
rect 5242 1517 5276 1551
rect 5310 1517 5344 1551
rect 5378 1517 5412 1551
rect 5446 1517 5480 1551
rect 5514 1517 5548 1551
rect 5582 1517 5616 1551
rect 5650 1517 5684 1551
rect 5718 1517 5752 1551
rect 5786 1517 5820 1551
rect 5854 1517 5888 1551
rect 5922 1517 5956 1551
rect 5990 1517 6024 1551
rect 6058 1517 6092 1551
rect 6126 1517 6160 1551
rect 6194 1517 6228 1551
rect 6262 1517 6296 1551
rect 6330 1517 6364 1551
rect 6398 1517 6432 1551
rect 6466 1517 6500 1551
rect 6534 1517 6568 1551
rect 6602 1517 6636 1551
rect 6670 1517 6704 1551
rect 6738 1517 6772 1551
rect 6806 1517 6840 1551
rect 6874 1517 6908 1551
rect 6942 1517 6976 1551
rect 7010 1517 7044 1551
rect 7078 1517 7112 1551
rect 7146 1517 7180 1551
rect 7214 1517 7248 1551
rect 7282 1517 7316 1551
rect 7350 1517 7384 1551
rect 7418 1517 7452 1551
rect 7486 1517 7520 1551
rect 7554 1517 7588 1551
rect 7622 1517 7656 1551
rect 7690 1517 7724 1551
rect 7758 1517 7792 1551
rect 7826 1517 7860 1551
rect 7894 1517 7928 1551
rect 7962 1517 7996 1551
rect 8030 1517 8064 1551
rect 8098 1517 8132 1551
rect 8166 1517 8200 1551
rect 8234 1517 8268 1551
rect 8302 1517 8336 1551
rect 8370 1517 8404 1551
rect 8438 1517 8472 1551
rect 8506 1517 8540 1551
rect 8574 1517 8608 1551
rect 8642 1517 8676 1551
rect 8710 1517 8744 1551
rect 8778 1517 8812 1551
rect 8846 1517 8880 1551
rect 8914 1517 8948 1551
rect 8982 1517 9016 1551
rect 9050 1517 9084 1551
rect 9118 1517 9152 1551
rect 9186 1517 9220 1551
rect 9254 1517 9288 1551
rect 9322 1517 9356 1551
rect 9390 1517 9424 1551
rect 9458 1517 9492 1551
rect 9526 1517 9560 1551
rect 9594 1517 9628 1551
rect 9662 1517 9696 1551
rect 9730 1517 9764 1551
rect 9798 1517 9832 1551
rect 9866 1517 9900 1551
rect 9934 1517 9968 1551
rect 10002 1517 10036 1551
rect 10070 1517 10104 1551
rect 10138 1517 10172 1551
rect 10206 1517 10240 1551
rect 10274 1517 10308 1551
rect 10342 1517 10376 1551
rect 10410 1517 10444 1551
rect 10478 1517 10512 1551
rect 10546 1517 10580 1551
rect 10614 1517 10648 1551
rect 10682 1517 10716 1551
rect 10750 1517 10784 1551
rect 10818 1517 10852 1551
rect 10886 1517 10920 1551
rect 10954 1517 10988 1551
rect 11022 1517 11056 1551
rect 11090 1517 11124 1551
rect 11158 1517 11192 1551
rect 11226 1517 11260 1551
rect 11294 1517 11328 1551
rect 11362 1517 11396 1551
rect 11430 1517 11464 1551
rect 11498 1517 11532 1551
rect 11566 1517 11600 1551
rect 11634 1517 11668 1551
rect 11702 1517 11736 1551
rect 11770 1517 11804 1551
rect 11838 1517 11872 1551
rect 11906 1517 11940 1551
rect 11974 1517 12008 1551
rect 12042 1517 12076 1551
rect 12110 1517 12144 1551
rect 12178 1517 12212 1551
rect 12246 1517 12280 1551
rect 12314 1517 12348 1551
rect 12382 1517 12416 1551
rect 12450 1517 12484 1551
rect 12518 1517 12552 1551
rect 12586 1517 12620 1551
rect 12654 1517 12688 1551
rect 12722 1517 12756 1551
rect 12790 1517 12824 1551
rect 12858 1517 12892 1551
rect 12926 1517 12960 1551
rect 12994 1517 13028 1551
rect 13062 1517 13096 1551
rect 13130 1517 13164 1551
rect 13198 1517 13232 1551
rect 13266 1517 13300 1551
rect 13334 1517 13368 1551
rect 13402 1517 13436 1551
rect 13470 1517 13504 1551
rect 13538 1517 13572 1551
rect 13606 1517 13640 1551
rect 13674 1517 13708 1551
rect 13742 1517 13776 1551
rect 13810 1517 13844 1551
rect 13878 1517 13912 1551
rect 13946 1517 13980 1551
rect 14014 1517 14048 1551
rect 14082 1517 14116 1551
rect 14150 1517 14184 1551
rect 14218 1517 14252 1551
rect 14286 1517 14320 1551
rect 14354 1517 14388 1551
rect 14422 1517 14456 1551
rect 14490 1517 14524 1551
rect 14558 1517 14592 1551
rect 14626 1517 14660 1551
rect 14694 1517 14728 1551
rect 14762 1517 14796 1551
rect 14830 1517 14864 1551
rect 14898 1517 14932 1551
rect 14966 1517 15000 1551
rect 15034 1517 15068 1551
rect 15102 1517 15136 1551
rect 15170 1517 15204 1551
rect 15238 1517 15272 1551
rect 15306 1517 15340 1551
rect 15374 1517 15408 1551
rect 15442 1517 15476 1551
rect 15510 1517 15544 1551
rect 15578 1517 15612 1551
rect 15646 1517 15680 1551
rect 15714 1517 15748 1551
rect 15782 1517 15816 1551
rect 15850 1517 15884 1551
rect 15918 1517 15952 1551
rect 15986 1517 16020 1551
rect 16054 1517 16088 1551
rect 16122 1517 16156 1551
rect 16190 1517 16224 1551
rect 16258 1517 16292 1551
rect 16326 1517 16360 1551
rect 16394 1517 16428 1551
rect 16462 1517 16496 1551
rect 16530 1517 16564 1551
rect 16598 1517 16632 1551
rect 16666 1517 16700 1551
rect 16734 1517 16768 1551
rect 16802 1517 16836 1551
rect 16870 1517 16904 1551
rect 16938 1517 16972 1551
rect 17006 1517 17040 1551
rect 17074 1517 17108 1551
rect 17142 1517 17176 1551
rect 17210 1517 17244 1551
rect 17278 1517 17312 1551
rect 17346 1517 17380 1551
rect 17414 1517 17448 1551
rect 17482 1517 17516 1551
rect 17550 1517 17584 1551
rect 17618 1517 17652 1551
rect 17686 1517 17720 1551
rect 17754 1517 17788 1551
rect 17822 1517 17856 1551
rect 17890 1517 17924 1551
rect 17958 1517 17992 1551
rect 18026 1517 18060 1551
rect 18094 1517 18128 1551
rect 18162 1517 18196 1551
rect 18230 1517 18264 1551
rect 18298 1517 18332 1551
rect 18366 1517 18400 1551
rect 18434 1517 18468 1551
rect 18502 1517 18536 1551
rect 18570 1517 18604 1551
rect 18638 1517 18672 1551
rect 18706 1517 18740 1551
rect 18774 1517 18808 1551
rect 18842 1517 18876 1551
rect 18910 1517 18944 1551
rect 18978 1517 19012 1551
rect 19046 1517 19080 1551
rect 19114 1517 19148 1551
rect 19182 1517 19216 1551
rect 19250 1517 19284 1551
rect 19318 1517 19352 1551
rect 19386 1517 19420 1551
rect 19454 1517 19488 1551
rect 19522 1517 19556 1551
rect 19590 1517 19624 1551
rect 19658 1517 19692 1551
rect 19726 1517 19760 1551
rect 19794 1517 19828 1551
rect 19862 1517 19896 1551
rect 19930 1517 19964 1551
rect 19998 1517 20032 1551
rect 20066 1517 20100 1551
rect 20134 1517 20168 1551
rect 20202 1517 20236 1551
rect 20270 1517 20304 1551
rect 20338 1517 20372 1551
rect 20406 1517 20440 1551
rect 20474 1517 20508 1551
rect 20542 1517 20576 1551
rect 20610 1517 20644 1551
rect 20678 1517 20712 1551
rect 20746 1517 20780 1551
rect 20814 1517 20848 1551
rect 20882 1517 20916 1551
rect 20950 1517 20984 1551
rect 21018 1517 21052 1551
rect 21086 1517 21120 1551
rect 21154 1517 21188 1551
rect 21222 1517 21256 1551
rect 21290 1517 21324 1551
rect 21358 1517 21392 1551
rect 21426 1517 21460 1551
rect 21494 1517 21528 1551
rect 21562 1517 21596 1551
rect 21630 1517 21664 1551
rect 21698 1517 21732 1551
rect 21766 1517 21800 1551
rect 21834 1517 21868 1551
rect 21902 1517 21936 1551
rect 21970 1517 22004 1551
rect 22038 1517 22072 1551
rect 22106 1517 22140 1551
rect 22174 1517 22208 1551
rect 22242 1517 22276 1551
rect 22310 1517 22344 1551
rect 22378 1517 22412 1551
rect 22446 1517 22480 1551
rect 22514 1517 22548 1551
rect 22582 1517 22616 1551
rect 22650 1517 22684 1551
rect 22718 1517 22752 1551
rect 22786 1517 22820 1551
rect 22854 1517 22888 1551
rect 22922 1517 22956 1551
rect 22990 1517 23024 1551
rect 23058 1517 23092 1551
rect 23126 1517 23160 1551
rect 23194 1517 23228 1551
rect 23262 1517 23296 1551
rect 23330 1517 23364 1551
rect 23398 1517 23432 1551
rect 23466 1517 23500 1551
rect 23534 1517 23568 1551
rect 23602 1517 23636 1551
rect 23670 1517 23704 1551
rect 23738 1517 23772 1551
rect 23806 1517 23840 1551
rect 23874 1517 23908 1551
rect 23942 1517 23976 1551
rect 24010 1517 24044 1551
rect 24078 1517 24112 1551
rect 24146 1517 24180 1551
rect 24214 1517 24248 1551
rect 24282 1517 24316 1551
rect 24350 1517 24384 1551
rect 24418 1517 24452 1551
rect 24486 1517 24520 1551
rect 24554 1517 24588 1551
rect 24622 1517 24656 1551
rect 24690 1517 24724 1551
rect 24758 1517 24792 1551
rect 24826 1517 24860 1551
rect 24894 1517 24928 1551
rect 24962 1517 24996 1551
rect 25030 1517 25064 1551
rect 25098 1517 25132 1551
rect 25166 1517 25200 1551
rect 25234 1517 25268 1551
rect 25302 1517 25336 1551
rect 25370 1517 25404 1551
rect 25438 1517 25472 1551
rect 25506 1517 25540 1551
rect 25574 1517 25608 1551
rect 25642 1517 25676 1551
rect 25710 1517 25744 1551
rect 25778 1517 25812 1551
rect 25846 1517 25880 1551
rect 25914 1517 25948 1551
rect 25982 1517 26016 1551
rect 26050 1517 26084 1551
rect 26118 1517 26152 1551
rect 26186 1517 26220 1551
rect 26254 1517 26288 1551
rect 26322 1517 26356 1551
rect 26390 1517 26424 1551
rect 26458 1517 26492 1551
rect 26526 1517 26560 1551
rect 26594 1517 26628 1551
rect 26662 1517 26696 1551
rect 26730 1517 26764 1551
rect 26798 1517 26832 1551
rect 26866 1517 26900 1551
rect 26934 1517 26968 1551
rect 27002 1517 27036 1551
rect 27070 1517 27104 1551
rect 27138 1517 27172 1551
rect 27206 1517 27240 1551
rect 27274 1517 27308 1551
rect 27342 1517 27376 1551
rect 27410 1517 27444 1551
rect 27478 1517 27508 1551
rect 1979 1487 27508 1517
rect 1975 1472 27508 1487
rect 1795 1415 1801 1449
rect 1975 1448 2010 1472
rect 2044 1448 2079 1472
rect 2113 1448 2148 1472
rect 1795 1376 1805 1415
rect 1907 1404 1945 1438
rect 27546 1404 27580 1414
rect 1907 1376 1942 1404
rect 1795 1342 1801 1376
rect 1835 1342 1873 1370
rect 1795 1270 1873 1342
rect 27686 1342 27692 7784
rect 27395 1270 27434 1302
rect 27468 1270 27507 1302
rect 27541 1270 27580 1302
rect 27614 1270 27692 1342
rect 1795 1264 27692 1270
rect 27905 8841 27911 8875
rect 28089 8841 28095 8875
rect 27905 8796 27915 8841
rect 28085 8796 28095 8841
rect 27905 8762 27911 8796
rect 28089 8762 28095 8796
rect 27905 8717 27915 8762
rect 28085 8717 28095 8762
rect 27905 8683 27911 8717
rect 28089 8683 28095 8717
rect 27905 8638 27915 8683
rect 28085 8638 28095 8683
rect 27905 8604 27911 8638
rect 28089 8604 28095 8638
rect 27905 8528 27915 8604
rect 28085 8528 28095 8604
rect 27905 8494 27911 8528
rect 28089 8494 28095 8528
rect 27905 8455 27915 8494
rect 28085 8455 28095 8494
rect 27905 8421 27911 8455
rect 28089 8421 28095 8455
rect 27905 8382 27915 8421
rect 28085 8382 28095 8421
rect 27905 8348 27911 8382
rect 28089 8348 28095 8382
rect 27905 8309 27915 8348
rect 28085 8309 28095 8348
rect 27905 8275 27911 8309
rect 28089 8275 28095 8309
rect 27905 8236 27915 8275
rect 28085 8236 28095 8275
rect 1347 1189 1353 1223
rect 1527 1222 1537 1261
rect 1347 1150 1357 1189
rect 1531 1188 1537 1222
rect 1347 1116 1353 1150
rect 1527 1149 1537 1188
rect 1347 1077 1357 1116
rect 1531 1115 1537 1149
rect 1527 1082 1537 1115
rect 27905 1082 27911 8236
rect 1347 1043 1353 1077
rect 1527 1076 27911 1082
rect 1347 1004 1357 1043
rect 1347 970 1353 1004
rect 23779 1042 23818 1076
rect 23852 1042 23891 1076
rect 23925 1042 23964 1076
rect 23998 1042 24037 1076
rect 24071 1042 24110 1076
rect 24144 1042 24183 1076
rect 24217 1042 24256 1076
rect 24290 1042 24329 1076
rect 24363 1042 24402 1076
rect 24436 1042 24475 1076
rect 24509 1042 24548 1076
rect 24582 1042 24621 1076
rect 24655 1042 24694 1076
rect 24728 1042 24767 1076
rect 24801 1042 24840 1076
rect 24874 1042 24913 1076
rect 24947 1042 24986 1076
rect 25020 1042 25059 1076
rect 25093 1042 25132 1076
rect 25166 1042 25205 1076
rect 25239 1042 25278 1076
rect 25312 1042 25351 1076
rect 25385 1042 25424 1076
rect 25458 1042 25497 1076
rect 25531 1042 25570 1076
rect 25604 1042 25643 1076
rect 25677 1042 25716 1076
rect 25750 1042 25789 1076
rect 25823 1042 25862 1076
rect 25896 1042 25935 1076
rect 25969 1042 26008 1076
rect 26042 1042 26081 1076
rect 26115 1042 26154 1076
rect 26188 1042 26227 1076
rect 26261 1042 26300 1076
rect 26334 1042 26373 1076
rect 26407 1042 26446 1076
rect 26480 1042 26519 1076
rect 26553 1042 26592 1076
rect 26626 1042 26665 1076
rect 26699 1042 26738 1076
rect 26772 1042 26811 1076
rect 26845 1042 26884 1076
rect 26918 1042 26957 1076
rect 26991 1042 27030 1076
rect 27064 1042 27103 1076
rect 27137 1042 27176 1076
rect 27210 1042 27249 1076
rect 27283 1042 27322 1076
rect 27356 1042 27395 1076
rect 27429 1042 27468 1076
rect 27502 1042 27541 1076
rect 27575 1042 27614 1076
rect 27648 1042 27687 1076
rect 27721 1042 27760 1076
rect 27794 1042 27833 1076
rect 27867 1042 27911 1076
rect 23779 1004 27911 1042
rect 23779 978 23818 1004
rect 23852 978 23891 1004
rect 23925 978 23964 1004
rect 23998 978 24037 1004
rect 24071 978 24110 1004
rect 24144 978 24183 1004
rect 24217 978 24256 1004
rect 24290 978 24329 1004
rect 24363 978 24402 1004
rect 24436 978 24475 1004
rect 24509 978 24548 1004
rect 24582 978 24621 1004
rect 24655 978 24694 1004
rect 24728 978 24767 1004
rect 24801 978 24840 1004
rect 24874 978 24913 1004
rect 24947 978 24986 1004
rect 25020 978 25059 1004
rect 25093 978 25132 1004
rect 25166 978 25205 1004
rect 25239 978 25278 1004
rect 25312 978 25351 1004
rect 25385 978 25424 1004
rect 25458 978 25497 1004
rect 25531 978 25570 1004
rect 25604 978 25643 1004
rect 25677 978 25716 1004
rect 25750 978 25789 1004
rect 25823 978 25862 1004
rect 25896 978 25935 1004
rect 25969 978 26008 1004
rect 26042 978 26081 1004
rect 26115 978 26154 1004
rect 26188 978 26227 1004
rect 26261 978 26300 1004
rect 26334 978 26373 1004
rect 26407 978 26446 1004
rect 26480 978 26519 1004
rect 26553 978 26592 1004
rect 26626 978 26665 1004
rect 26699 978 26738 1004
rect 26772 978 26811 1004
rect 26845 978 26884 1004
rect 26918 978 26957 1004
rect 26991 978 27030 1004
rect 27064 978 27103 1004
rect 27137 978 27176 1004
rect 27210 978 27249 1004
rect 27283 978 27322 1004
rect 27356 978 27395 1004
rect 27429 978 27468 1004
rect 27502 978 27541 1004
rect 27575 978 27614 1004
rect 27648 978 27687 1004
rect 27721 978 27760 1004
rect 27794 978 27833 1004
rect 27867 978 27911 1004
rect 1347 892 1357 970
rect 28089 930 28095 8236
rect 1357 876 1561 882
rect 1595 876 1630 898
rect 1664 876 1699 898
rect 1733 876 1768 898
rect 1802 876 1837 898
rect 1871 876 1906 898
rect 1940 876 1975 898
rect 2009 876 2044 898
rect 2078 876 2113 898
rect 2147 876 2182 898
rect 2216 876 2251 898
rect 2285 876 2320 898
rect 2354 876 2389 898
rect 2423 876 2458 898
rect 2492 876 2527 898
rect 2561 876 2596 898
rect 2630 876 2665 898
rect 2699 876 2734 898
rect 2768 876 2803 898
rect 2837 876 2872 898
rect 2906 876 2941 898
rect 2975 876 3010 898
rect 3044 876 3079 898
rect 3113 876 3148 898
rect 3182 876 3217 898
rect 3251 876 3286 898
rect 3320 876 3355 898
rect 3389 876 3424 898
rect 3458 876 3493 898
rect 3527 876 3562 898
rect 3596 876 3631 898
rect 3665 876 3700 898
rect 3734 876 3769 898
rect 3803 876 3838 898
rect 3872 876 3907 898
rect 3941 876 3976 898
rect 4010 876 4045 898
rect 4079 876 4114 898
rect 4148 876 4183 898
rect 1357 842 4183 876
rect 28085 892 28095 930
rect 1357 808 1561 842
rect 1595 808 1630 842
rect 1664 808 1699 842
rect 1733 808 1768 842
rect 1802 808 1837 842
rect 1871 808 1906 842
rect 1940 808 1975 842
rect 2009 808 2044 842
rect 2078 808 2113 842
rect 2147 808 2182 842
rect 2216 808 2251 842
rect 2285 808 2320 842
rect 2354 808 2389 842
rect 2423 808 2458 842
rect 2492 808 2527 842
rect 2561 808 2596 842
rect 2630 808 2665 842
rect 2699 808 2734 842
rect 2768 808 2803 842
rect 2837 808 2872 842
rect 2906 808 2941 842
rect 2975 808 3010 842
rect 3044 808 3079 842
rect 3113 808 3148 842
rect 3182 808 3217 842
rect 3251 808 3286 842
rect 3320 808 3355 842
rect 3389 808 3424 842
rect 3458 808 3493 842
rect 3527 808 3562 842
rect 3596 808 3631 842
rect 3665 808 3700 842
rect 3734 808 3769 842
rect 3803 808 3838 842
rect 3872 808 3907 842
rect 3941 808 3976 842
rect 4010 808 4045 842
rect 4079 808 4114 842
rect 4148 808 4183 842
rect 27881 808 28085 842
rect 144 -1453 548 -1441
rect 144 -1487 165 -1453
rect 199 -1487 253 -1453
rect 287 -1487 340 -1453
rect 374 -1487 427 -1453
rect 461 -1487 514 -1453
rect 144 -1539 548 -1487
rect 144 -1573 165 -1539
rect 199 -1573 253 -1539
rect 287 -1573 340 -1539
rect 374 -1573 427 -1539
rect 461 -1573 514 -1539
rect 144 -1577 548 -1573
<< viali >>
rect 1425 9212 1459 9226
rect 1425 9192 1459 9212
rect 1498 9192 1532 9226
rect 1571 9192 1605 9226
rect 1644 9192 1678 9226
rect 1717 9192 1751 9226
rect 1790 9192 1824 9226
rect 1863 9192 1897 9226
rect 1936 9192 1970 9226
rect 2009 9192 2043 9226
rect 2082 9192 2116 9226
rect 2155 9192 2189 9226
rect 2228 9192 2262 9226
rect 2301 9192 2335 9226
rect 2374 9192 2408 9226
rect 2447 9192 2481 9226
rect 2520 9192 2554 9226
rect 2593 9192 2627 9226
rect 2666 9192 2700 9226
rect 2739 9192 2773 9226
rect 2812 9192 2846 9226
rect 2885 9192 2919 9226
rect 2958 9192 2992 9226
rect 3031 9192 3065 9226
rect 3104 9192 3138 9226
rect 3177 9192 3211 9226
rect 3250 9192 3284 9226
rect 3323 9192 3357 9226
rect 3396 9192 3430 9226
rect 3469 9192 3503 9226
rect 3542 9192 3576 9226
rect 3615 9192 3649 9226
rect 3688 9192 3722 9226
rect 3761 9192 3795 9226
rect 3834 9192 3868 9226
rect 3907 9192 3941 9226
rect 3980 9192 4014 9226
rect 4053 9192 4087 9226
rect 4126 9192 4160 9226
rect 4199 9192 4233 9226
rect 4272 9192 4306 9226
rect 4345 9192 4379 9226
rect 4418 9192 4452 9226
rect 4491 9192 4525 9226
rect 4564 9192 4598 9226
rect 4637 9192 4671 9226
rect 4710 9192 4744 9226
rect 4783 9192 4817 9226
rect 4856 9192 4890 9226
rect 4929 9192 4963 9226
rect 5002 9192 5036 9226
rect 5075 9192 5109 9226
rect 5148 9192 5182 9226
rect 5221 9192 5255 9226
rect 5294 9192 5328 9226
rect 5367 9192 5401 9226
rect 5440 9192 5474 9226
rect 1353 1992 1357 9154
rect 1357 9082 1459 9154
rect 1498 9144 1532 9154
rect 1498 9120 1527 9144
rect 1527 9120 1532 9144
rect 1571 9120 1605 9154
rect 1644 9120 1678 9154
rect 1717 9120 1751 9154
rect 1790 9120 1824 9154
rect 1863 9120 1897 9154
rect 1936 9120 1970 9154
rect 2009 9120 2043 9154
rect 2082 9120 2116 9154
rect 2155 9120 2189 9154
rect 2228 9120 2262 9154
rect 2301 9120 2335 9154
rect 2374 9120 2408 9154
rect 2447 9120 2481 9154
rect 2520 9120 2554 9154
rect 2593 9120 2627 9154
rect 2666 9120 2700 9154
rect 2739 9120 2773 9154
rect 2812 9120 2846 9154
rect 2885 9120 2919 9154
rect 2958 9120 2992 9154
rect 3031 9120 3065 9154
rect 3104 9120 3138 9154
rect 3177 9120 3211 9154
rect 3250 9120 3284 9154
rect 3323 9120 3357 9154
rect 3396 9120 3430 9154
rect 3469 9120 3503 9154
rect 3542 9120 3576 9154
rect 3615 9120 3649 9154
rect 3688 9120 3722 9154
rect 3761 9120 3795 9154
rect 3834 9120 3868 9154
rect 3907 9120 3941 9154
rect 3980 9120 4014 9154
rect 4053 9120 4087 9154
rect 4126 9120 4160 9154
rect 4199 9120 4233 9154
rect 4272 9120 4306 9154
rect 4345 9120 4379 9154
rect 4418 9120 4452 9154
rect 4491 9120 4525 9154
rect 4564 9120 4598 9154
rect 4637 9120 4671 9154
rect 4710 9120 4744 9154
rect 4783 9120 4817 9154
rect 4856 9120 4890 9154
rect 4929 9120 4963 9154
rect 5002 9120 5036 9154
rect 5075 9120 5109 9154
rect 5148 9120 5182 9154
rect 5221 9120 5255 9154
rect 5294 9120 5328 9154
rect 5367 9120 5401 9154
rect 5440 9120 5474 9154
rect 5513 9120 27867 9226
rect 27911 9160 27945 9194
rect 27983 9160 28017 9194
rect 28055 9160 28089 9194
rect 5585 9110 27867 9120
rect 27911 9110 27945 9114
rect 1357 2064 1527 9082
rect 1527 2064 1531 9082
rect 1570 9048 1604 9082
rect 1643 9048 1677 9082
rect 1716 9048 1750 9082
rect 1789 9048 1823 9082
rect 1862 9048 1896 9082
rect 1935 9048 1969 9082
rect 2008 9048 2042 9082
rect 2081 9048 2115 9082
rect 2154 9048 2188 9082
rect 2227 9048 2261 9082
rect 2300 9048 2334 9082
rect 2373 9048 2407 9082
rect 2446 9048 2480 9082
rect 2519 9048 2553 9082
rect 2592 9048 2626 9082
rect 2665 9048 2699 9082
rect 2738 9048 2772 9082
rect 2811 9048 2845 9082
rect 2884 9048 2918 9082
rect 2957 9048 2991 9082
rect 3030 9048 3064 9082
rect 3103 9048 3137 9082
rect 3176 9048 3210 9082
rect 3249 9048 3283 9082
rect 3322 9048 3356 9082
rect 3395 9048 3429 9082
rect 3468 9048 3502 9082
rect 3541 9048 3575 9082
rect 3614 9048 3648 9082
rect 3687 9048 3721 9082
rect 3760 9048 3794 9082
rect 3833 9048 3867 9082
rect 3906 9048 3940 9082
rect 3979 9048 4013 9082
rect 4052 9048 4086 9082
rect 4125 9048 4159 9082
rect 4198 9048 4232 9082
rect 4271 9048 4305 9082
rect 4344 9048 4378 9082
rect 4417 9048 4451 9082
rect 4490 9048 4524 9082
rect 4563 9048 4597 9082
rect 4636 9048 4670 9082
rect 4709 9048 4743 9082
rect 4782 9048 4816 9082
rect 4855 9048 4889 9082
rect 4928 9048 4962 9082
rect 5001 9048 5035 9082
rect 5074 9048 5108 9082
rect 5147 9048 5181 9082
rect 5220 9048 5254 9082
rect 5293 9048 5327 9082
rect 5366 9048 5400 9082
rect 5439 9048 5473 9082
rect 5512 9048 5546 9082
rect 5585 9048 27867 9110
rect 27911 9080 27945 9110
rect 27983 9080 28017 9114
rect 28055 9080 28089 9114
rect 27911 9000 27915 9034
rect 27915 9000 27945 9034
rect 27983 9000 28017 9034
rect 28055 9000 28085 9034
rect 28085 9000 28089 9034
rect 27911 8920 27915 8954
rect 27915 8920 27945 8954
rect 27983 8920 28017 8954
rect 28055 8920 28085 8954
rect 28085 8920 28089 8954
rect 1357 1992 1459 2064
rect 1497 1991 1527 2025
rect 1527 1991 1531 2025
rect 1353 1919 1357 1953
rect 1357 1919 1387 1953
rect 1425 1919 1459 1953
rect 1497 1918 1527 1952
rect 1527 1918 1531 1952
rect 1353 1846 1357 1880
rect 1357 1846 1387 1880
rect 1425 1846 1459 1880
rect 1497 1845 1527 1879
rect 1527 1845 1531 1879
rect 1353 1773 1357 1807
rect 1357 1773 1387 1807
rect 1425 1773 1459 1807
rect 1497 1772 1527 1806
rect 1527 1772 1531 1806
rect 1353 1700 1357 1734
rect 1357 1700 1387 1734
rect 1425 1700 1459 1734
rect 1497 1699 1527 1733
rect 1527 1699 1531 1733
rect 1353 1627 1357 1661
rect 1357 1627 1387 1661
rect 1425 1627 1459 1661
rect 1497 1626 1527 1660
rect 1527 1626 1531 1660
rect 1353 1554 1357 1588
rect 1357 1554 1387 1588
rect 1425 1554 1459 1588
rect 1497 1553 1527 1587
rect 1527 1553 1531 1587
rect 1353 1481 1357 1515
rect 1357 1481 1387 1515
rect 1425 1481 1459 1515
rect 1497 1480 1527 1514
rect 1527 1480 1531 1514
rect 1353 1408 1357 1442
rect 1357 1408 1387 1442
rect 1425 1408 1459 1442
rect 1497 1407 1527 1441
rect 1527 1407 1531 1441
rect 1353 1335 1357 1369
rect 1357 1335 1387 1369
rect 1425 1335 1459 1369
rect 1497 1334 1527 1368
rect 1527 1334 1531 1368
rect 1353 1262 1357 1296
rect 1357 1262 1387 1296
rect 1425 1262 1459 1296
rect 1497 1261 1527 1295
rect 1527 1261 1531 1295
rect 1873 8843 1907 8847
rect 1946 8843 1980 8847
rect 2019 8843 2053 8847
rect 2092 8843 27614 8847
rect 1873 8813 1907 8843
rect 1946 8813 1980 8843
rect 2019 8813 2053 8843
rect 1801 8741 1805 8775
rect 1805 8741 1839 8775
rect 1839 8741 1873 8775
rect 1873 8741 1907 8775
rect 1946 8741 1980 8775
rect 2019 8741 2053 8775
rect 2092 8741 27407 8843
rect 27407 8809 27442 8843
rect 27442 8809 27476 8843
rect 27476 8809 27511 8843
rect 27511 8809 27545 8843
rect 27545 8809 27580 8843
rect 27580 8809 27614 8843
rect 27407 8775 27614 8809
rect 27407 8741 27442 8775
rect 27442 8741 27476 8775
rect 27476 8741 27511 8775
rect 27511 8741 27545 8775
rect 27545 8741 27580 8775
rect 27580 8741 27614 8775
rect 27652 8741 27682 8775
rect 27682 8741 27686 8775
rect 1801 8706 1907 8741
rect 1801 8672 1805 8706
rect 1805 8672 1839 8706
rect 1839 8672 1873 8706
rect 1873 8672 1907 8706
rect 1907 8673 1941 8703
rect 1941 8673 1979 8703
rect 2018 8673 2052 8703
rect 2091 8673 2125 8703
rect 2164 8673 27339 8741
rect 27339 8707 27542 8741
rect 27339 8673 27374 8707
rect 27374 8673 27408 8707
rect 27408 8673 27443 8707
rect 27443 8673 27477 8707
rect 27477 8673 27512 8707
rect 1907 8672 1979 8673
rect 1801 8638 1979 8672
rect 2018 8669 2052 8673
rect 2091 8669 2125 8673
rect 2164 8669 27512 8673
rect 27512 8669 27542 8707
rect 27580 8667 27614 8701
rect 27652 8667 27682 8701
rect 27682 8667 27686 8701
rect 1801 8637 1941 8638
rect 1801 8603 1805 8637
rect 1805 8603 1839 8637
rect 1839 8603 1873 8637
rect 1873 8603 1907 8637
rect 1907 8604 1941 8637
rect 1941 8604 1975 8638
rect 1975 8604 1979 8638
rect 1907 8603 1979 8604
rect 1801 8569 1979 8603
rect 1801 8568 1941 8569
rect 1801 8534 1805 8568
rect 1805 8534 1839 8568
rect 1839 8534 1873 8568
rect 1873 8534 1907 8568
rect 1907 8535 1941 8568
rect 1941 8535 1975 8569
rect 1975 8535 1979 8569
rect 1907 8534 1979 8535
rect 1801 8500 1979 8534
rect 1801 8499 1941 8500
rect 1801 8465 1805 8499
rect 1805 8465 1839 8499
rect 1839 8465 1873 8499
rect 1873 8465 1907 8499
rect 1907 8466 1941 8499
rect 1941 8466 1975 8500
rect 1975 8466 1979 8500
rect 1907 8465 1979 8466
rect 1801 8431 1979 8465
rect 1801 8430 1941 8431
rect 1801 8396 1805 8430
rect 1805 8396 1839 8430
rect 1839 8396 1873 8430
rect 1873 8396 1907 8430
rect 1907 8397 1941 8430
rect 1941 8397 1975 8431
rect 1975 8397 1979 8431
rect 1907 8396 1979 8397
rect 1801 8362 1979 8396
rect 1801 8361 1941 8362
rect 1801 8327 1805 8361
rect 1805 8327 1839 8361
rect 1839 8327 1873 8361
rect 1873 8327 1907 8361
rect 1907 8328 1941 8361
rect 1941 8328 1975 8362
rect 1975 8328 1979 8362
rect 1907 8327 1979 8328
rect 1801 8293 1979 8327
rect 1801 8292 1941 8293
rect 1801 8258 1805 8292
rect 1805 8258 1839 8292
rect 1839 8258 1873 8292
rect 1873 8258 1907 8292
rect 1907 8259 1941 8292
rect 1941 8259 1975 8293
rect 1975 8259 1979 8293
rect 1907 8258 1979 8259
rect 1801 8224 1979 8258
rect 1801 8223 1941 8224
rect 1801 8189 1805 8223
rect 1805 8189 1839 8223
rect 1839 8189 1873 8223
rect 1873 8189 1907 8223
rect 1907 8190 1941 8223
rect 1941 8190 1975 8224
rect 1975 8190 1979 8224
rect 1907 8189 1979 8190
rect 1801 8155 1979 8189
rect 1801 8154 1941 8155
rect 1801 8120 1805 8154
rect 1805 8120 1839 8154
rect 1839 8120 1873 8154
rect 1873 8120 1907 8154
rect 1907 8121 1941 8154
rect 1941 8121 1975 8155
rect 1975 8121 1979 8155
rect 1907 8120 1979 8121
rect 1801 8086 1979 8120
rect 1801 8085 1941 8086
rect 1801 8051 1805 8085
rect 1805 8051 1839 8085
rect 1839 8051 1873 8085
rect 1873 8051 1907 8085
rect 1907 8052 1941 8085
rect 1941 8052 1975 8086
rect 1975 8052 1979 8086
rect 1907 8051 1979 8052
rect 1801 8017 1979 8051
rect 1801 8016 1941 8017
rect 1801 7982 1805 8016
rect 1805 7982 1839 8016
rect 1839 7982 1873 8016
rect 1873 7982 1907 8016
rect 1907 7983 1941 8016
rect 1941 7983 1975 8017
rect 1975 7983 1979 8017
rect 1907 7982 1979 7983
rect 1801 7948 1979 7982
rect 1801 7947 1941 7948
rect 1801 7913 1805 7947
rect 1805 7913 1839 7947
rect 1839 7913 1873 7947
rect 1873 7913 1907 7947
rect 1907 7914 1941 7947
rect 1941 7914 1975 7948
rect 1975 7914 1979 7948
rect 1907 7913 1979 7914
rect 1801 7879 1979 7913
rect 1801 7878 1941 7879
rect 1801 7844 1805 7878
rect 1805 7844 1839 7878
rect 1839 7844 1873 7878
rect 1873 7844 1907 7878
rect 1907 7845 1941 7878
rect 1941 7845 1975 7879
rect 1975 7845 1979 7879
rect 1907 7844 1979 7845
rect 1801 7810 1979 7844
rect 1801 7809 1941 7810
rect 1801 7775 1805 7809
rect 1805 7775 1839 7809
rect 1839 7775 1873 7809
rect 1873 7775 1907 7809
rect 1907 7776 1941 7809
rect 1941 7776 1975 7810
rect 1975 7776 1979 7810
rect 1907 7775 1979 7776
rect 1801 7741 1979 7775
rect 1801 7740 1941 7741
rect 1801 7706 1805 7740
rect 1805 7706 1839 7740
rect 1839 7706 1873 7740
rect 1873 7706 1907 7740
rect 1907 7707 1941 7740
rect 1941 7707 1975 7741
rect 1975 7707 1979 7741
rect 1907 7706 1979 7707
rect 1801 7672 1979 7706
rect 1801 7671 1941 7672
rect 1801 7637 1805 7671
rect 1805 7637 1839 7671
rect 1839 7637 1873 7671
rect 1873 7637 1907 7671
rect 1907 7638 1941 7671
rect 1941 7638 1975 7672
rect 1975 7638 1979 7672
rect 1907 7637 1979 7638
rect 1801 7603 1979 7637
rect 1801 7602 1941 7603
rect 1801 7568 1805 7602
rect 1805 7568 1839 7602
rect 1839 7568 1873 7602
rect 1873 7568 1907 7602
rect 1907 7569 1941 7602
rect 1941 7569 1975 7603
rect 1975 7569 1979 7603
rect 1907 7568 1979 7569
rect 1801 7534 1979 7568
rect 1801 7533 1941 7534
rect 1801 7499 1805 7533
rect 1805 7499 1839 7533
rect 1839 7499 1873 7533
rect 1873 7499 1907 7533
rect 1907 7500 1941 7533
rect 1941 7500 1975 7534
rect 1975 7500 1979 7534
rect 1907 7499 1979 7500
rect 1801 7465 1979 7499
rect 1801 7464 1941 7465
rect 1801 7430 1805 7464
rect 1805 7430 1839 7464
rect 1839 7430 1873 7464
rect 1873 7430 1907 7464
rect 1907 7431 1941 7464
rect 1941 7431 1975 7465
rect 1975 7431 1979 7465
rect 1907 7430 1979 7431
rect 1801 7396 1979 7430
rect 1801 7395 1941 7396
rect 1801 7361 1805 7395
rect 1805 7361 1839 7395
rect 1839 7361 1873 7395
rect 1873 7361 1907 7395
rect 1907 7362 1941 7395
rect 1941 7362 1975 7396
rect 1975 7362 1979 7396
rect 1907 7361 1979 7362
rect 1801 7327 1979 7361
rect 1801 7326 1941 7327
rect 1801 7292 1805 7326
rect 1805 7292 1839 7326
rect 1839 7292 1873 7326
rect 1873 7292 1907 7326
rect 1907 7293 1941 7326
rect 1941 7293 1975 7327
rect 1975 7293 1979 7327
rect 1907 7292 1979 7293
rect 1801 7258 1979 7292
rect 1801 7257 1941 7258
rect 1801 7223 1805 7257
rect 1805 7223 1839 7257
rect 1839 7223 1873 7257
rect 1873 7223 1907 7257
rect 1907 7224 1941 7257
rect 1941 7224 1975 7258
rect 1975 7224 1979 7258
rect 1907 7223 1979 7224
rect 1801 7189 1979 7223
rect 1801 7188 1941 7189
rect 1801 7154 1805 7188
rect 1805 7154 1839 7188
rect 1839 7154 1873 7188
rect 1873 7154 1907 7188
rect 1907 7155 1941 7188
rect 1941 7155 1975 7189
rect 1975 7155 1979 7189
rect 1907 7154 1979 7155
rect 1801 7120 1979 7154
rect 1801 7119 1941 7120
rect 1801 7085 1805 7119
rect 1805 7085 1839 7119
rect 1839 7085 1873 7119
rect 1873 7085 1907 7119
rect 1907 7086 1941 7119
rect 1941 7086 1975 7120
rect 1975 7086 1979 7120
rect 1907 7085 1979 7086
rect 1801 7051 1979 7085
rect 1801 7050 1941 7051
rect 1801 7016 1805 7050
rect 1805 7016 1839 7050
rect 1839 7016 1873 7050
rect 1873 7016 1907 7050
rect 1907 7017 1941 7050
rect 1941 7017 1975 7051
rect 1975 7017 1979 7051
rect 1907 7016 1979 7017
rect 1801 6982 1979 7016
rect 1801 6981 1941 6982
rect 1801 6947 1805 6981
rect 1805 6947 1839 6981
rect 1839 6947 1873 6981
rect 1873 6947 1907 6981
rect 1907 6948 1941 6981
rect 1941 6948 1975 6982
rect 1975 6948 1979 6982
rect 1907 6947 1979 6948
rect 1801 6913 1979 6947
rect 1801 6912 1941 6913
rect 1801 6878 1805 6912
rect 1805 6878 1839 6912
rect 1839 6878 1873 6912
rect 1873 6878 1907 6912
rect 1907 6879 1941 6912
rect 1941 6879 1975 6913
rect 1975 6879 1979 6913
rect 1907 6878 1979 6879
rect 1801 6844 1979 6878
rect 1801 6843 1941 6844
rect 1801 6809 1805 6843
rect 1805 6809 1839 6843
rect 1839 6809 1873 6843
rect 1873 6809 1907 6843
rect 1907 6810 1941 6843
rect 1941 6810 1975 6844
rect 1975 6810 1979 6844
rect 1907 6809 1979 6810
rect 1801 6775 1979 6809
rect 1801 6774 1941 6775
rect 1801 6740 1805 6774
rect 1805 6740 1839 6774
rect 1839 6740 1873 6774
rect 1873 6740 1907 6774
rect 1907 6741 1941 6774
rect 1941 6741 1975 6775
rect 1975 6741 1979 6775
rect 1907 6740 1979 6741
rect 1801 6706 1979 6740
rect 1801 6705 1941 6706
rect 1801 6671 1805 6705
rect 1805 6671 1839 6705
rect 1839 6671 1873 6705
rect 1873 6671 1907 6705
rect 1907 6672 1941 6705
rect 1941 6672 1975 6706
rect 1975 6672 1979 6706
rect 1907 6671 1979 6672
rect 1801 6637 1979 6671
rect 1801 6636 1941 6637
rect 1801 6602 1805 6636
rect 1805 6602 1839 6636
rect 1839 6602 1873 6636
rect 1873 6602 1907 6636
rect 1907 6603 1941 6636
rect 1941 6603 1975 6637
rect 1975 6603 1979 6637
rect 1907 6602 1979 6603
rect 1801 6568 1979 6602
rect 1801 6567 1941 6568
rect 1801 6533 1805 6567
rect 1805 6533 1839 6567
rect 1839 6533 1873 6567
rect 1873 6533 1907 6567
rect 1907 6534 1941 6567
rect 1941 6534 1975 6568
rect 1975 6534 1979 6568
rect 1907 6533 1979 6534
rect 1801 6499 1979 6533
rect 1801 6498 1941 6499
rect 1801 6464 1805 6498
rect 1805 6464 1839 6498
rect 1839 6464 1873 6498
rect 1873 6464 1907 6498
rect 1907 6465 1941 6498
rect 1941 6465 1975 6499
rect 1975 6465 1979 6499
rect 1907 6464 1979 6465
rect 1801 6430 1979 6464
rect 1801 6429 1941 6430
rect 1801 6395 1805 6429
rect 1805 6395 1839 6429
rect 1839 6395 1873 6429
rect 1873 6395 1907 6429
rect 1907 6396 1941 6429
rect 1941 6396 1975 6430
rect 1975 6396 1979 6430
rect 1907 6395 1979 6396
rect 1801 6361 1979 6395
rect 1801 6360 1941 6361
rect 1801 6326 1805 6360
rect 1805 6326 1839 6360
rect 1839 6326 1873 6360
rect 1873 6326 1907 6360
rect 1907 6327 1941 6360
rect 1941 6327 1975 6361
rect 1975 6327 1979 6361
rect 1907 6326 1979 6327
rect 1801 6292 1979 6326
rect 1801 6291 1941 6292
rect 1801 6257 1805 6291
rect 1805 6257 1839 6291
rect 1839 6257 1873 6291
rect 1873 6257 1907 6291
rect 1907 6258 1941 6291
rect 1941 6258 1975 6292
rect 1975 6258 1979 6292
rect 1907 6257 1979 6258
rect 1801 6223 1979 6257
rect 1801 6222 1941 6223
rect 1801 6188 1805 6222
rect 1805 6188 1839 6222
rect 1839 6188 1873 6222
rect 1873 6188 1907 6222
rect 1907 6189 1941 6222
rect 1941 6189 1975 6223
rect 1975 6189 1979 6223
rect 1907 6188 1979 6189
rect 1801 6154 1979 6188
rect 1801 6153 1941 6154
rect 1801 6119 1805 6153
rect 1805 6119 1839 6153
rect 1839 6119 1873 6153
rect 1873 6119 1907 6153
rect 1907 6120 1941 6153
rect 1941 6120 1975 6154
rect 1975 6120 1979 6154
rect 1907 6119 1979 6120
rect 1801 6085 1979 6119
rect 1801 6084 1941 6085
rect 1801 6050 1805 6084
rect 1805 6050 1839 6084
rect 1839 6050 1873 6084
rect 1873 6050 1907 6084
rect 1907 6051 1941 6084
rect 1941 6051 1975 6085
rect 1975 6051 1979 6085
rect 1907 6050 1979 6051
rect 1801 6016 1979 6050
rect 1801 6015 1941 6016
rect 1801 5437 1805 6015
rect 1805 5947 1907 6015
rect 1907 5982 1941 6015
rect 1941 5982 1975 6016
rect 1975 5982 1979 6016
rect 1907 5947 1979 5982
rect 1805 5437 1975 5947
rect 1975 5437 1979 5947
rect 1801 5429 1979 5437
rect 27508 8595 27512 8629
rect 27512 8595 27542 8629
rect 27580 8593 27614 8627
rect 27652 8593 27682 8627
rect 27682 8593 27686 8627
rect 27508 8521 27512 8555
rect 27512 8521 27542 8555
rect 27580 8519 27614 8553
rect 27652 8519 27682 8553
rect 27682 8519 27686 8553
rect 1801 5369 1907 5429
rect 1945 5369 1979 5390
rect 1801 5357 1805 5369
rect 1805 5357 1839 5369
rect 1839 5357 1873 5369
rect 1873 5357 1907 5369
rect 1945 5356 1975 5369
rect 1975 5356 1979 5369
rect 1801 5300 1835 5318
rect 1873 5300 1907 5318
rect 1945 5300 1979 5317
rect 1801 5284 1805 5300
rect 1805 5284 1835 5300
rect 1873 5284 1907 5300
rect 1945 5283 1975 5300
rect 1975 5283 1979 5300
rect 1801 5231 1835 5245
rect 1873 5231 1907 5245
rect 1945 5231 1979 5244
rect 1801 5211 1805 5231
rect 1805 5211 1835 5231
rect 1873 5211 1907 5231
rect 1945 5210 1975 5231
rect 1975 5210 1979 5231
rect 1801 5162 1835 5172
rect 1873 5162 1907 5172
rect 1945 5162 1979 5171
rect 1801 5138 1805 5162
rect 1805 5138 1835 5162
rect 1873 5138 1907 5162
rect 1945 5137 1975 5162
rect 1975 5137 1979 5162
rect 1801 5093 1835 5099
rect 1873 5093 1907 5099
rect 1945 5093 1979 5098
rect 1801 5065 1805 5093
rect 1805 5065 1835 5093
rect 1873 5065 1907 5093
rect 1945 5064 1975 5093
rect 1975 5064 1979 5093
rect 1801 5024 1835 5026
rect 1873 5024 1907 5026
rect 1945 5024 1979 5025
rect 1801 4992 1805 5024
rect 1805 4992 1835 5024
rect 1873 4992 1907 5024
rect 1945 4991 1975 5024
rect 1975 4991 1979 5024
rect 1801 4921 1805 4953
rect 1805 4921 1835 4953
rect 1873 4921 1907 4953
rect 1945 4921 1975 4952
rect 1975 4921 1979 4952
rect 1801 4919 1835 4921
rect 1873 4919 1907 4921
rect 1945 4918 1979 4921
rect 1801 4852 1805 4880
rect 1805 4852 1835 4880
rect 1873 4852 1907 4880
rect 1945 4852 1975 4879
rect 1975 4852 1979 4879
rect 1801 4846 1835 4852
rect 1873 4846 1907 4852
rect 1945 4845 1979 4852
rect 1801 4783 1805 4807
rect 1805 4783 1835 4807
rect 1873 4783 1907 4807
rect 1945 4783 1975 4806
rect 1975 4783 1979 4806
rect 1801 4773 1835 4783
rect 1873 4773 1907 4783
rect 1945 4772 1979 4783
rect 1801 4714 1805 4734
rect 1805 4714 1835 4734
rect 1873 4714 1907 4734
rect 1945 4714 1975 4733
rect 1975 4714 1979 4733
rect 1801 4700 1835 4714
rect 1873 4700 1907 4714
rect 1945 4699 1979 4714
rect 1801 4645 1805 4661
rect 1805 4645 1835 4661
rect 1873 4645 1907 4661
rect 1945 4645 1975 4660
rect 1975 4645 1979 4660
rect 1801 4627 1835 4645
rect 1873 4627 1907 4645
rect 1945 4626 1979 4645
rect 1801 4576 1805 4588
rect 1805 4576 1835 4588
rect 1873 4576 1907 4588
rect 1945 4576 1975 4587
rect 1975 4576 1979 4587
rect 1801 4554 1835 4576
rect 1873 4554 1907 4576
rect 1945 4553 1979 4576
rect 1801 4507 1805 4515
rect 1805 4507 1835 4515
rect 1873 4507 1907 4515
rect 1945 4507 1975 4514
rect 1975 4507 1979 4514
rect 1801 4481 1835 4507
rect 1873 4481 1907 4507
rect 1945 4480 1979 4507
rect 1801 4438 1805 4442
rect 1805 4438 1835 4442
rect 1873 4438 1907 4442
rect 1945 4438 1975 4441
rect 1975 4438 1979 4441
rect 1801 4408 1835 4438
rect 1873 4408 1907 4438
rect 1945 4407 1979 4438
rect 1801 4335 1835 4369
rect 1873 4335 1907 4369
rect 1945 4334 1979 4368
rect 1801 4265 1835 4296
rect 1873 4265 1907 4296
rect 1945 4265 1979 4295
rect 1801 4262 1805 4265
rect 1805 4262 1835 4265
rect 1873 4262 1907 4265
rect 1945 4261 1975 4265
rect 1975 4261 1979 4265
rect 1801 4196 1835 4223
rect 1873 4196 1907 4223
rect 1945 4196 1979 4222
rect 1801 4189 1805 4196
rect 1805 4189 1835 4196
rect 1873 4189 1907 4196
rect 1945 4188 1975 4196
rect 1975 4188 1979 4196
rect 1801 4127 1835 4150
rect 1873 4127 1907 4150
rect 1945 4127 1979 4149
rect 1801 4116 1805 4127
rect 1805 4116 1835 4127
rect 1873 4116 1907 4127
rect 1945 4115 1975 4127
rect 1975 4115 1979 4127
rect 1801 4058 1835 4077
rect 1873 4058 1907 4077
rect 1945 4058 1979 4076
rect 1801 4043 1805 4058
rect 1805 4043 1835 4058
rect 1873 4043 1907 4058
rect 1945 4042 1975 4058
rect 1975 4042 1979 4058
rect 1801 3989 1835 4004
rect 1873 3989 1907 4004
rect 1945 3989 1979 4003
rect 1801 3970 1805 3989
rect 1805 3970 1835 3989
rect 1873 3970 1907 3989
rect 1945 3969 1975 3989
rect 1975 3969 1979 3989
rect 1801 3920 1835 3931
rect 1873 3920 1907 3931
rect 1945 3920 1979 3930
rect 1801 3897 1805 3920
rect 1805 3897 1835 3920
rect 1873 3897 1907 3920
rect 1945 3896 1975 3920
rect 1975 3896 1979 3920
rect 1801 3824 1805 3858
rect 1805 3824 1835 3858
rect 1873 3824 1907 3858
rect 1945 3823 1975 3857
rect 1975 3823 1979 3857
rect 1801 3751 1805 3785
rect 1805 3751 1835 3785
rect 1873 3751 1907 3785
rect 1945 3750 1975 3784
rect 1975 3750 1979 3784
rect 1801 3678 1805 3712
rect 1805 3678 1835 3712
rect 1873 3678 1907 3712
rect 1945 3677 1975 3711
rect 1975 3677 1979 3711
rect 1801 3605 1805 3639
rect 1805 3605 1835 3639
rect 1873 3605 1907 3639
rect 1945 3604 1975 3638
rect 1975 3604 1979 3638
rect 1801 3532 1805 3566
rect 1805 3532 1835 3566
rect 1873 3532 1907 3566
rect 1945 3531 1975 3565
rect 1975 3531 1979 3565
rect 1801 3459 1805 3493
rect 1805 3459 1835 3493
rect 1873 3459 1907 3493
rect 1945 3458 1975 3492
rect 1975 3458 1979 3492
rect 1801 3386 1805 3420
rect 1805 3386 1835 3420
rect 1873 3386 1907 3420
rect 1945 3385 1975 3419
rect 1975 3385 1979 3419
rect 1801 3313 1805 3347
rect 1805 3313 1835 3347
rect 1873 3313 1907 3347
rect 1945 3312 1975 3346
rect 1975 3312 1979 3346
rect 1801 3240 1805 3274
rect 1805 3240 1835 3274
rect 1873 3240 1907 3274
rect 1945 3239 1975 3273
rect 1975 3239 1979 3273
rect 1801 3167 1805 3201
rect 1805 3167 1835 3201
rect 1873 3167 1907 3201
rect 1945 3166 1975 3200
rect 1975 3166 1979 3200
rect 1801 3094 1805 3128
rect 1805 3094 1835 3128
rect 1873 3094 1907 3128
rect 1945 3093 1975 3127
rect 1975 3093 1979 3127
rect 1801 3021 1805 3055
rect 1805 3021 1835 3055
rect 1873 3021 1907 3055
rect 1945 3020 1975 3054
rect 1975 3020 1979 3054
rect 1801 2948 1805 2982
rect 1805 2948 1835 2982
rect 1873 2948 1907 2982
rect 1945 2947 1975 2981
rect 1975 2947 1979 2981
rect 1801 2875 1805 2909
rect 1805 2875 1835 2909
rect 1873 2875 1907 2909
rect 1945 2874 1975 2908
rect 1975 2874 1979 2908
rect 1801 2802 1805 2836
rect 1805 2802 1835 2836
rect 1873 2802 1907 2836
rect 1945 2801 1975 2835
rect 1975 2801 1979 2835
rect 1801 2729 1805 2763
rect 1805 2729 1835 2763
rect 1873 2729 1907 2763
rect 1945 2728 1975 2762
rect 1975 2728 1979 2762
rect 1801 2656 1805 2690
rect 1805 2656 1835 2690
rect 1873 2656 1907 2690
rect 1945 2655 1975 2689
rect 1975 2655 1979 2689
rect 1801 2583 1805 2617
rect 1805 2583 1835 2617
rect 1873 2583 1907 2617
rect 1945 2582 1975 2616
rect 1975 2582 1979 2616
rect 1801 2510 1805 2544
rect 1805 2510 1835 2544
rect 1873 2510 1907 2544
rect 1945 2509 1975 2543
rect 1975 2509 1979 2543
rect 1801 2437 1805 2471
rect 1805 2437 1835 2471
rect 1873 2437 1907 2471
rect 1945 2436 1975 2470
rect 1975 2436 1979 2470
rect 1801 2364 1805 2398
rect 1805 2364 1835 2398
rect 1873 2364 1907 2398
rect 1945 2363 1975 2397
rect 1975 2363 1979 2397
rect 1801 2291 1805 2325
rect 1805 2291 1835 2325
rect 1873 2291 1907 2325
rect 1945 2290 1975 2324
rect 1975 2290 1979 2324
rect 1801 2218 1805 2252
rect 1805 2218 1835 2252
rect 1873 2218 1907 2252
rect 2259 8458 2293 8461
rect 2332 8458 2366 8461
rect 2405 8458 2439 8461
rect 2478 8458 2512 8461
rect 2551 8458 2585 8461
rect 2624 8458 2658 8461
rect 2697 8458 2731 8461
rect 2770 8458 2804 8461
rect 2843 8458 2877 8461
rect 2916 8458 2950 8461
rect 2989 8458 3023 8461
rect 3062 8458 27216 8461
rect 2259 8427 2273 8458
rect 2273 8427 2293 8458
rect 2332 8427 2341 8458
rect 2341 8427 2366 8458
rect 2405 8427 2439 8458
rect 2478 8427 2512 8458
rect 2551 8427 2585 8458
rect 2624 8427 2658 8458
rect 2697 8427 2731 8458
rect 2770 8427 2804 8458
rect 2843 8427 2877 8458
rect 2916 8427 2950 8458
rect 2989 8427 3023 8458
rect 2187 5259 2191 8389
rect 2191 8317 2293 8389
rect 2332 8356 2341 8389
rect 2341 8356 2366 8389
rect 2405 8356 2439 8389
rect 2332 8355 2366 8356
rect 2405 8355 2409 8356
rect 2409 8355 2439 8356
rect 2478 8355 2512 8389
rect 2551 8355 2585 8389
rect 2624 8355 2658 8389
rect 2697 8355 2731 8389
rect 2770 8355 2804 8389
rect 2843 8355 2877 8389
rect 2916 8355 2950 8389
rect 2989 8355 3023 8389
rect 3062 8356 27195 8458
rect 27195 8356 27216 8458
rect 27254 8357 27288 8389
rect 3062 8355 27127 8356
rect 27127 8355 27216 8356
rect 27254 8355 27263 8357
rect 27263 8355 27288 8357
rect 2191 5331 2361 8317
rect 2361 5331 2365 8317
rect 2404 8288 2409 8317
rect 2409 8288 2438 8317
rect 2477 8288 2511 8317
rect 2550 8288 2584 8317
rect 2623 8288 2657 8317
rect 2696 8288 2730 8317
rect 2769 8288 2803 8317
rect 2842 8288 2876 8317
rect 2915 8288 2949 8317
rect 2988 8288 3022 8317
rect 3061 8288 3095 8317
rect 3134 8288 27127 8355
rect 27127 8288 27144 8355
rect 27182 8289 27216 8315
rect 27254 8289 27288 8315
rect 2404 8283 2438 8288
rect 2477 8283 2511 8288
rect 2550 8283 2584 8288
rect 2623 8283 2657 8288
rect 2696 8283 2730 8288
rect 2769 8283 2803 8288
rect 2842 8283 2876 8288
rect 2915 8283 2949 8288
rect 2988 8283 3022 8288
rect 3061 8283 3095 8288
rect 3134 8283 27144 8288
rect 27182 8281 27216 8289
rect 27254 8281 27263 8289
rect 27263 8281 27288 8289
rect 2191 5259 2293 5331
rect 2331 5258 2361 5292
rect 2361 5258 2365 5292
rect 2187 5186 2191 5220
rect 2191 5186 2221 5220
rect 2259 5186 2293 5220
rect 2331 5185 2361 5219
rect 2361 5185 2365 5219
rect 2187 5113 2191 5147
rect 2191 5113 2221 5147
rect 2259 5113 2293 5147
rect 2331 5112 2361 5146
rect 2361 5112 2365 5146
rect 2187 5040 2191 5074
rect 2191 5040 2221 5074
rect 2259 5040 2293 5074
rect 2331 5039 2361 5073
rect 2361 5039 2365 5073
rect 2187 4967 2191 5001
rect 2191 4967 2221 5001
rect 2259 4967 2293 5001
rect 2331 4966 2361 5000
rect 2361 4966 2365 5000
rect 2187 4894 2191 4928
rect 2191 4894 2221 4928
rect 2259 4894 2293 4928
rect 2331 4893 2361 4927
rect 2361 4893 2365 4927
rect 2187 4821 2191 4855
rect 2191 4821 2221 4855
rect 2259 4821 2293 4855
rect 2331 4820 2361 4854
rect 2361 4820 2365 4854
rect 2187 4748 2191 4782
rect 2191 4748 2221 4782
rect 2259 4748 2293 4782
rect 2331 4747 2361 4781
rect 2361 4747 2365 4781
rect 2187 4675 2191 4709
rect 2191 4675 2221 4709
rect 2259 4675 2293 4709
rect 2331 4674 2361 4708
rect 2361 4674 2365 4708
rect 2187 4602 2191 4636
rect 2191 4602 2221 4636
rect 2259 4602 2293 4636
rect 2331 4601 2361 4635
rect 2361 4601 2365 4635
rect 2187 4529 2191 4563
rect 2191 4529 2221 4563
rect 2259 4529 2293 4563
rect 2331 4528 2361 4562
rect 2361 4528 2365 4562
rect 2187 4456 2191 4490
rect 2191 4456 2221 4490
rect 2259 4456 2293 4490
rect 2331 4455 2361 4489
rect 2361 4455 2365 4489
rect 2187 4383 2191 4417
rect 2191 4383 2221 4417
rect 2259 4383 2293 4417
rect 2331 4382 2361 4416
rect 2361 4382 2365 4416
rect 2187 4310 2191 4344
rect 2191 4310 2221 4344
rect 2259 4310 2293 4344
rect 2331 4309 2361 4343
rect 2361 4309 2365 4343
rect 2187 4237 2191 4271
rect 2191 4237 2221 4271
rect 2259 4237 2293 4271
rect 2331 4236 2361 4270
rect 2361 4236 2365 4270
rect 2187 4164 2191 4198
rect 2191 4164 2221 4198
rect 2259 4164 2293 4198
rect 2331 4163 2361 4197
rect 2361 4163 2365 4197
rect 2187 4091 2191 4125
rect 2191 4091 2221 4125
rect 2259 4091 2293 4125
rect 2331 4090 2361 4124
rect 2361 4090 2365 4124
rect 2187 4018 2191 4052
rect 2191 4018 2221 4052
rect 2259 4018 2293 4052
rect 2331 4017 2361 4051
rect 2361 4017 2365 4051
rect 2187 3945 2191 3979
rect 2191 3945 2221 3979
rect 2259 3945 2293 3979
rect 2331 3944 2361 3978
rect 2361 3944 2365 3978
rect 2187 3872 2191 3906
rect 2191 3872 2221 3906
rect 2259 3872 2293 3906
rect 2331 3871 2361 3905
rect 2361 3871 2365 3905
rect 2187 3799 2191 3833
rect 2191 3799 2221 3833
rect 2259 3799 2293 3833
rect 2331 3798 2361 3832
rect 2361 3798 2365 3832
rect 2187 3726 2191 3760
rect 2191 3726 2221 3760
rect 2259 3726 2293 3760
rect 2331 3725 2361 3759
rect 2361 3725 2365 3759
rect 2187 3653 2191 3687
rect 2191 3653 2221 3687
rect 2259 3653 2293 3687
rect 2331 3652 2361 3686
rect 2361 3652 2365 3686
rect 2187 3580 2191 3614
rect 2191 3580 2221 3614
rect 2259 3580 2293 3614
rect 2331 3579 2361 3613
rect 2361 3579 2365 3613
rect 2187 3507 2191 3541
rect 2191 3507 2221 3541
rect 2259 3507 2293 3541
rect 2331 3506 2361 3540
rect 2361 3506 2365 3540
rect 2187 3434 2191 3468
rect 2191 3434 2221 3468
rect 2259 3434 2293 3468
rect 2331 3433 2361 3467
rect 2361 3433 2365 3467
rect 2187 3361 2191 3395
rect 2191 3361 2221 3395
rect 2259 3361 2293 3395
rect 2331 3360 2361 3394
rect 2361 3360 2365 3394
rect 2187 3288 2191 3322
rect 2191 3288 2221 3322
rect 2259 3288 2293 3322
rect 2331 3287 2361 3321
rect 2361 3287 2365 3321
rect 2187 3215 2191 3249
rect 2191 3215 2221 3249
rect 2259 3215 2293 3249
rect 2331 3214 2361 3248
rect 2361 3214 2365 3248
rect 2187 3142 2191 3176
rect 2191 3142 2221 3176
rect 2259 3142 2293 3176
rect 2331 3141 2361 3175
rect 2361 3141 2365 3175
rect 2187 3069 2191 3103
rect 2191 3069 2221 3103
rect 2259 3069 2293 3103
rect 2331 3068 2361 3102
rect 2361 3068 2365 3102
rect 2187 2996 2191 3030
rect 2191 2996 2221 3030
rect 2259 2996 2293 3030
rect 2331 2995 2361 3029
rect 2361 2995 2365 3029
rect 2187 2923 2191 2957
rect 2191 2923 2221 2957
rect 2259 2923 2293 2957
rect 2331 2922 2361 2956
rect 2361 2922 2365 2956
rect 2187 2850 2221 2884
rect 2259 2850 2293 2884
rect 2331 2849 2365 2883
rect 2187 2790 2221 2811
rect 2259 2790 2293 2811
rect 2331 2790 2365 2810
rect 2187 2777 2191 2790
rect 2191 2777 2221 2790
rect 2259 2777 2293 2790
rect 2331 2776 2361 2790
rect 2361 2776 2365 2790
rect 2187 2704 2191 2738
rect 2191 2704 2221 2738
rect 2259 2704 2293 2738
rect 2331 2703 2361 2737
rect 2361 2703 2365 2737
rect 2187 2631 2191 2665
rect 2191 2631 2221 2665
rect 2259 2631 2293 2665
rect 2331 2630 2361 2664
rect 2361 2630 2365 2664
rect 2187 2558 2191 2592
rect 2191 2558 2221 2592
rect 2259 2558 2293 2592
rect 2331 2557 2361 2591
rect 2361 2557 2365 2591
rect 2187 2485 2191 2519
rect 2191 2485 2221 2519
rect 2259 2485 2293 2519
rect 2331 2484 2361 2518
rect 2361 2484 2365 2518
rect 27110 8221 27144 8243
rect 27110 8209 27144 8221
rect 27182 8207 27216 8241
rect 27254 8207 27263 8241
rect 27263 8207 27288 8241
rect 27110 8135 27144 8169
rect 27182 8133 27216 8167
rect 27254 8133 27263 8167
rect 27263 8133 27288 8167
rect 27110 8061 27144 8095
rect 27182 8059 27216 8093
rect 27254 8059 27263 8093
rect 27263 8059 27288 8093
rect 27110 7987 27144 8021
rect 27182 7985 27216 8019
rect 27254 7985 27263 8019
rect 27263 7985 27288 8019
rect 27110 7913 27144 7947
rect 27182 7912 27216 7946
rect 27254 7912 27263 7946
rect 27263 7912 27288 7946
rect 27110 7839 27144 7873
rect 27182 7839 27216 7873
rect 27254 7839 27263 7873
rect 27263 7839 27288 7873
rect 27110 7729 27144 7763
rect 27182 7729 27216 7763
rect 27254 7729 27263 7763
rect 27263 7729 27288 7763
rect 27110 7656 27144 7690
rect 27182 7656 27216 7690
rect 27254 7656 27263 7690
rect 27263 7656 27288 7690
rect 27110 7583 27144 7617
rect 27182 7583 27216 7617
rect 27254 7583 27263 7617
rect 27263 7583 27288 7617
rect 27110 7510 27144 7544
rect 27182 7510 27216 7544
rect 27254 7510 27263 7544
rect 27263 7510 27288 7544
rect 27110 7437 27144 7471
rect 27182 7437 27216 7471
rect 27254 7437 27263 7471
rect 27263 7437 27288 7471
rect 27110 7364 27144 7398
rect 27182 7364 27216 7398
rect 27254 7364 27263 7398
rect 27263 7364 27288 7398
rect 27110 7291 27144 7325
rect 27182 7291 27216 7325
rect 27254 7291 27263 7325
rect 27263 7291 27288 7325
rect 27110 7218 27144 7252
rect 27182 7218 27216 7252
rect 27254 7218 27263 7252
rect 27263 7218 27288 7252
rect 27110 7145 27144 7179
rect 27182 7145 27216 7179
rect 27254 7145 27263 7179
rect 27263 7145 27288 7179
rect 27110 7072 27144 7106
rect 27182 7072 27216 7106
rect 27254 7072 27263 7106
rect 27263 7072 27288 7106
rect 27110 6999 27144 7033
rect 27182 6999 27216 7033
rect 27254 6999 27263 7033
rect 27263 6999 27288 7033
rect 27110 6926 27144 6960
rect 27182 6926 27216 6960
rect 27254 6926 27263 6960
rect 27263 6926 27288 6960
rect 27110 6853 27144 6887
rect 27182 6853 27216 6887
rect 27254 6853 27263 6887
rect 27263 6853 27288 6887
rect 27110 6780 27144 6814
rect 27182 6780 27216 6814
rect 27254 6780 27263 6814
rect 27263 6780 27288 6814
rect 27110 6707 27144 6741
rect 27182 6707 27216 6741
rect 27254 6707 27263 6741
rect 27263 6707 27288 6741
rect 27110 6634 27144 6668
rect 27182 6634 27216 6668
rect 27254 6634 27263 6668
rect 27263 6634 27288 6668
rect 27110 6561 27144 6595
rect 27182 6561 27216 6595
rect 27254 6561 27263 6595
rect 27263 6561 27288 6595
rect 27110 6488 27144 6522
rect 27182 6488 27216 6522
rect 27254 6488 27263 6522
rect 27263 6488 27288 6522
rect 27110 6415 27144 6449
rect 27182 6415 27216 6449
rect 27254 6415 27263 6449
rect 27263 6415 27288 6449
rect 27110 6342 27144 6376
rect 27182 6342 27216 6376
rect 27254 6342 27263 6376
rect 27263 6342 27288 6376
rect 27110 6269 27144 6303
rect 27182 6269 27216 6303
rect 27254 6269 27263 6303
rect 27263 6269 27288 6303
rect 27110 6196 27144 6230
rect 27182 6196 27216 6230
rect 27254 6196 27263 6230
rect 27263 6196 27288 6230
rect 27110 6123 27144 6157
rect 27182 6123 27216 6157
rect 27254 6123 27263 6157
rect 27263 6123 27288 6157
rect 27110 6050 27144 6084
rect 27182 6050 27216 6084
rect 27254 6050 27263 6084
rect 27263 6050 27288 6084
rect 27110 5977 27144 6011
rect 27182 5977 27216 6011
rect 27254 5977 27263 6011
rect 27263 5977 27288 6011
rect 27110 5904 27144 5938
rect 27182 5904 27216 5938
rect 27254 5904 27263 5938
rect 27263 5904 27288 5938
rect 27110 5831 27144 5865
rect 27182 5831 27216 5865
rect 27254 5831 27263 5865
rect 27263 5831 27288 5865
rect 27110 5758 27144 5792
rect 27182 5758 27216 5792
rect 27254 5758 27263 5792
rect 27263 5758 27288 5792
rect 27110 5685 27144 5719
rect 27182 5685 27216 5719
rect 27254 5685 27263 5719
rect 27263 5685 27288 5719
rect 27110 5612 27144 5646
rect 27182 5612 27216 5646
rect 27254 5612 27263 5646
rect 27263 5612 27288 5646
rect 27110 5539 27144 5573
rect 27182 5539 27216 5573
rect 27254 5539 27263 5573
rect 27263 5539 27288 5573
rect 27110 5466 27144 5500
rect 27182 5466 27216 5500
rect 27254 5466 27263 5500
rect 27263 5466 27288 5500
rect 27110 5393 27144 5427
rect 27182 5393 27216 5427
rect 27254 5393 27263 5427
rect 27263 5393 27288 5427
rect 27110 5320 27144 5354
rect 27182 5320 27216 5354
rect 27254 5320 27263 5354
rect 27263 5320 27288 5354
rect 27110 5247 27144 5281
rect 27182 5247 27216 5281
rect 27254 5247 27263 5281
rect 27263 5247 27288 5281
rect 27110 5174 27144 5208
rect 27182 5174 27216 5208
rect 27254 5174 27263 5208
rect 27263 5174 27288 5208
rect 27110 5101 27144 5135
rect 27182 5101 27216 5135
rect 27254 5101 27263 5135
rect 27263 5101 27288 5135
rect 27110 5028 27144 5062
rect 27182 5028 27216 5062
rect 27254 5028 27263 5062
rect 27263 5028 27288 5062
rect 27110 4955 27144 4989
rect 27182 4955 27216 4989
rect 27254 4955 27263 4989
rect 27263 4955 27288 4989
rect 27110 4882 27144 4916
rect 27182 4882 27216 4916
rect 27254 4882 27263 4916
rect 27263 4882 27288 4916
rect 27110 4809 27144 4843
rect 27182 4809 27216 4843
rect 27254 4809 27263 4843
rect 27263 4809 27288 4843
rect 27110 4736 27144 4770
rect 27182 4736 27216 4770
rect 27254 4736 27263 4770
rect 27263 4736 27288 4770
rect 27110 4663 27144 4697
rect 27182 4663 27216 4697
rect 27254 4663 27263 4697
rect 27263 4663 27288 4697
rect 27110 4590 27144 4624
rect 27182 4590 27216 4624
rect 27254 4590 27263 4624
rect 27263 4590 27288 4624
rect 27110 4517 27144 4551
rect 27182 4517 27216 4551
rect 27254 4517 27263 4551
rect 27263 4517 27288 4551
rect 27110 4444 27144 4478
rect 27182 4444 27216 4478
rect 27254 4444 27263 4478
rect 27263 4444 27288 4478
rect 27110 4371 27144 4405
rect 27182 4371 27216 4405
rect 27254 4371 27263 4405
rect 27263 4371 27288 4405
rect 27110 4298 27144 4332
rect 27182 4298 27216 4332
rect 27254 4298 27263 4332
rect 27263 4298 27288 4332
rect 27110 4225 27144 4259
rect 27182 4225 27216 4259
rect 27254 4225 27263 4259
rect 27263 4225 27288 4259
rect 27110 4152 27144 4186
rect 27182 4152 27216 4186
rect 27254 4152 27263 4186
rect 27263 4152 27288 4186
rect 27110 4079 27144 4113
rect 27182 4079 27216 4113
rect 27254 4079 27263 4113
rect 27263 4079 27288 4113
rect 27110 4006 27144 4040
rect 27182 4006 27216 4040
rect 27254 4006 27263 4040
rect 27263 4006 27288 4040
rect 27110 3933 27144 3967
rect 27182 3933 27216 3967
rect 27254 3933 27263 3967
rect 27263 3933 27288 3967
rect 27110 3860 27144 3894
rect 27182 3860 27216 3894
rect 27254 3860 27263 3894
rect 27263 3860 27288 3894
rect 27110 3787 27144 3821
rect 27182 3787 27216 3821
rect 27254 3787 27263 3821
rect 27263 3787 27288 3821
rect 27110 3714 27144 3748
rect 27182 3714 27216 3748
rect 27254 3714 27263 3748
rect 27263 3714 27288 3748
rect 27110 3641 27144 3675
rect 27182 3641 27216 3675
rect 27254 3641 27263 3675
rect 27263 3641 27288 3675
rect 27110 3568 27144 3602
rect 27182 3568 27216 3602
rect 27254 3568 27263 3602
rect 27263 3568 27288 3602
rect 27110 3495 27144 3529
rect 27182 3495 27216 3529
rect 27254 3495 27263 3529
rect 27263 3495 27288 3529
rect 27110 3422 27144 3456
rect 27182 3422 27216 3456
rect 27254 3422 27263 3456
rect 27263 3422 27288 3456
rect 27110 3349 27144 3383
rect 27182 3349 27216 3383
rect 27254 3349 27263 3383
rect 27263 3349 27288 3383
rect 27110 3276 27144 3310
rect 27182 3276 27216 3310
rect 27254 3276 27263 3310
rect 27263 3276 27288 3310
rect 2187 2416 2191 2446
rect 2191 2416 2221 2446
rect 2259 2416 2293 2446
rect 2331 2441 26341 2445
rect 26380 2441 26414 2445
rect 26453 2441 26487 2445
rect 26526 2441 26560 2445
rect 26599 2441 26633 2445
rect 26672 2441 26706 2445
rect 26745 2441 26779 2445
rect 26818 2441 26852 2445
rect 26891 2441 26925 2445
rect 26964 2441 26998 2445
rect 27037 2441 27071 2445
rect 2187 2412 2221 2416
rect 2259 2412 2293 2416
rect 2331 2373 26341 2441
rect 26380 2411 26414 2441
rect 26453 2411 26487 2441
rect 26526 2411 26560 2441
rect 26599 2411 26633 2441
rect 26672 2411 26706 2441
rect 26745 2411 26779 2441
rect 26818 2411 26852 2441
rect 26891 2411 26925 2441
rect 26964 2411 26998 2441
rect 27037 2411 27045 2441
rect 27045 2411 27071 2441
rect 27110 2411 27263 3237
rect 2187 2348 2191 2373
rect 2191 2348 2221 2373
rect 2187 2339 2221 2348
rect 2259 2271 26413 2373
rect 26452 2339 26486 2373
rect 26525 2339 26559 2373
rect 26598 2339 26632 2373
rect 26671 2339 26705 2373
rect 26744 2339 26778 2373
rect 26817 2339 26851 2373
rect 26890 2339 26924 2373
rect 26963 2339 26997 2373
rect 27036 2339 27070 2373
rect 27109 2339 27113 2373
rect 27113 2339 27143 2373
rect 27182 2339 27263 2411
rect 27263 2339 27288 3237
rect 26452 2271 26486 2301
rect 26525 2271 26559 2301
rect 26598 2271 26632 2301
rect 26671 2271 26705 2301
rect 26744 2271 26778 2301
rect 26817 2271 26851 2301
rect 26890 2271 26924 2301
rect 26963 2271 26997 2301
rect 27036 2271 27070 2301
rect 27109 2271 27113 2301
rect 27113 2271 27143 2301
rect 2259 2267 26413 2271
rect 26452 2267 26486 2271
rect 26525 2267 26559 2271
rect 26598 2267 26632 2271
rect 26671 2267 26705 2271
rect 26744 2267 26778 2271
rect 26817 2267 26851 2271
rect 26890 2267 26924 2271
rect 26963 2267 26997 2271
rect 27036 2267 27070 2271
rect 27109 2267 27143 2271
rect 27182 2267 27216 2301
rect 27508 8447 27512 8481
rect 27512 8447 27542 8481
rect 27580 8445 27614 8479
rect 27652 8445 27682 8479
rect 27682 8445 27686 8479
rect 27508 8373 27512 8407
rect 27512 8373 27542 8407
rect 27580 8371 27614 8405
rect 27652 8371 27682 8405
rect 27682 8371 27686 8405
rect 27508 8299 27512 8333
rect 27512 8299 27542 8333
rect 27580 8298 27614 8332
rect 27652 8298 27682 8332
rect 27682 8298 27686 8332
rect 27508 8225 27512 8259
rect 27512 8225 27542 8259
rect 27580 8225 27614 8259
rect 27652 8225 27682 8259
rect 27682 8225 27686 8259
rect 27508 8115 27512 8149
rect 27512 8115 27542 8149
rect 27580 8115 27614 8149
rect 27652 8115 27682 8149
rect 27682 8115 27686 8149
rect 27508 8042 27512 8076
rect 27512 8042 27542 8076
rect 27580 8042 27614 8076
rect 27652 8042 27682 8076
rect 27682 8042 27686 8076
rect 27508 7969 27512 8003
rect 27512 7969 27542 8003
rect 27580 7969 27614 8003
rect 27652 7969 27682 8003
rect 27682 7969 27686 8003
rect 27508 7896 27512 7930
rect 27512 7896 27542 7930
rect 27580 7896 27614 7930
rect 27652 7896 27682 7930
rect 27682 7896 27686 7930
rect 27508 7823 27512 7857
rect 27512 7823 27542 7857
rect 27580 7823 27614 7857
rect 27652 7823 27682 7857
rect 27682 7823 27686 7857
rect 1945 2217 1975 2251
rect 1975 2217 1979 2251
rect 1801 2145 1805 2179
rect 1805 2145 1835 2179
rect 1873 2145 1907 2179
rect 1945 2144 1975 2178
rect 1975 2144 1979 2178
rect 1801 2072 1805 2106
rect 1805 2072 1835 2106
rect 1873 2072 1907 2106
rect 1945 2071 1975 2105
rect 1975 2071 1979 2105
rect 1801 1999 1805 2033
rect 1805 1999 1835 2033
rect 1873 1999 1907 2033
rect 1945 1998 1975 2032
rect 1975 1998 1979 2032
rect 27508 3301 27512 7784
rect 27512 3301 27682 7784
rect 27508 3266 27580 3301
rect 27508 3232 27512 3266
rect 27512 3232 27546 3266
rect 27546 3233 27580 3266
rect 27580 3233 27682 3301
rect 27682 3233 27686 7784
rect 27546 3232 27686 3233
rect 27508 3198 27686 3232
rect 27508 3197 27580 3198
rect 27508 3163 27512 3197
rect 27512 3163 27546 3197
rect 27546 3164 27580 3197
rect 27580 3164 27614 3198
rect 27614 3164 27648 3198
rect 27648 3164 27682 3198
rect 27682 3164 27686 3198
rect 27546 3163 27686 3164
rect 27508 3129 27686 3163
rect 27508 3128 27580 3129
rect 27508 3094 27512 3128
rect 27512 3094 27546 3128
rect 27546 3095 27580 3128
rect 27580 3095 27614 3129
rect 27614 3095 27648 3129
rect 27648 3095 27682 3129
rect 27682 3095 27686 3129
rect 27546 3094 27686 3095
rect 27508 3060 27686 3094
rect 27508 3059 27580 3060
rect 27508 3025 27512 3059
rect 27512 3025 27546 3059
rect 27546 3026 27580 3059
rect 27580 3026 27614 3060
rect 27614 3026 27648 3060
rect 27648 3026 27682 3060
rect 27682 3026 27686 3060
rect 27546 3025 27686 3026
rect 27508 2991 27686 3025
rect 27508 2990 27580 2991
rect 27508 2956 27512 2990
rect 27512 2956 27546 2990
rect 27546 2957 27580 2990
rect 27580 2957 27614 2991
rect 27614 2957 27648 2991
rect 27648 2957 27682 2991
rect 27682 2957 27686 2991
rect 27546 2956 27686 2957
rect 27508 2922 27686 2956
rect 27508 2921 27580 2922
rect 27508 2887 27512 2921
rect 27512 2887 27546 2921
rect 27546 2888 27580 2921
rect 27580 2888 27614 2922
rect 27614 2888 27648 2922
rect 27648 2888 27682 2922
rect 27682 2888 27686 2922
rect 27546 2887 27686 2888
rect 27508 2853 27686 2887
rect 27508 2852 27580 2853
rect 27508 2818 27512 2852
rect 27512 2818 27546 2852
rect 27546 2819 27580 2852
rect 27580 2819 27614 2853
rect 27614 2819 27648 2853
rect 27648 2819 27682 2853
rect 27682 2819 27686 2853
rect 27546 2818 27686 2819
rect 27508 2784 27686 2818
rect 27508 2783 27580 2784
rect 27508 2749 27512 2783
rect 27512 2749 27546 2783
rect 27546 2750 27580 2783
rect 27580 2750 27614 2784
rect 27614 2750 27648 2784
rect 27648 2750 27682 2784
rect 27682 2750 27686 2784
rect 27546 2749 27686 2750
rect 27508 2715 27686 2749
rect 27508 2714 27580 2715
rect 27508 2680 27512 2714
rect 27512 2680 27546 2714
rect 27546 2681 27580 2714
rect 27580 2681 27614 2715
rect 27614 2681 27648 2715
rect 27648 2681 27682 2715
rect 27682 2681 27686 2715
rect 27546 2680 27686 2681
rect 27508 2646 27686 2680
rect 27508 2645 27580 2646
rect 27508 2611 27512 2645
rect 27512 2611 27546 2645
rect 27546 2612 27580 2645
rect 27580 2612 27614 2646
rect 27614 2612 27648 2646
rect 27648 2612 27682 2646
rect 27682 2612 27686 2646
rect 27546 2611 27686 2612
rect 27508 2577 27686 2611
rect 27508 2576 27580 2577
rect 27508 2542 27512 2576
rect 27512 2542 27546 2576
rect 27546 2543 27580 2576
rect 27580 2543 27614 2577
rect 27614 2543 27648 2577
rect 27648 2543 27682 2577
rect 27682 2543 27686 2577
rect 27546 2542 27686 2543
rect 27508 2508 27686 2542
rect 27508 2507 27580 2508
rect 27508 2473 27512 2507
rect 27512 2473 27546 2507
rect 27546 2474 27580 2507
rect 27580 2474 27614 2508
rect 27614 2474 27648 2508
rect 27648 2474 27682 2508
rect 27682 2474 27686 2508
rect 27546 2473 27686 2474
rect 27508 2439 27686 2473
rect 27508 2438 27580 2439
rect 27508 2404 27512 2438
rect 27512 2404 27546 2438
rect 27546 2405 27580 2438
rect 27580 2405 27614 2439
rect 27614 2405 27648 2439
rect 27648 2405 27682 2439
rect 27682 2405 27686 2439
rect 27546 2404 27686 2405
rect 27508 2370 27686 2404
rect 27508 2369 27580 2370
rect 27508 2335 27512 2369
rect 27512 2335 27546 2369
rect 27546 2336 27580 2369
rect 27580 2336 27614 2370
rect 27614 2336 27648 2370
rect 27648 2336 27682 2370
rect 27682 2336 27686 2370
rect 27546 2335 27686 2336
rect 27508 2301 27686 2335
rect 27508 2300 27580 2301
rect 27508 2266 27512 2300
rect 27512 2266 27546 2300
rect 27546 2267 27580 2300
rect 27580 2267 27614 2301
rect 27614 2267 27648 2301
rect 27648 2267 27682 2301
rect 27682 2267 27686 2301
rect 27546 2266 27686 2267
rect 27508 2232 27686 2266
rect 27508 2231 27580 2232
rect 27508 2197 27512 2231
rect 27512 2197 27546 2231
rect 27546 2198 27580 2231
rect 27580 2198 27614 2232
rect 27614 2198 27648 2232
rect 27648 2198 27682 2232
rect 27682 2198 27686 2232
rect 27546 2197 27686 2198
rect 27508 2163 27686 2197
rect 27508 2162 27580 2163
rect 27508 2128 27512 2162
rect 27512 2128 27546 2162
rect 27546 2129 27580 2162
rect 27580 2129 27614 2163
rect 27614 2129 27648 2163
rect 27648 2129 27682 2163
rect 27682 2129 27686 2163
rect 27546 2128 27686 2129
rect 27508 2094 27686 2128
rect 27508 2093 27580 2094
rect 27508 2059 27512 2093
rect 27512 2059 27546 2093
rect 27546 2060 27580 2093
rect 27580 2060 27614 2094
rect 27614 2060 27648 2094
rect 27648 2060 27682 2094
rect 27682 2060 27686 2094
rect 27546 2059 27686 2060
rect 27508 2025 27686 2059
rect 27508 2024 27580 2025
rect 27508 1990 27512 2024
rect 27512 1990 27546 2024
rect 27546 1991 27580 2024
rect 27580 1991 27614 2025
rect 27614 1991 27648 2025
rect 27648 1991 27682 2025
rect 27682 1991 27686 2025
rect 27546 1990 27686 1991
rect 1801 1926 1805 1960
rect 1805 1926 1835 1960
rect 1873 1926 1907 1960
rect 1945 1925 1975 1959
rect 1975 1925 1979 1959
rect 27508 1956 27686 1990
rect 27508 1955 27580 1956
rect 27508 1921 27512 1955
rect 27512 1921 27546 1955
rect 27546 1922 27580 1955
rect 27580 1922 27614 1956
rect 27614 1922 27648 1956
rect 27648 1922 27682 1956
rect 27682 1922 27686 1956
rect 27546 1921 27686 1922
rect 27508 1887 27686 1921
rect 1801 1853 1805 1887
rect 1805 1853 1835 1887
rect 1873 1853 1907 1887
rect 27508 1886 27580 1887
rect 1945 1852 1975 1886
rect 1975 1852 1979 1886
rect 27508 1852 27512 1886
rect 27512 1852 27546 1886
rect 27546 1853 27580 1886
rect 27580 1853 27614 1887
rect 27614 1853 27648 1887
rect 27648 1853 27682 1887
rect 27682 1853 27686 1887
rect 27546 1852 27686 1853
rect 1801 1780 1805 1814
rect 1805 1780 1835 1814
rect 1873 1780 1907 1814
rect 27508 1818 27686 1852
rect 27508 1817 27580 1818
rect 1945 1779 1975 1813
rect 1975 1779 1979 1813
rect 27508 1783 27512 1817
rect 27512 1783 27546 1817
rect 27546 1784 27580 1817
rect 27580 1784 27614 1818
rect 27614 1784 27648 1818
rect 27648 1784 27682 1818
rect 27682 1784 27686 1818
rect 27546 1783 27686 1784
rect 1801 1707 1805 1741
rect 1805 1707 1835 1741
rect 1873 1707 1907 1741
rect 1945 1706 1975 1740
rect 1975 1706 1979 1740
rect 27508 1749 27686 1783
rect 27508 1748 27580 1749
rect 27508 1714 27512 1748
rect 27512 1714 27546 1748
rect 27546 1715 27580 1748
rect 27580 1715 27614 1749
rect 27614 1715 27648 1749
rect 27648 1715 27682 1749
rect 27682 1715 27686 1749
rect 27546 1714 27686 1715
rect 1801 1634 1805 1668
rect 1805 1634 1835 1668
rect 1873 1634 1907 1668
rect 1945 1633 1975 1667
rect 1975 1633 1979 1667
rect 27508 1680 27686 1714
rect 27508 1679 27580 1680
rect 27508 1645 27512 1679
rect 27512 1645 27546 1679
rect 27546 1646 27580 1679
rect 27580 1646 27614 1680
rect 27614 1646 27648 1680
rect 27648 1646 27682 1680
rect 27682 1646 27686 1680
rect 27546 1645 27686 1646
rect 1801 1561 1805 1595
rect 1805 1561 1835 1595
rect 1873 1561 1907 1595
rect 1945 1560 1975 1594
rect 1975 1560 1979 1594
rect 27508 1611 27686 1645
rect 27508 1610 27580 1611
rect 27508 1576 27512 1610
rect 27512 1576 27546 1610
rect 27546 1577 27580 1610
rect 27580 1577 27614 1611
rect 27614 1577 27648 1611
rect 27648 1577 27682 1611
rect 27682 1577 27686 1611
rect 27546 1576 27686 1577
rect 1801 1488 1805 1522
rect 1805 1488 1835 1522
rect 1873 1488 1907 1522
rect 1945 1487 1975 1521
rect 1975 1487 1979 1521
rect 27508 1542 27686 1576
rect 27508 1541 27580 1542
rect 27508 1507 27512 1541
rect 27512 1507 27546 1541
rect 27546 1508 27580 1541
rect 27580 1508 27614 1542
rect 27614 1508 27648 1542
rect 27648 1508 27682 1542
rect 27682 1508 27686 1542
rect 27546 1507 27686 1508
rect 27508 1473 27686 1507
rect 27508 1472 27580 1473
rect 1801 1415 1805 1449
rect 1805 1415 1835 1449
rect 1873 1415 1907 1449
rect 1945 1438 1975 1448
rect 1975 1438 2010 1448
rect 2010 1438 2044 1448
rect 2044 1438 2079 1448
rect 2079 1438 2113 1448
rect 2113 1438 2148 1448
rect 1945 1404 2148 1438
rect 2148 1404 27323 1448
rect 27362 1414 27396 1448
rect 27435 1414 27469 1448
rect 27508 1414 27546 1472
rect 27546 1439 27580 1472
rect 27580 1439 27614 1473
rect 27614 1439 27648 1473
rect 27648 1439 27682 1473
rect 27682 1439 27686 1473
rect 27546 1414 27686 1439
rect 27580 1404 27686 1414
rect 1945 1376 1976 1404
rect 1801 1370 1805 1376
rect 1805 1370 1835 1376
rect 1873 1370 1907 1376
rect 1907 1370 1942 1376
rect 1942 1370 1976 1376
rect 1976 1370 2011 1404
rect 2011 1370 2045 1404
rect 2045 1370 2080 1404
rect 2080 1376 27323 1404
rect 1801 1342 1835 1370
rect 1873 1336 2080 1370
rect 1873 1302 1907 1336
rect 1907 1302 1942 1336
rect 1942 1302 1976 1336
rect 1976 1302 2011 1336
rect 2011 1302 2045 1336
rect 2045 1302 2080 1336
rect 2080 1302 27395 1376
rect 27434 1342 27468 1376
rect 27507 1342 27541 1376
rect 27580 1342 27614 1404
rect 27614 1370 27648 1404
rect 27648 1370 27682 1404
rect 27682 1370 27686 1404
rect 27614 1342 27686 1370
rect 27434 1302 27468 1304
rect 27507 1302 27541 1304
rect 27580 1302 27614 1304
rect 1873 1270 27395 1302
rect 27434 1270 27468 1302
rect 27507 1270 27541 1302
rect 27580 1270 27614 1302
rect 27911 8841 27915 8875
rect 27915 8841 27945 8875
rect 27983 8841 28017 8875
rect 28055 8841 28085 8875
rect 28085 8841 28089 8875
rect 27911 8762 27915 8796
rect 27915 8762 27945 8796
rect 27983 8762 28017 8796
rect 28055 8762 28085 8796
rect 28085 8762 28089 8796
rect 27911 8683 27915 8717
rect 27915 8683 27945 8717
rect 27983 8683 28017 8717
rect 28055 8683 28085 8717
rect 28085 8683 28089 8717
rect 27911 8604 27915 8638
rect 27915 8604 27945 8638
rect 27983 8604 28017 8638
rect 28055 8604 28085 8638
rect 28085 8604 28089 8638
rect 27911 8494 27915 8528
rect 27915 8494 27945 8528
rect 27983 8494 28017 8528
rect 28055 8494 28085 8528
rect 28085 8494 28089 8528
rect 27911 8421 27915 8455
rect 27915 8421 27945 8455
rect 27983 8421 28017 8455
rect 28055 8421 28085 8455
rect 28085 8421 28089 8455
rect 27911 8348 27915 8382
rect 27915 8348 27945 8382
rect 27983 8348 28017 8382
rect 28055 8348 28085 8382
rect 28085 8348 28089 8382
rect 27911 8275 27915 8309
rect 27915 8275 27945 8309
rect 27983 8275 28017 8309
rect 28055 8275 28085 8309
rect 28085 8275 28089 8309
rect 1353 1189 1357 1223
rect 1357 1189 1387 1223
rect 1425 1189 1459 1223
rect 1497 1188 1527 1222
rect 1527 1188 1531 1222
rect 1353 1116 1357 1150
rect 1357 1116 1387 1150
rect 1425 1116 1459 1150
rect 1497 1115 1527 1149
rect 1527 1115 1531 1149
rect 1353 1043 1357 1077
rect 1357 1043 1387 1077
rect 1425 1043 1459 1077
rect 1497 1004 1527 1076
rect 1353 970 1357 1004
rect 1357 970 1387 1004
rect 1425 978 1527 1004
rect 1527 978 23779 1076
rect 23818 1042 23852 1076
rect 23891 1042 23925 1076
rect 23964 1042 23998 1076
rect 24037 1042 24071 1076
rect 24110 1042 24144 1076
rect 24183 1042 24217 1076
rect 24256 1042 24290 1076
rect 24329 1042 24363 1076
rect 24402 1042 24436 1076
rect 24475 1042 24509 1076
rect 24548 1042 24582 1076
rect 24621 1042 24655 1076
rect 24694 1042 24728 1076
rect 24767 1042 24801 1076
rect 24840 1042 24874 1076
rect 24913 1042 24947 1076
rect 24986 1042 25020 1076
rect 25059 1042 25093 1076
rect 25132 1042 25166 1076
rect 25205 1042 25239 1076
rect 25278 1042 25312 1076
rect 25351 1042 25385 1076
rect 25424 1042 25458 1076
rect 25497 1042 25531 1076
rect 25570 1042 25604 1076
rect 25643 1042 25677 1076
rect 25716 1042 25750 1076
rect 25789 1042 25823 1076
rect 25862 1042 25896 1076
rect 25935 1042 25969 1076
rect 26008 1042 26042 1076
rect 26081 1042 26115 1076
rect 26154 1042 26188 1076
rect 26227 1042 26261 1076
rect 26300 1042 26334 1076
rect 26373 1042 26407 1076
rect 26446 1042 26480 1076
rect 26519 1042 26553 1076
rect 26592 1042 26626 1076
rect 26665 1042 26699 1076
rect 26738 1042 26772 1076
rect 26811 1042 26845 1076
rect 26884 1042 26918 1076
rect 26957 1042 26991 1076
rect 27030 1042 27064 1076
rect 27103 1042 27137 1076
rect 27176 1042 27210 1076
rect 27249 1042 27283 1076
rect 27322 1042 27356 1076
rect 27395 1042 27429 1076
rect 27468 1042 27502 1076
rect 27541 1042 27575 1076
rect 27614 1042 27648 1076
rect 27687 1042 27721 1076
rect 27760 1042 27794 1076
rect 27833 1042 27867 1076
rect 23818 978 23852 1004
rect 23891 978 23925 1004
rect 23964 978 23998 1004
rect 24037 978 24071 1004
rect 24110 978 24144 1004
rect 24183 978 24217 1004
rect 24256 978 24290 1004
rect 24329 978 24363 1004
rect 24402 978 24436 1004
rect 24475 978 24509 1004
rect 24548 978 24582 1004
rect 24621 978 24655 1004
rect 24694 978 24728 1004
rect 24767 978 24801 1004
rect 24840 978 24874 1004
rect 24913 978 24947 1004
rect 24986 978 25020 1004
rect 25059 978 25093 1004
rect 25132 978 25166 1004
rect 25205 978 25239 1004
rect 25278 978 25312 1004
rect 25351 978 25385 1004
rect 25424 978 25458 1004
rect 25497 978 25531 1004
rect 25570 978 25604 1004
rect 25643 978 25677 1004
rect 25716 978 25750 1004
rect 25789 978 25823 1004
rect 25862 978 25896 1004
rect 25935 978 25969 1004
rect 26008 978 26042 1004
rect 26081 978 26115 1004
rect 26154 978 26188 1004
rect 26227 978 26261 1004
rect 26300 978 26334 1004
rect 26373 978 26407 1004
rect 26446 978 26480 1004
rect 26519 978 26553 1004
rect 26592 978 26626 1004
rect 26665 978 26699 1004
rect 26738 978 26772 1004
rect 26811 978 26845 1004
rect 26884 978 26918 1004
rect 26957 978 26991 1004
rect 27030 978 27064 1004
rect 27103 978 27137 1004
rect 27176 978 27210 1004
rect 27249 978 27283 1004
rect 27322 978 27356 1004
rect 27395 978 27429 1004
rect 27468 978 27502 1004
rect 27541 978 27575 1004
rect 27614 978 27648 1004
rect 27687 978 27721 1004
rect 27760 978 27794 1004
rect 27833 978 27867 1004
rect 27911 978 27915 8236
rect 27915 978 28085 8236
rect 1425 898 1595 978
rect 1595 944 1630 978
rect 1630 944 1664 978
rect 1664 944 1699 978
rect 1699 944 1733 978
rect 1733 944 1768 978
rect 1768 944 1802 978
rect 1802 944 1837 978
rect 1837 944 1871 978
rect 1871 944 1906 978
rect 1906 944 1940 978
rect 1940 944 1975 978
rect 1975 944 2009 978
rect 2009 944 2044 978
rect 2044 944 2078 978
rect 2078 944 2113 978
rect 2113 944 2147 978
rect 2147 944 2182 978
rect 2182 944 2216 978
rect 2216 944 2251 978
rect 2251 944 2285 978
rect 2285 944 2320 978
rect 2320 944 2354 978
rect 2354 944 2389 978
rect 2389 944 2423 978
rect 2423 944 2458 978
rect 2458 944 2492 978
rect 2492 944 2527 978
rect 2527 944 2561 978
rect 2561 944 2596 978
rect 2596 944 2630 978
rect 2630 944 2665 978
rect 2665 944 2699 978
rect 2699 944 2734 978
rect 2734 944 2768 978
rect 2768 944 2803 978
rect 2803 944 2837 978
rect 2837 944 2872 978
rect 2872 944 2906 978
rect 2906 944 2941 978
rect 2941 944 2975 978
rect 2975 944 3010 978
rect 3010 944 3044 978
rect 3044 944 3079 978
rect 3079 944 3113 978
rect 3113 944 3148 978
rect 3148 944 3182 978
rect 3182 944 3217 978
rect 3217 944 3251 978
rect 3251 944 3286 978
rect 3286 944 3320 978
rect 3320 944 3355 978
rect 3355 944 3389 978
rect 3389 944 3424 978
rect 3424 944 3458 978
rect 3458 944 3493 978
rect 3493 944 3527 978
rect 3527 944 3562 978
rect 3562 944 3596 978
rect 3596 944 3631 978
rect 3631 944 3665 978
rect 3665 944 3700 978
rect 3700 944 3734 978
rect 3734 944 3769 978
rect 3769 944 3803 978
rect 3803 944 3838 978
rect 3838 944 3872 978
rect 3872 944 3907 978
rect 3907 944 3941 978
rect 3941 944 3976 978
rect 3976 944 4010 978
rect 4010 944 4045 978
rect 4045 944 4079 978
rect 4079 944 4114 978
rect 4114 944 4148 978
rect 4148 944 4183 978
rect 1595 910 4183 944
rect 1595 898 1630 910
rect 1630 898 1664 910
rect 1664 898 1699 910
rect 1699 898 1733 910
rect 1733 898 1768 910
rect 1768 898 1802 910
rect 1802 898 1837 910
rect 1837 898 1871 910
rect 1871 898 1906 910
rect 1906 898 1940 910
rect 1940 898 1975 910
rect 1975 898 2009 910
rect 2009 898 2044 910
rect 2044 898 2078 910
rect 2078 898 2113 910
rect 2113 898 2147 910
rect 2147 898 2182 910
rect 2182 898 2216 910
rect 2216 898 2251 910
rect 2251 898 2285 910
rect 2285 898 2320 910
rect 2320 898 2354 910
rect 2354 898 2389 910
rect 2389 898 2423 910
rect 2423 898 2458 910
rect 2458 898 2492 910
rect 2492 898 2527 910
rect 2527 898 2561 910
rect 2561 898 2596 910
rect 2596 898 2630 910
rect 2630 898 2665 910
rect 2665 898 2699 910
rect 2699 898 2734 910
rect 2734 898 2768 910
rect 2768 898 2803 910
rect 2803 898 2837 910
rect 2837 898 2872 910
rect 2872 898 2906 910
rect 2906 898 2941 910
rect 2941 898 2975 910
rect 2975 898 3010 910
rect 3010 898 3044 910
rect 3044 898 3079 910
rect 3079 898 3113 910
rect 3113 898 3148 910
rect 3148 898 3182 910
rect 3182 898 3217 910
rect 3217 898 3251 910
rect 3251 898 3286 910
rect 3286 898 3320 910
rect 3320 898 3355 910
rect 3355 898 3389 910
rect 3389 898 3424 910
rect 3424 898 3458 910
rect 3458 898 3493 910
rect 3493 898 3527 910
rect 3527 898 3562 910
rect 3562 898 3596 910
rect 3596 898 3631 910
rect 3631 898 3665 910
rect 3665 898 3700 910
rect 3700 898 3734 910
rect 3734 898 3769 910
rect 3769 898 3803 910
rect 3803 898 3838 910
rect 3838 898 3872 910
rect 3872 898 3907 910
rect 3907 898 3941 910
rect 3941 898 3976 910
rect 3976 898 4010 910
rect 4010 898 4045 910
rect 4045 898 4079 910
rect 4079 898 4114 910
rect 4114 898 4148 910
rect 4148 898 4183 910
rect 4183 898 23779 978
rect 23818 970 23852 978
rect 23891 970 23925 978
rect 23964 970 23998 978
rect 24037 970 24071 978
rect 24110 970 24144 978
rect 24183 970 24217 978
rect 24256 970 24290 978
rect 24329 970 24363 978
rect 24402 970 24436 978
rect 24475 970 24509 978
rect 24548 970 24582 978
rect 24621 970 24655 978
rect 24694 970 24728 978
rect 24767 970 24801 978
rect 24840 970 24874 978
rect 24913 970 24947 978
rect 24986 970 25020 978
rect 25059 970 25093 978
rect 25132 970 25166 978
rect 25205 970 25239 978
rect 25278 970 25312 978
rect 25351 970 25385 978
rect 25424 970 25458 978
rect 25497 970 25531 978
rect 25570 970 25604 978
rect 25643 970 25677 978
rect 25716 970 25750 978
rect 25789 970 25823 978
rect 25862 970 25896 978
rect 25935 970 25969 978
rect 26008 970 26042 978
rect 26081 970 26115 978
rect 26154 970 26188 978
rect 26227 970 26261 978
rect 26300 970 26334 978
rect 26373 970 26407 978
rect 26446 970 26480 978
rect 26519 970 26553 978
rect 26592 970 26626 978
rect 26665 970 26699 978
rect 26738 970 26772 978
rect 26811 970 26845 978
rect 26884 970 26918 978
rect 26957 970 26991 978
rect 27030 970 27064 978
rect 27103 970 27137 978
rect 27176 970 27210 978
rect 27249 970 27283 978
rect 27322 970 27356 978
rect 27395 970 27429 978
rect 27468 970 27502 978
rect 27541 970 27575 978
rect 27614 970 27648 978
rect 27687 970 27721 978
rect 27760 970 27794 978
rect 27833 970 27867 978
rect 23818 898 23852 932
rect 23891 898 23925 932
rect 23964 898 23998 932
rect 24037 898 24071 932
rect 24110 898 24144 932
rect 24183 898 24217 932
rect 24256 898 24290 932
rect 24329 898 24363 932
rect 24402 898 24436 932
rect 24475 898 24509 932
rect 24548 898 24582 932
rect 24621 898 24655 932
rect 24694 898 24728 932
rect 24767 898 24801 932
rect 24840 898 24874 932
rect 24913 898 24947 932
rect 24986 898 25020 932
rect 25059 898 25093 932
rect 25132 898 25166 932
rect 25205 898 25239 932
rect 25278 898 25312 932
rect 25351 898 25385 932
rect 25424 898 25458 932
rect 25497 898 25531 932
rect 25570 898 25604 932
rect 25643 898 25677 932
rect 25716 898 25750 932
rect 25789 898 25823 932
rect 25862 898 25896 932
rect 25935 898 25969 932
rect 26008 898 26042 932
rect 26081 898 26115 932
rect 26154 898 26188 932
rect 26227 898 26261 932
rect 26300 898 26334 932
rect 26373 898 26407 932
rect 26446 898 26480 932
rect 26519 898 26553 932
rect 26592 898 26626 932
rect 26665 898 26699 932
rect 26738 898 26772 932
rect 26811 898 26845 932
rect 26884 898 26918 932
rect 26957 898 26991 932
rect 27030 898 27064 932
rect 27103 898 27137 932
rect 27176 898 27210 932
rect 27249 898 27283 932
rect 27322 898 27356 932
rect 27395 898 27429 932
rect 27468 898 27502 932
rect 27541 898 27575 932
rect 27614 898 27648 932
rect 27687 898 27721 932
rect 27760 898 27794 932
rect 27833 898 27867 932
rect 27911 930 28085 978
rect 28085 930 28089 8236
rect 165 -1487 199 -1453
rect 253 -1487 287 -1453
rect 340 -1487 374 -1453
rect 427 -1487 461 -1453
rect 514 -1487 548 -1453
rect 165 -1573 199 -1539
rect 253 -1573 287 -1539
rect 340 -1573 374 -1539
rect 427 -1573 461 -1539
rect 514 -1573 548 -1539
<< metal1 >>
rect 17183 21928 17189 21980
rect 17241 21928 17305 21980
rect 17357 21928 18040 21980
rect 18081 21921 18199 21927
rect 18133 21869 18147 21921
rect 18081 21766 18199 21869
rect 18133 21714 18147 21766
rect 18081 21708 18199 21714
rect 18368 21695 18420 21928
rect 18368 21631 18420 21643
rect 17181 21573 17187 21625
rect 17239 21573 17254 21625
rect 17306 21573 17321 21625
rect 17373 21573 17388 21625
rect 17440 21573 17454 21625
rect 17506 21573 17520 21625
rect 17572 21573 17586 21625
rect 17638 21573 17652 21625
rect 17704 21573 17718 21625
rect 17770 21573 17784 21625
rect 17836 21573 17850 21625
rect 17902 21573 17916 21625
rect 17968 21573 17982 21625
rect 18034 21573 18040 21625
rect 18368 21338 18420 21579
tri 18368 21320 18386 21338 ne
rect 18386 21320 18420 21338
tri 18420 21320 18468 21368 sw
tri 18386 21286 18420 21320 ne
rect 18420 21286 18468 21320
tri 18420 21238 18468 21286 ne
tri 18468 21238 18550 21320 sw
tri 18468 21208 18498 21238 ne
rect 18498 20199 18550 21238
rect 18498 20135 18550 20147
rect 18498 20077 18550 20083
tri 3410 18618 3531 18739 se
rect 3410 18428 3531 18618
tri 2244 18307 2365 18428 nw
tri 3410 18307 3531 18428 ne
tri 2496 18095 2577 18176 nw
tri 2921 18095 3002 18176 ne
rect 2210 11817 2244 11910
tri 2244 11817 2337 11910 sw
rect 23854 10165 23869 10217
rect 25956 10137 26074 10268
rect 3534 9876 3540 9928
rect 3592 9876 3604 9928
rect 3656 9922 18566 9928
rect 3656 9876 18514 9922
tri 18486 9848 18514 9876 ne
rect 18514 9858 18566 9870
rect 18514 9800 18566 9806
tri 2865 9590 2886 9611 sw
rect 2865 9584 2886 9590
tri 2886 9584 2892 9590 sw
rect 2865 9576 2892 9584
tri 2892 9576 2900 9584 sw
tri 18085 9576 18093 9584 se
rect 18093 9576 18124 9584
rect 18085 9532 18124 9576
rect 23854 9538 23985 9590
rect 1347 9226 28095 9232
rect 1347 9192 1425 9226
rect 1459 9192 1498 9226
rect 1532 9192 1571 9226
rect 1605 9192 1644 9226
rect 1678 9192 1717 9226
rect 1751 9192 1790 9226
rect 1824 9192 1863 9226
rect 1897 9192 1936 9226
rect 1970 9192 2009 9226
rect 2043 9192 2082 9226
rect 2116 9192 2155 9226
rect 2189 9192 2228 9226
rect 2262 9192 2301 9226
rect 2335 9192 2374 9226
rect 2408 9192 2447 9226
rect 2481 9192 2520 9226
rect 2554 9192 2593 9226
rect 2627 9192 2666 9226
rect 2700 9192 2739 9226
rect 2773 9192 2812 9226
rect 2846 9192 2885 9226
rect 2919 9192 2958 9226
rect 2992 9192 3031 9226
rect 3065 9192 3104 9226
rect 3138 9192 3177 9226
rect 3211 9192 3250 9226
rect 3284 9192 3323 9226
rect 3357 9192 3396 9226
rect 3430 9192 3469 9226
rect 3503 9192 3542 9226
rect 3576 9192 3615 9226
rect 3649 9192 3688 9226
rect 3722 9192 3761 9226
rect 3795 9192 3834 9226
rect 3868 9192 3907 9226
rect 3941 9192 3980 9226
rect 4014 9192 4053 9226
rect 4087 9192 4126 9226
rect 4160 9192 4199 9226
rect 4233 9192 4272 9226
rect 4306 9192 4345 9226
rect 4379 9192 4418 9226
rect 4452 9192 4491 9226
rect 4525 9192 4564 9226
rect 4598 9192 4637 9226
rect 4671 9192 4710 9226
rect 4744 9192 4783 9226
rect 4817 9192 4856 9226
rect 4890 9192 4929 9226
rect 4963 9192 5002 9226
rect 5036 9192 5075 9226
rect 5109 9192 5148 9226
rect 5182 9192 5221 9226
rect 5255 9192 5294 9226
rect 5328 9192 5367 9226
rect 5401 9192 5440 9226
rect 5474 9192 5513 9226
rect 1347 9154 5513 9192
rect 1347 1992 1353 9154
rect 1459 9120 1498 9154
rect 1532 9120 1571 9154
rect 1605 9120 1644 9154
rect 1678 9120 1717 9154
rect 1751 9120 1790 9154
rect 1824 9120 1863 9154
rect 1897 9120 1936 9154
rect 1970 9120 2009 9154
rect 2043 9120 2082 9154
rect 2116 9120 2155 9154
rect 2189 9120 2228 9154
rect 2262 9120 2301 9154
rect 2335 9120 2374 9154
rect 2408 9120 2447 9154
rect 2481 9120 2520 9154
rect 2554 9120 2593 9154
rect 2627 9120 2666 9154
rect 2700 9120 2739 9154
rect 2773 9120 2812 9154
rect 2846 9120 2885 9154
rect 2919 9120 2958 9154
rect 2992 9120 3031 9154
rect 3065 9120 3104 9154
rect 3138 9120 3177 9154
rect 3211 9120 3250 9154
rect 3284 9120 3323 9154
rect 3357 9120 3396 9154
rect 3430 9120 3469 9154
rect 3503 9120 3542 9154
rect 3576 9120 3615 9154
rect 3649 9120 3688 9154
rect 3722 9120 3761 9154
rect 3795 9120 3834 9154
rect 3868 9120 3907 9154
rect 3941 9120 3980 9154
rect 4014 9120 4053 9154
rect 4087 9120 4126 9154
rect 4160 9120 4199 9154
rect 4233 9120 4272 9154
rect 4306 9120 4345 9154
rect 4379 9120 4418 9154
rect 4452 9120 4491 9154
rect 4525 9120 4564 9154
rect 4598 9120 4637 9154
rect 4671 9120 4710 9154
rect 4744 9120 4783 9154
rect 4817 9120 4856 9154
rect 4890 9120 4929 9154
rect 4963 9120 5002 9154
rect 5036 9120 5075 9154
rect 5109 9120 5148 9154
rect 5182 9120 5221 9154
rect 5255 9120 5294 9154
rect 5328 9120 5367 9154
rect 5401 9120 5440 9154
rect 5474 9120 5513 9154
rect 27867 9194 28095 9226
rect 27867 9160 27911 9194
rect 27945 9160 27983 9194
rect 28017 9160 28055 9194
rect 28089 9160 28095 9194
rect 1459 9082 5585 9120
rect 1531 9048 1570 9082
rect 1604 9048 1643 9082
rect 1677 9048 1716 9082
rect 1750 9048 1789 9082
rect 1823 9048 1862 9082
rect 1896 9048 1935 9082
rect 1969 9048 2008 9082
rect 2042 9048 2081 9082
rect 2115 9048 2154 9082
rect 2188 9048 2227 9082
rect 2261 9048 2300 9082
rect 2334 9048 2373 9082
rect 2407 9048 2446 9082
rect 2480 9048 2519 9082
rect 2553 9048 2592 9082
rect 2626 9048 2665 9082
rect 2699 9048 2738 9082
rect 2772 9048 2811 9082
rect 2845 9048 2884 9082
rect 2918 9048 2957 9082
rect 2991 9048 3030 9082
rect 3064 9048 3103 9082
rect 3137 9048 3176 9082
rect 3210 9048 3249 9082
rect 3283 9048 3322 9082
rect 3356 9048 3395 9082
rect 3429 9048 3468 9082
rect 3502 9048 3541 9082
rect 3575 9048 3614 9082
rect 3648 9048 3687 9082
rect 3721 9048 3760 9082
rect 3794 9048 3833 9082
rect 3867 9048 3906 9082
rect 3940 9048 3979 9082
rect 4013 9048 4052 9082
rect 4086 9048 4125 9082
rect 4159 9048 4198 9082
rect 4232 9048 4271 9082
rect 4305 9048 4344 9082
rect 4378 9048 4417 9082
rect 4451 9048 4490 9082
rect 4524 9048 4563 9082
rect 4597 9048 4636 9082
rect 4670 9048 4709 9082
rect 4743 9048 4782 9082
rect 4816 9048 4855 9082
rect 4889 9048 4928 9082
rect 4962 9048 5001 9082
rect 5035 9048 5074 9082
rect 5108 9048 5147 9082
rect 5181 9048 5220 9082
rect 5254 9048 5293 9082
rect 5327 9048 5366 9082
rect 5400 9048 5439 9082
rect 5473 9048 5512 9082
rect 5546 9048 5585 9082
rect 27867 9114 28095 9160
rect 27867 9080 27911 9114
rect 27945 9080 27983 9114
rect 28017 9080 28055 9114
rect 28089 9080 28095 9114
rect 27867 9048 28095 9080
rect 1531 9042 28095 9048
rect 1531 2064 1537 9042
rect 27905 9034 28095 9042
tri 23290 9011 23291 9012 se
tri 18221 9004 18228 9011 sw
tri 23283 9004 23290 9011 se
rect 23290 9004 23291 9011
rect 18221 9003 18228 9004
tri 18228 9003 18229 9004 sw
rect 18221 8960 18229 9003
rect 27905 9000 27911 9034
rect 27945 9000 27983 9034
rect 28017 9000 28055 9034
rect 28089 9000 28095 9034
tri 18221 8959 18222 8960 nw
rect 27905 8954 28095 9000
rect 2905 8928 3034 8936
tri 3034 8928 3042 8936 sw
tri 23459 8928 23467 8936 se
rect 2905 8927 3042 8928
tri 3042 8927 3043 8928 sw
rect 27905 8920 27911 8954
rect 27945 8920 27983 8954
rect 28017 8920 28055 8954
rect 28089 8920 28095 8954
rect 27905 8875 28095 8920
rect 1459 2025 1537 2064
rect 1459 1992 1497 2025
rect 1347 1991 1497 1992
rect 1531 1991 1537 2025
rect 1347 1953 1537 1991
rect 1347 1919 1353 1953
rect 1387 1919 1425 1953
rect 1459 1952 1537 1953
rect 1459 1919 1497 1952
rect 1347 1918 1497 1919
rect 1531 1918 1537 1952
rect 1347 1880 1537 1918
rect 1347 1846 1353 1880
rect 1387 1846 1425 1880
rect 1459 1879 1537 1880
rect 1459 1846 1497 1879
rect 1347 1845 1497 1846
rect 1531 1845 1537 1879
rect 1347 1807 1537 1845
rect 1347 1773 1353 1807
rect 1387 1773 1425 1807
rect 1459 1806 1537 1807
rect 1459 1773 1497 1806
rect 1347 1772 1497 1773
rect 1531 1772 1537 1806
rect 1347 1734 1537 1772
rect 1347 1700 1353 1734
rect 1387 1700 1425 1734
rect 1459 1733 1537 1734
rect 1459 1700 1497 1733
rect 1347 1699 1497 1700
rect 1531 1699 1537 1733
rect 1347 1661 1537 1699
rect 1347 1627 1353 1661
rect 1387 1627 1425 1661
rect 1459 1660 1537 1661
rect 1459 1627 1497 1660
rect 1347 1626 1497 1627
rect 1531 1626 1537 1660
rect 1347 1588 1537 1626
rect 1347 1554 1353 1588
rect 1387 1554 1425 1588
rect 1459 1587 1537 1588
rect 1459 1554 1497 1587
rect 1347 1553 1497 1554
rect 1531 1553 1537 1587
rect 1347 1515 1537 1553
rect 1347 1481 1353 1515
rect 1387 1481 1425 1515
rect 1459 1514 1537 1515
rect 1459 1481 1497 1514
rect 1347 1480 1497 1481
rect 1531 1480 1537 1514
rect 1347 1442 1537 1480
rect 1347 1408 1353 1442
rect 1387 1408 1425 1442
rect 1459 1441 1537 1442
rect 1459 1408 1497 1441
rect 1347 1407 1497 1408
rect 1531 1407 1537 1441
rect 1347 1369 1537 1407
rect 1347 1335 1353 1369
rect 1387 1335 1425 1369
rect 1459 1368 1537 1369
rect 1459 1335 1497 1368
rect 1347 1334 1497 1335
rect 1531 1334 1537 1368
rect 1347 1296 1537 1334
rect 1347 1262 1353 1296
rect 1387 1262 1425 1296
rect 1459 1295 1537 1296
rect 1459 1262 1497 1295
rect 1347 1261 1497 1262
rect 1531 1261 1537 1295
rect 1795 8847 27692 8853
rect 1795 8813 1873 8847
rect 1907 8813 1946 8847
rect 1980 8813 2019 8847
rect 2053 8813 2092 8847
rect 1795 8775 2092 8813
rect 1795 5357 1801 8775
rect 1907 8741 1946 8775
rect 1980 8741 2019 8775
rect 2053 8741 2092 8775
rect 27614 8775 27692 8847
rect 27614 8741 27652 8775
rect 27686 8741 27692 8775
rect 1907 8703 2164 8741
rect 1979 8669 2018 8703
rect 2052 8669 2091 8703
rect 2125 8669 2164 8703
rect 27542 8701 27692 8741
rect 27542 8669 27580 8701
rect 1979 8667 27580 8669
rect 27614 8667 27652 8701
rect 27686 8667 27692 8701
rect 1979 8663 27692 8667
rect 1979 5429 1985 8663
tri 23172 8629 23174 8631 se
tri 23166 8623 23172 8629 se
rect 23172 8623 23174 8629
rect 27502 8629 27692 8663
rect 27502 8595 27508 8629
rect 27542 8627 27692 8629
rect 27542 8595 27580 8627
rect 27502 8593 27580 8595
rect 27614 8593 27652 8627
rect 27686 8593 27692 8627
rect 3049 8555 3052 8579
tri 3052 8555 3076 8579 nw
rect 27502 8555 27692 8593
tri 3049 8552 3052 8555 nw
tri 23341 8552 23344 8555 se
tri 23338 8549 23341 8552 se
rect 23341 8549 23344 8552
rect 3089 8547 3217 8549
tri 3217 8547 3219 8549 sw
tri 23336 8547 23338 8549 se
rect 23338 8547 23344 8549
rect 3089 8503 3223 8547
rect 3089 8497 3217 8503
tri 3217 8497 3223 8503 nw
rect 27502 8521 27508 8555
rect 27542 8553 27692 8555
rect 27542 8521 27580 8553
rect 27502 8519 27580 8521
rect 27614 8519 27652 8553
rect 27686 8519 27692 8553
rect 27502 8481 27692 8519
rect 1907 5390 1985 5429
rect 1907 5357 1945 5390
rect 1795 5356 1945 5357
rect 1979 5356 1985 5390
rect 1795 5318 1985 5356
rect 1795 5284 1801 5318
rect 1835 5284 1873 5318
rect 1907 5317 1985 5318
rect 1907 5284 1945 5317
rect 1795 5283 1945 5284
rect 1979 5283 1985 5317
rect 1795 5245 1985 5283
rect 1795 5211 1801 5245
rect 1835 5211 1873 5245
rect 1907 5244 1985 5245
rect 1907 5211 1945 5244
rect 1795 5210 1945 5211
rect 1979 5210 1985 5244
rect 1795 5172 1985 5210
rect 1795 5138 1801 5172
rect 1835 5138 1873 5172
rect 1907 5171 1985 5172
rect 1907 5138 1945 5171
rect 1795 5137 1945 5138
rect 1979 5137 1985 5171
rect 1795 5099 1985 5137
rect 1795 5065 1801 5099
rect 1835 5065 1873 5099
rect 1907 5098 1985 5099
rect 1907 5065 1945 5098
rect 1795 5064 1945 5065
rect 1979 5064 1985 5098
rect 1795 5026 1985 5064
rect 1795 4992 1801 5026
rect 1835 4992 1873 5026
rect 1907 5025 1985 5026
rect 1907 4992 1945 5025
rect 1795 4991 1945 4992
rect 1979 4991 1985 5025
rect 1795 4953 1985 4991
rect 1795 4919 1801 4953
rect 1835 4919 1873 4953
rect 1907 4952 1985 4953
rect 1907 4919 1945 4952
rect 1795 4918 1945 4919
rect 1979 4918 1985 4952
rect 1795 4880 1985 4918
rect 1795 4846 1801 4880
rect 1835 4846 1873 4880
rect 1907 4879 1985 4880
rect 1907 4846 1945 4879
rect 1795 4845 1945 4846
rect 1979 4845 1985 4879
rect 1795 4807 1985 4845
rect 1795 4773 1801 4807
rect 1835 4773 1873 4807
rect 1907 4806 1985 4807
rect 1907 4773 1945 4806
rect 1795 4772 1945 4773
rect 1979 4772 1985 4806
rect 1795 4734 1985 4772
rect 1795 4700 1801 4734
rect 1835 4700 1873 4734
rect 1907 4733 1985 4734
rect 1907 4700 1945 4733
rect 1795 4699 1945 4700
rect 1979 4699 1985 4733
rect 1795 4661 1985 4699
rect 1795 4627 1801 4661
rect 1835 4627 1873 4661
rect 1907 4660 1985 4661
rect 1907 4627 1945 4660
rect 1795 4626 1945 4627
rect 1979 4626 1985 4660
rect 1795 4588 1985 4626
rect 1795 4554 1801 4588
rect 1835 4554 1873 4588
rect 1907 4587 1985 4588
rect 1907 4554 1945 4587
rect 1795 4553 1945 4554
rect 1979 4553 1985 4587
rect 1795 4515 1985 4553
rect 1795 4481 1801 4515
rect 1835 4481 1873 4515
rect 1907 4514 1985 4515
rect 1907 4481 1945 4514
rect 1795 4480 1945 4481
rect 1979 4480 1985 4514
rect 1795 4442 1985 4480
rect 1795 4408 1801 4442
rect 1835 4408 1873 4442
rect 1907 4441 1985 4442
rect 1907 4408 1945 4441
rect 1795 4407 1945 4408
rect 1979 4407 1985 4441
rect 1795 4369 1985 4407
rect 1795 4335 1801 4369
rect 1835 4335 1873 4369
rect 1907 4368 1985 4369
rect 1907 4335 1945 4368
rect 1795 4334 1945 4335
rect 1979 4334 1985 4368
rect 1795 4296 1985 4334
rect 1795 4262 1801 4296
rect 1835 4262 1873 4296
rect 1907 4295 1985 4296
rect 1907 4262 1945 4295
rect 1795 4261 1945 4262
rect 1979 4261 1985 4295
rect 1795 4223 1985 4261
rect 1795 4189 1801 4223
rect 1835 4189 1873 4223
rect 1907 4222 1985 4223
rect 1907 4189 1945 4222
rect 1795 4188 1945 4189
rect 1979 4188 1985 4222
rect 1795 4150 1985 4188
rect 1795 4116 1801 4150
rect 1835 4116 1873 4150
rect 1907 4149 1985 4150
rect 1907 4116 1945 4149
rect 1795 4115 1945 4116
rect 1979 4115 1985 4149
rect 1795 4077 1985 4115
rect 1795 4043 1801 4077
rect 1835 4043 1873 4077
rect 1907 4076 1985 4077
rect 1907 4043 1945 4076
rect 1795 4042 1945 4043
rect 1979 4042 1985 4076
rect 1795 4004 1985 4042
rect 1795 3970 1801 4004
rect 1835 3970 1873 4004
rect 1907 4003 1985 4004
rect 1907 3970 1945 4003
rect 1795 3969 1945 3970
rect 1979 3969 1985 4003
rect 1795 3931 1985 3969
rect 1795 3897 1801 3931
rect 1835 3897 1873 3931
rect 1907 3930 1985 3931
rect 1907 3897 1945 3930
rect 1795 3896 1945 3897
rect 1979 3896 1985 3930
rect 1795 3858 1985 3896
rect 1795 3824 1801 3858
rect 1835 3824 1873 3858
rect 1907 3857 1985 3858
rect 1907 3824 1945 3857
rect 1795 3823 1945 3824
rect 1979 3823 1985 3857
rect 1795 3785 1985 3823
rect 1795 3751 1801 3785
rect 1835 3751 1873 3785
rect 1907 3784 1985 3785
rect 1907 3751 1945 3784
rect 1795 3750 1945 3751
rect 1979 3750 1985 3784
rect 1795 3712 1985 3750
rect 1795 3678 1801 3712
rect 1835 3678 1873 3712
rect 1907 3711 1985 3712
rect 1907 3678 1945 3711
rect 1795 3677 1945 3678
rect 1979 3677 1985 3711
rect 1795 3639 1985 3677
rect 1795 3605 1801 3639
rect 1835 3605 1873 3639
rect 1907 3638 1985 3639
rect 1907 3605 1945 3638
rect 1795 3604 1945 3605
rect 1979 3604 1985 3638
rect 1795 3566 1985 3604
rect 1795 3532 1801 3566
rect 1835 3532 1873 3566
rect 1907 3565 1985 3566
rect 1907 3532 1945 3565
rect 1795 3531 1945 3532
rect 1979 3531 1985 3565
rect 1795 3493 1985 3531
rect 1795 3459 1801 3493
rect 1835 3459 1873 3493
rect 1907 3492 1985 3493
rect 1907 3459 1945 3492
rect 1795 3458 1945 3459
rect 1979 3458 1985 3492
rect 1795 3420 1985 3458
rect 1795 3386 1801 3420
rect 1835 3386 1873 3420
rect 1907 3419 1985 3420
rect 1907 3386 1945 3419
rect 1795 3385 1945 3386
rect 1979 3385 1985 3419
rect 1795 3347 1985 3385
rect 1795 3313 1801 3347
rect 1835 3313 1873 3347
rect 1907 3346 1985 3347
rect 1907 3313 1945 3346
rect 1795 3312 1945 3313
rect 1979 3312 1985 3346
rect 1795 3274 1985 3312
rect 1795 3240 1801 3274
rect 1835 3240 1873 3274
rect 1907 3273 1985 3274
rect 1907 3240 1945 3273
rect 1795 3239 1945 3240
rect 1979 3239 1985 3273
rect 1795 3201 1985 3239
rect 1795 3167 1801 3201
rect 1835 3167 1873 3201
rect 1907 3200 1985 3201
rect 1907 3167 1945 3200
rect 1795 3166 1945 3167
rect 1979 3166 1985 3200
rect 1795 3128 1985 3166
rect 1795 3094 1801 3128
rect 1835 3094 1873 3128
rect 1907 3127 1985 3128
rect 1907 3094 1945 3127
rect 1795 3093 1945 3094
rect 1979 3093 1985 3127
rect 1795 3055 1985 3093
rect 1795 3021 1801 3055
rect 1835 3021 1873 3055
rect 1907 3054 1985 3055
rect 1907 3021 1945 3054
rect 1795 3020 1945 3021
rect 1979 3020 1985 3054
rect 1795 2982 1985 3020
rect 1795 2948 1801 2982
rect 1835 2948 1873 2982
rect 1907 2981 1985 2982
rect 1907 2948 1945 2981
rect 1795 2947 1945 2948
rect 1979 2947 1985 2981
rect 1795 2909 1985 2947
rect 1795 2875 1801 2909
rect 1835 2875 1873 2909
rect 1907 2908 1985 2909
rect 1907 2875 1945 2908
rect 1795 2874 1945 2875
rect 1979 2874 1985 2908
rect 1795 2836 1985 2874
rect 1795 2802 1801 2836
rect 1835 2802 1873 2836
rect 1907 2835 1985 2836
rect 1907 2802 1945 2835
rect 1795 2801 1945 2802
rect 1979 2801 1985 2835
rect 1795 2763 1985 2801
rect 1795 2729 1801 2763
rect 1835 2729 1873 2763
rect 1907 2762 1985 2763
rect 1907 2729 1945 2762
rect 1795 2728 1945 2729
rect 1979 2728 1985 2762
rect 1795 2690 1985 2728
rect 1795 2656 1801 2690
rect 1835 2656 1873 2690
rect 1907 2689 1985 2690
rect 1907 2656 1945 2689
rect 1795 2655 1945 2656
rect 1979 2655 1985 2689
rect 1795 2617 1985 2655
rect 1795 2583 1801 2617
rect 1835 2583 1873 2617
rect 1907 2616 1985 2617
rect 1907 2583 1945 2616
rect 1795 2582 1945 2583
rect 1979 2582 1985 2616
rect 1795 2544 1985 2582
rect 1795 2510 1801 2544
rect 1835 2510 1873 2544
rect 1907 2543 1985 2544
rect 1907 2510 1945 2543
rect 1795 2509 1945 2510
rect 1979 2509 1985 2543
rect 1795 2471 1985 2509
rect 1795 2437 1801 2471
rect 1835 2437 1873 2471
rect 1907 2470 1985 2471
rect 1907 2437 1945 2470
rect 1795 2436 1945 2437
rect 1979 2436 1985 2470
rect 1795 2398 1985 2436
rect 1795 2364 1801 2398
rect 1835 2364 1873 2398
rect 1907 2397 1985 2398
rect 1907 2364 1945 2397
rect 1795 2363 1945 2364
rect 1979 2363 1985 2397
rect 1795 2325 1985 2363
rect 1795 2291 1801 2325
rect 1835 2291 1873 2325
rect 1907 2324 1985 2325
rect 1907 2291 1945 2324
rect 1795 2290 1945 2291
rect 1979 2290 1985 2324
rect 1795 2252 1985 2290
rect 2181 8461 27294 8467
rect 2181 8427 2259 8461
rect 2293 8427 2332 8461
rect 2366 8427 2405 8461
rect 2439 8427 2478 8461
rect 2512 8427 2551 8461
rect 2585 8427 2624 8461
rect 2658 8427 2697 8461
rect 2731 8427 2770 8461
rect 2804 8427 2843 8461
rect 2877 8427 2916 8461
rect 2950 8427 2989 8461
rect 3023 8427 3062 8461
rect 2181 8389 3062 8427
rect 2181 5259 2187 8389
rect 2293 8355 2332 8389
rect 2366 8355 2405 8389
rect 2439 8355 2478 8389
rect 2512 8355 2551 8389
rect 2585 8355 2624 8389
rect 2658 8355 2697 8389
rect 2731 8355 2770 8389
rect 2804 8355 2843 8389
rect 2877 8355 2916 8389
rect 2950 8355 2989 8389
rect 3023 8355 3062 8389
rect 27216 8389 27294 8461
rect 27216 8355 27254 8389
rect 27288 8355 27294 8389
rect 2293 8317 3134 8355
rect 2365 8283 2404 8317
rect 2438 8283 2477 8317
rect 2511 8283 2550 8317
rect 2584 8283 2623 8317
rect 2657 8283 2696 8317
rect 2730 8283 2769 8317
rect 2803 8283 2842 8317
rect 2876 8283 2915 8317
rect 2949 8283 2988 8317
rect 3022 8283 3061 8317
rect 3095 8283 3134 8317
rect 27144 8315 27294 8355
rect 27144 8283 27182 8315
rect 2365 8281 27182 8283
rect 27216 8281 27254 8315
rect 27288 8281 27294 8315
rect 2365 8277 27294 8281
rect 2365 5331 2371 8277
rect 27104 8243 27294 8277
rect 8951 8188 8957 8240
rect 9009 8188 9021 8240
rect 9073 8188 9079 8240
rect 12171 8188 12177 8240
rect 12229 8188 12241 8240
rect 12293 8188 12299 8240
rect 15391 8188 15397 8240
rect 15449 8188 15461 8240
rect 15513 8188 15519 8240
rect 18611 8188 18617 8240
rect 18669 8188 18681 8240
rect 18733 8188 18739 8240
rect 21831 8188 21837 8240
rect 21889 8188 21901 8240
rect 21953 8188 21959 8240
rect 25051 8188 25057 8240
rect 25109 8188 25121 8240
rect 25173 8188 25179 8240
rect 26914 8236 26998 8242
rect 26914 8184 26930 8236
rect 26982 8184 26998 8236
rect 26914 8172 26998 8184
rect 6978 8083 6990 8129
tri 6978 8077 6984 8083 ne
rect 6984 8077 6990 8083
rect 7042 8077 7054 8129
rect 7106 8083 7118 8129
rect 7106 8077 7112 8083
tri 7112 8077 7118 8083 nw
rect 26914 8120 26930 8172
rect 26982 8120 26998 8172
rect 26914 8108 26998 8120
rect 26914 8056 26930 8108
rect 26982 8056 26998 8108
rect 4430 8002 4436 8054
rect 4488 8002 4500 8054
rect 4552 8002 4558 8054
rect 26914 8050 26998 8056
rect 27104 8209 27110 8243
rect 27144 8241 27294 8243
rect 27144 8209 27182 8241
rect 27104 8207 27182 8209
rect 27216 8207 27254 8241
rect 27288 8207 27294 8241
rect 27104 8169 27294 8207
rect 27104 8135 27110 8169
rect 27144 8167 27294 8169
rect 27144 8135 27182 8167
rect 27104 8133 27182 8135
rect 27216 8133 27254 8167
rect 27288 8133 27294 8167
rect 27104 8095 27294 8133
rect 27104 8061 27110 8095
rect 27144 8093 27294 8095
rect 27144 8061 27182 8093
rect 27104 8059 27182 8061
rect 27216 8059 27254 8093
rect 27288 8059 27294 8093
rect 27104 8021 27294 8059
rect 27104 7987 27110 8021
rect 27144 8019 27294 8021
rect 27144 7987 27182 8019
rect 27104 7985 27182 7987
rect 27216 7985 27254 8019
rect 27288 7985 27294 8019
rect 3298 7880 3304 7932
rect 3356 7880 3368 7932
rect 3420 7922 3426 7932
tri 3426 7922 3436 7932 sw
rect 3615 7922 3621 7974
rect 3673 7922 3685 7974
rect 3737 7922 3743 7974
rect 3420 7913 3436 7922
tri 3436 7913 3445 7922 sw
rect 3420 7912 3445 7913
tri 3445 7912 3446 7913 sw
rect 3420 7907 3446 7912
tri 3446 7907 3451 7912 sw
rect 3420 7896 3562 7907
tri 3562 7896 3573 7907 sw
tri 3764 7896 3775 7907 se
rect 3775 7896 17133 7907
rect 3420 7891 3573 7896
tri 3573 7891 3578 7896 sw
tri 3759 7891 3764 7896 se
rect 3764 7891 17133 7896
rect 3420 7880 17133 7891
rect 3315 7875 17133 7880
tri 3522 7873 3524 7875 ne
rect 3524 7873 3811 7875
tri 3811 7873 3813 7875 nw
tri 17107 7873 17109 7875 ne
rect 17109 7873 17133 7875
tri 3524 7859 3538 7873 ne
rect 3538 7859 3797 7873
tri 3797 7859 3811 7873 nw
tri 17109 7859 17123 7873 ne
rect 17123 7859 17133 7873
tri 17123 7855 17127 7859 ne
rect 17127 7855 17133 7859
rect 17185 7855 17200 7907
rect 17252 7855 17267 7907
rect 17319 7855 17333 7907
rect 17385 7855 17391 7907
rect 24210 7856 24216 7972
rect 24332 7956 26705 7972
rect 24332 7904 25661 7956
rect 25713 7904 25725 7956
rect 25777 7904 26705 7956
rect 24332 7887 26705 7904
rect 27104 7947 27294 7985
rect 27104 7913 27110 7947
rect 27144 7946 27294 7947
rect 27144 7913 27182 7946
rect 27104 7912 27182 7913
rect 27216 7912 27254 7946
rect 27288 7912 27294 7946
rect 24332 7873 24355 7887
tri 24355 7873 24369 7887 nw
rect 27104 7873 27294 7912
rect 24332 7856 24338 7873
tri 24338 7856 24355 7873 nw
rect 3371 7793 3377 7845
rect 3429 7793 3441 7845
rect 3493 7839 3499 7845
tri 3499 7839 3505 7845 sw
tri 3829 7839 3835 7845 se
rect 3835 7839 10253 7845
tri 10253 7839 10259 7845 sw
rect 27104 7839 27110 7873
rect 27144 7839 27182 7873
rect 27216 7839 27254 7873
rect 27288 7839 27294 7873
rect 3493 7823 3505 7839
tri 3505 7823 3521 7839 sw
tri 3813 7823 3829 7839 se
rect 3829 7823 10259 7839
tri 10259 7823 10275 7839 sw
rect 3493 7821 3521 7823
tri 3521 7821 3523 7823 sw
tri 3811 7821 3813 7823 se
rect 3813 7821 10275 7823
rect 3493 7814 10275 7821
tri 10275 7814 10284 7823 sw
rect 3493 7813 10284 7814
rect 3493 7793 3838 7813
tri 3838 7793 3858 7813 nw
tri 10200 7793 10220 7813 ne
rect 10220 7793 10284 7813
tri 10220 7784 10229 7793 ne
rect 10229 7784 10284 7793
tri 10229 7779 10234 7784 ne
tri 3520 7708 3534 7722 ne
rect 7137 7656 7143 7708
rect 7195 7656 7207 7708
rect 7259 7656 8501 7708
rect 8553 7656 8565 7708
rect 8617 7656 8623 7708
rect 10234 7656 10284 7784
rect 27104 7763 27294 7839
rect 27104 7729 27110 7763
rect 27144 7729 27182 7763
rect 27216 7729 27254 7763
rect 27288 7729 27294 7763
rect 27104 7690 27294 7729
tri 10284 7656 10294 7666 sw
rect 27104 7656 27110 7690
rect 27144 7656 27182 7690
rect 27216 7656 27254 7690
rect 27288 7656 27294 7690
rect 10234 7630 10294 7656
tri 10294 7630 10320 7656 sw
tri 8693 7627 8696 7630 se
rect 8696 7627 8702 7630
rect 8693 7581 8702 7627
tri 8693 7578 8696 7581 ne
rect 8696 7578 8702 7581
rect 8754 7578 8771 7630
rect 8823 7578 8839 7630
rect 8891 7627 8897 7630
tri 8897 7627 8900 7630 sw
rect 8891 7581 8900 7627
rect 10234 7627 10320 7630
tri 10320 7627 10323 7630 sw
tri 14304 7627 14307 7630 se
rect 14307 7627 14313 7630
rect 10234 7613 10332 7627
tri 10234 7583 10264 7613 ne
rect 10264 7583 10332 7613
tri 10264 7581 10266 7583 ne
rect 10266 7581 10332 7583
rect 14304 7581 14313 7627
rect 8891 7578 8897 7581
tri 8897 7578 8900 7581 nw
tri 14304 7578 14307 7581 ne
rect 14307 7578 14313 7581
rect 14365 7578 14382 7630
rect 14434 7578 14450 7630
rect 14502 7627 14508 7630
tri 14508 7627 14511 7630 sw
rect 14502 7581 14511 7627
rect 14502 7578 14508 7581
tri 14508 7578 14511 7581 nw
tri 17122 7627 17125 7630 se
rect 17125 7627 17133 7630
rect 17122 7581 17133 7627
tri 17122 7578 17125 7581 ne
rect 17125 7578 17133 7581
rect 17185 7578 17200 7630
rect 17252 7578 17267 7630
rect 17319 7578 17333 7630
rect 17385 7627 17391 7630
tri 17391 7627 17394 7630 sw
rect 17385 7581 17394 7627
rect 17385 7578 17391 7581
tri 17391 7578 17394 7581 nw
tri 20373 7627 20376 7630 se
rect 20376 7627 20382 7630
rect 20373 7581 20382 7627
tri 20373 7578 20376 7581 ne
rect 20376 7578 20382 7581
rect 20434 7578 20451 7630
rect 20503 7578 20519 7630
rect 20571 7627 20577 7630
tri 20577 7627 20580 7630 sw
rect 20571 7581 20580 7627
rect 20571 7578 20577 7581
tri 20577 7578 20580 7581 nw
tri 23767 7627 23770 7630 se
rect 23770 7627 23776 7630
rect 23767 7581 23776 7627
tri 23767 7578 23770 7581 ne
rect 23770 7578 23776 7581
rect 23828 7578 23845 7630
rect 23897 7578 23913 7630
rect 23965 7627 23971 7630
tri 23971 7627 23974 7630 sw
rect 23965 7581 23974 7627
rect 23965 7578 23971 7581
tri 23971 7578 23974 7581 nw
rect 27104 7617 27294 7656
rect 27104 7583 27110 7617
rect 27144 7583 27182 7617
rect 27216 7583 27254 7617
rect 27288 7583 27294 7617
rect 27104 7544 27294 7583
rect 27104 7510 27110 7544
rect 27144 7510 27182 7544
rect 27216 7510 27254 7544
rect 27288 7510 27294 7544
rect 3543 7424 3549 7476
rect 3601 7424 3613 7476
rect 3665 7471 3671 7476
tri 3671 7471 3676 7476 sw
rect 27104 7471 27294 7510
rect 3665 7425 4161 7471
tri 27102 7437 27104 7439 se
rect 27104 7437 27110 7471
rect 27144 7437 27182 7471
rect 27216 7437 27254 7471
rect 27288 7437 27294 7471
tri 27090 7425 27102 7437 se
rect 27102 7425 27294 7437
rect 3665 7424 3672 7425
tri 3672 7424 3673 7425 nw
tri 27089 7424 27090 7425 se
rect 27090 7424 27294 7425
tri 27080 7415 27089 7424 se
rect 27089 7415 27294 7424
rect 2475 7405 2488 7415
tri 2488 7405 2498 7415 sw
tri 27076 7411 27080 7415 se
rect 27080 7411 27294 7415
rect 2475 7398 2498 7405
tri 2498 7398 2505 7405 sw
tri 2675 7398 2682 7405 se
rect 2682 7398 2728 7405
tri 2728 7398 2735 7405 sw
rect 27076 7398 27294 7411
rect 2475 7396 2505 7398
tri 2505 7396 2507 7398 sw
tri 2673 7396 2675 7398 se
rect 2675 7396 2735 7398
tri 2735 7396 2737 7398 sw
rect 2475 7376 2507 7396
tri 2507 7376 2527 7396 sw
tri 2653 7376 2673 7396 se
rect 2673 7376 2737 7396
tri 2737 7376 2757 7396 sw
rect 2488 7371 3638 7376
tri 3638 7371 3643 7376 sw
rect 2488 7364 3643 7371
tri 3643 7364 3650 7371 sw
rect 2488 7344 3650 7364
tri 3650 7344 3670 7364 sw
rect 3927 7344 3933 7396
rect 3985 7344 3997 7396
rect 4049 7344 4055 7396
rect 27076 7364 27110 7398
rect 27144 7364 27182 7398
rect 27216 7364 27254 7398
rect 27288 7364 27294 7398
tri 2654 7325 2673 7344 ne
rect 2673 7325 2737 7344
tri 2737 7325 2756 7344 nw
tri 3615 7325 3634 7344 ne
rect 3634 7325 3670 7344
tri 3670 7325 3689 7344 sw
rect 27076 7325 27294 7364
tri 2673 7316 2682 7325 ne
rect 2682 7316 2728 7325
tri 2728 7316 2737 7325 nw
tri 3634 7316 3643 7325 ne
rect 3643 7316 3689 7325
tri 3689 7316 3698 7325 sw
tri 3643 7291 3668 7316 ne
rect 3668 7291 23776 7316
tri 3668 7285 3674 7291 ne
rect 3674 7285 23776 7291
rect 2488 7284 3630 7285
tri 3630 7284 3631 7285 sw
tri 3674 7284 3675 7285 ne
rect 3675 7284 23776 7285
rect 2488 7257 3631 7284
rect 2474 7256 3631 7257
tri 3631 7256 3659 7284 sw
tri 23750 7264 23770 7284 ne
rect 23770 7264 23776 7284
rect 23828 7264 23845 7316
rect 23897 7264 23913 7316
rect 23965 7284 24423 7316
rect 23965 7264 23971 7284
tri 23971 7264 23991 7284 nw
tri 24341 7264 24361 7284 ne
rect 24361 7264 24423 7284
tri 24361 7256 24369 7264 ne
rect 24369 7256 24423 7264
rect 2474 7253 20382 7256
rect 2474 7252 2522 7253
tri 2522 7252 2523 7253 nw
tri 3093 7252 3094 7253 ne
rect 3094 7252 3202 7253
tri 3202 7252 3203 7253 nw
tri 3607 7252 3608 7253 ne
rect 3608 7252 20382 7253
rect 2474 7231 2501 7252
tri 2501 7231 2522 7252 nw
tri 3094 7231 3115 7252 ne
rect 3115 7231 3181 7252
tri 3181 7231 3202 7252 nw
tri 3608 7231 3629 7252 ne
rect 3629 7231 20382 7252
rect 2474 7224 2494 7231
tri 2494 7224 2501 7231 nw
tri 3115 7224 3122 7231 ne
rect 3122 7224 3174 7231
tri 3174 7224 3181 7231 nw
tri 3629 7224 3636 7231 ne
rect 3636 7224 20382 7231
rect 2474 7221 2491 7224
tri 2491 7221 2494 7224 nw
tri 3122 7221 3125 7224 ne
rect 3125 7221 3171 7224
tri 3171 7221 3174 7224 nw
tri 20356 7221 20359 7224 ne
rect 20359 7221 20382 7224
rect 2474 7218 2488 7221
tri 2488 7218 2491 7221 nw
tri 20359 7218 20362 7221 ne
rect 20362 7218 20382 7221
tri 20362 7204 20376 7218 ne
rect 20376 7204 20382 7218
rect 20434 7204 20451 7256
rect 20503 7204 20519 7256
rect 20571 7252 23732 7256
tri 23732 7252 23736 7256 sw
tri 24369 7254 24371 7256 ne
rect 20571 7231 23736 7252
tri 23736 7231 23757 7252 sw
rect 20571 7224 24327 7231
rect 20571 7218 20591 7224
tri 20591 7218 20597 7224 nw
tri 23675 7218 23681 7224 ne
rect 23681 7218 24327 7224
rect 20571 7204 20577 7218
tri 20577 7204 20591 7218 nw
tri 23681 7204 23695 7218 ne
rect 23695 7204 24327 7218
tri 23695 7199 23700 7204 ne
rect 23700 7199 24327 7204
tri 24234 7196 24237 7199 ne
rect 24237 7196 24327 7199
rect 3625 7190 8702 7196
rect 3677 7164 8702 7190
rect 3677 7145 3708 7164
tri 3708 7145 3727 7164 nw
tri 8676 7145 8695 7164 ne
rect 8695 7145 8702 7164
rect 3677 7144 3707 7145
tri 3707 7144 3708 7145 nw
tri 8695 7144 8696 7145 ne
rect 8696 7144 8702 7145
rect 8754 7144 8771 7196
rect 8823 7144 8839 7196
rect 8891 7144 8897 7196
rect 8949 7144 8955 7196
rect 9007 7144 9019 7196
rect 9071 7144 9561 7196
rect 9613 7144 9625 7196
rect 9677 7144 12781 7196
rect 12833 7144 12845 7196
rect 12897 7144 14082 7196
rect 14134 7144 14146 7196
rect 14198 7163 14650 7196
rect 14198 7158 14272 7163
tri 14272 7158 14277 7163 nw
tri 14523 7158 14528 7163 ne
rect 14528 7158 14650 7163
rect 14198 7145 14259 7158
tri 14259 7145 14272 7158 nw
tri 14528 7145 14541 7158 ne
rect 14541 7145 14650 7158
rect 14198 7144 14258 7145
tri 14258 7144 14259 7145 nw
tri 14541 7144 14542 7145 ne
rect 14542 7144 14650 7145
rect 14702 7144 14714 7196
rect 14766 7144 16001 7196
rect 16053 7144 16065 7196
rect 16117 7144 19221 7196
rect 19273 7144 19285 7196
rect 19337 7144 20162 7196
rect 20214 7144 20226 7196
rect 20278 7179 20320 7196
tri 20320 7179 20337 7196 sw
tri 20604 7179 20621 7196 se
rect 20621 7179 20730 7196
rect 20278 7175 20337 7179
tri 20337 7175 20341 7179 sw
tri 20600 7175 20604 7179 se
rect 20604 7175 20730 7179
rect 20278 7144 20730 7175
rect 20782 7144 20794 7196
rect 20846 7144 22441 7196
rect 22493 7144 22505 7196
rect 22557 7144 23499 7196
rect 23551 7144 23563 7196
rect 23615 7144 23621 7196
tri 24237 7179 24254 7196 ne
rect 24254 7179 24327 7196
tri 24254 7164 24269 7179 ne
rect 24269 7164 24327 7179
tri 24269 7158 24275 7164 ne
rect 3677 7138 3697 7144
rect 3625 7134 3697 7138
tri 3697 7134 3707 7144 nw
rect 3625 7126 3677 7134
tri 3677 7114 3697 7134 nw
tri 14287 7114 14307 7134 se
rect 14307 7114 14313 7134
rect 3625 7068 3677 7074
rect 3863 7108 14313 7114
rect 3915 7082 14313 7108
rect 14365 7082 14382 7134
rect 14434 7082 14450 7134
rect 14502 7114 14508 7134
tri 14508 7114 14528 7134 sw
rect 14502 7082 24231 7114
rect 3915 7072 3955 7082
tri 3955 7072 3965 7082 nw
tri 24149 7072 24159 7082 ne
rect 24159 7072 24231 7082
rect 3915 7056 3935 7072
rect 3863 7052 3935 7056
tri 3935 7052 3955 7072 nw
tri 24159 7052 24179 7072 ne
rect 3863 7050 3933 7052
tri 3933 7050 3935 7052 nw
rect 3863 7044 3925 7050
rect 3915 7042 3925 7044
tri 3925 7042 3933 7050 nw
tri 4802 7042 4810 7050 se
rect 4810 7042 5126 7050
tri 5126 7042 5134 7050 sw
tri 10177 7042 10185 7050 se
rect 10185 7042 10584 7050
tri 10584 7042 10592 7050 sw
tri 11108 7042 11116 7050 se
rect 11116 7042 11515 7050
tri 11515 7042 11523 7050 sw
tri 16661 7042 16669 7050 se
rect 16669 7042 17069 7050
tri 17069 7042 17077 7050 sw
tri 17591 7042 17599 7050 se
rect 17599 7042 17999 7050
tri 17999 7042 18007 7050 sw
tri 23230 7042 23238 7050 se
rect 23238 7042 23552 7050
tri 23552 7042 23560 7050 sw
rect 3915 7033 3916 7042
tri 3916 7033 3925 7042 nw
tri 3915 7032 3916 7033 nw
rect 3863 6986 3915 6992
rect 4765 6963 5170 7042
tri 4765 6960 4768 6963 ne
rect 4768 6962 5170 6963
rect 4768 6960 5168 6962
tri 5168 6960 5170 6962 nw
rect 10141 6962 10592 7042
rect 11072 6962 11523 7042
rect 16626 6962 17137 7042
rect 17556 6962 18067 7042
rect 23230 6962 23596 7042
tri 10141 6960 10143 6962 ne
rect 10143 6960 10626 6962
tri 10626 6960 10628 6962 nw
tri 11072 6960 11074 6962 ne
rect 11074 6960 11557 6962
tri 11557 6960 11559 6962 nw
tri 16626 6960 16628 6962 ne
rect 16628 6960 17111 6962
tri 17111 6960 17113 6962 nw
tri 17556 6960 17558 6962 ne
rect 17558 6960 18041 6962
tri 18041 6960 18043 6962 nw
tri 23194 6960 23196 6962 ne
rect 23196 6960 23594 6962
tri 23594 6960 23596 6962 nw
tri 4768 6936 4792 6960 ne
rect 4792 6936 5134 6960
tri 3654 6926 3664 6936 ne
rect 3664 6926 3707 6936
tri 4792 6926 4802 6936 ne
rect 4802 6926 5134 6936
tri 5134 6926 5168 6960 nw
tri 10143 6926 10177 6960 ne
rect 10177 6926 10592 6960
tri 10592 6926 10626 6960 nw
tri 11074 6926 11108 6960 ne
rect 11108 6926 11523 6960
tri 11523 6926 11557 6960 nw
tri 16628 6926 16662 6960 ne
rect 16662 6926 17077 6960
tri 17077 6926 17111 6960 nw
tri 17558 6926 17592 6960 ne
rect 17592 6926 18007 6960
tri 18007 6926 18041 6960 nw
tri 23196 6926 23230 6960 ne
rect 23230 6926 23560 6960
tri 23560 6926 23594 6960 nw
tri 3664 6918 3672 6926 ne
rect 3672 6918 3707 6926
tri 4802 6918 4810 6926 ne
rect 4810 6918 5126 6926
tri 5126 6918 5134 6926 nw
tri 10177 6918 10185 6926 ne
rect 10185 6918 10584 6926
tri 10584 6918 10592 6926 nw
tri 11108 6918 11116 6926 ne
rect 11116 6918 11515 6926
tri 11515 6918 11523 6926 nw
tri 16662 6918 16670 6926 ne
rect 16670 6918 17069 6926
tri 17069 6918 17077 6926 nw
tri 17592 6918 17600 6926 ne
rect 17600 6918 17999 6926
tri 17999 6918 18007 6926 nw
tri 23230 6918 23238 6926 ne
rect 23238 6918 23552 6926
tri 23552 6918 23560 6926 nw
tri 3672 6907 3683 6918 ne
rect 3683 6907 3707 6918
rect 24179 6907 24231 7072
tri 3683 6887 3703 6907 ne
rect 3703 6887 3707 6907
tri 3703 6883 3707 6887 ne
tri 2488 6707 2498 6717 sw
rect 2488 6675 2498 6707
tri 2498 6675 2530 6707 sw
rect 2488 6668 2530 6675
tri 2530 6668 2537 6675 sw
tri 3290 6668 3297 6675 se
rect 3297 6668 3349 6675
tri 3349 6668 3356 6675 sw
rect 2488 6664 2537 6668
tri 2537 6664 2541 6668 sw
tri 3286 6664 3290 6668 se
rect 3290 6664 3356 6668
tri 3356 6664 3360 6668 sw
tri 2650 6595 2669 6614 ne
rect 2669 6595 2741 6614
tri 2741 6595 2760 6614 nw
tri 3265 6595 3284 6614 ne
rect 3284 6595 3356 6614
tri 3356 6595 3375 6614 nw
tri 2669 6582 2682 6595 ne
rect 2682 6582 2728 6595
tri 2728 6582 2741 6595 nw
tri 3284 6582 3297 6595 ne
rect 3297 6582 3343 6595
tri 3343 6582 3356 6595 nw
tri 3845 6529 3863 6547 se
tri 3118 6522 3125 6529 se
rect 3125 6522 3171 6529
tri 3171 6522 3178 6529 sw
tri 3838 6522 3845 6529 se
rect 3845 6522 3863 6529
tri 3093 6497 3118 6522 se
rect 3118 6497 3178 6522
tri 3178 6497 3203 6522 sw
tri 3813 6497 3838 6522 se
rect 3838 6497 3863 6522
tri 3841 6449 3844 6452 ne
rect 3844 6449 3863 6452
tri 3844 6447 3846 6449 ne
rect 3846 6447 3863 6449
rect 2494 6430 2531 6447
tri 2531 6430 2548 6447 nw
tri 3846 6430 3863 6447 ne
rect 2494 6415 2516 6430
tri 2516 6415 2531 6430 nw
rect 2494 6401 2498 6415
tri 2494 6397 2498 6401 ne
tri 2498 6397 2516 6415 nw
tri 3654 6123 3661 6130 ne
rect 3661 6123 3707 6130
tri 3661 6084 3700 6123 ne
rect 3700 6084 3707 6123
tri 3700 6077 3707 6084 ne
tri 16636 5977 16669 6010 se
rect 16669 5977 17068 6010
tri 17068 5977 17101 6010 sw
tri 16632 5973 16636 5977 se
rect 16636 5973 17101 5977
tri 17101 5973 17105 5977 sw
tri 2488 5904 2505 5921 sw
rect 2488 5868 2505 5904
tri 2505 5868 2541 5904 sw
tri 3507 5868 3543 5904 se
rect 16632 5867 17105 5973
tri 16632 5865 16634 5867 ne
rect 16634 5865 17103 5867
tri 17103 5865 17105 5867 nw
tri 16634 5831 16668 5865 ne
rect 16668 5831 17069 5865
tri 17069 5831 17103 5865 nw
tri 16668 5830 16669 5831 ne
rect 16669 5830 17068 5831
tri 17068 5830 17069 5831 nw
tri 2650 5792 2676 5818 ne
rect 2676 5792 2734 5818
tri 2734 5792 2760 5818 nw
tri 3507 5792 3533 5818 ne
rect 3533 5792 3543 5818
tri 2676 5786 2682 5792 ne
rect 2682 5786 2728 5792
tri 2728 5786 2734 5792 nw
tri 3533 5786 3539 5792 ne
rect 3539 5786 3543 5792
tri 3539 5782 3543 5786 ne
tri 3111 5719 3125 5733 se
rect 3125 5719 3171 5733
tri 3171 5719 3185 5733 sw
tri 3093 5701 3111 5719 se
rect 3111 5701 3185 5719
tri 3185 5701 3203 5719 sw
rect 2503 5646 2551 5651
tri 2551 5646 2556 5651 nw
tri 3406 5646 3411 5651 ne
rect 3411 5646 3459 5651
rect 2503 5612 2517 5646
tri 2517 5612 2551 5646 nw
tri 3411 5612 3445 5646 ne
rect 3445 5612 3459 5646
tri 2503 5598 2517 5612 nw
tri 3445 5598 3459 5612 ne
tri 4329 5477 4349 5497 ne
rect 4401 5466 4414 5497
tri 4414 5466 4445 5497 nw
tri 23748 5466 23779 5497 ne
rect 23779 5466 23783 5497
rect 4401 5462 4410 5466
tri 4410 5462 4414 5466 nw
tri 23779 5462 23783 5466 ne
rect 4401 5454 4402 5462
tri 4402 5454 4410 5462 nw
tri 3706 5453 3707 5454 se
tri 4401 5453 4402 5454 nw
tri 3680 5427 3706 5453 se
rect 3706 5427 3707 5453
tri 3667 5414 3680 5427 se
rect 3680 5414 3707 5427
rect 2293 5292 2371 5331
rect 2293 5259 2331 5292
rect 2181 5258 2331 5259
rect 2365 5258 2371 5292
rect 2181 5220 2371 5258
rect 2181 5186 2187 5220
rect 2221 5186 2259 5220
rect 2293 5219 2371 5220
rect 2293 5186 2331 5219
rect 2181 5185 2331 5186
rect 2365 5185 2371 5219
rect 2181 5147 2371 5185
rect 2181 5113 2187 5147
rect 2221 5113 2259 5147
rect 2293 5146 2371 5147
rect 2293 5113 2331 5146
rect 2181 5112 2331 5113
rect 2365 5112 2371 5146
rect 3707 5160 3910 5166
rect 2181 5074 2371 5112
tri 3599 5101 3625 5127 se
tri 3585 5087 3599 5101 se
rect 3599 5087 3625 5101
rect 3759 5108 3858 5160
rect 3707 5096 3910 5108
rect 2181 5040 2187 5074
rect 2221 5040 2259 5074
rect 2293 5073 2371 5074
rect 2293 5040 2331 5073
rect 2181 5039 2331 5040
rect 2365 5039 2371 5073
rect 2181 5001 2371 5039
rect 3759 5044 3858 5096
rect 3707 5038 3910 5044
tri 23761 5038 23783 5060 se
rect 23783 5038 23793 5060
tri 23760 5037 23761 5038 se
rect 23761 5037 23793 5038
rect 2181 4967 2187 5001
rect 2221 4967 2259 5001
rect 2293 5000 2371 5001
rect 2293 4967 2331 5000
rect 2181 4966 2331 4967
rect 2365 4966 2371 5000
rect 2503 5028 2534 5037
tri 2534 5028 2543 5037 nw
tri 2646 5028 2655 5037 ne
rect 2655 5028 2682 5037
rect 2503 5001 2507 5028
tri 2507 5001 2534 5028 nw
tri 2655 5001 2682 5028 ne
rect 2728 5035 2762 5037
tri 2762 5035 2764 5037 nw
tri 3601 5035 3603 5037 ne
rect 3603 5035 3625 5037
tri 23758 5035 23760 5037 se
rect 23760 5035 23793 5037
rect 2728 5028 2755 5035
tri 2755 5028 2762 5035 nw
tri 3603 5028 3610 5035 ne
rect 3610 5028 3625 5035
tri 2728 5001 2755 5028 nw
tri 3610 5013 3625 5028 ne
tri 2503 4997 2507 5001 nw
rect 2181 4928 2371 4966
rect 2181 4894 2187 4928
rect 2221 4894 2259 4928
rect 2293 4927 2371 4928
rect 2293 4894 2331 4927
rect 2181 4893 2331 4894
rect 2365 4893 2371 4927
rect 2181 4855 2371 4893
rect 2181 4821 2187 4855
rect 2221 4821 2259 4855
rect 2293 4854 2371 4855
rect 2293 4821 2331 4854
rect 2181 4820 2331 4821
rect 2365 4820 2371 4854
rect 3543 4961 3867 4967
rect 3595 4909 3867 4961
rect 3543 4897 3867 4909
rect 3595 4845 3867 4897
rect 3543 4839 3867 4845
rect 2181 4782 2371 4820
rect 2181 4748 2187 4782
rect 2221 4748 2259 4782
rect 2293 4781 2371 4782
rect 2293 4748 2331 4781
rect 2181 4747 2331 4748
rect 2365 4747 2371 4781
rect 2181 4709 2371 4747
rect 2181 4675 2187 4709
rect 2221 4675 2259 4709
rect 2293 4708 2371 4709
rect 2293 4675 2331 4708
rect 2181 4674 2331 4675
rect 2365 4674 2371 4708
rect 2181 4636 2371 4674
tri 4322 4663 4332 4673 ne
rect 4332 4663 4418 4673
tri 4418 4663 4428 4673 nw
tri 4332 4646 4349 4663 ne
rect 4349 4646 4401 4663
tri 4401 4646 4418 4663 nw
rect 2181 4602 2187 4636
rect 2221 4602 2259 4636
rect 2293 4635 2371 4636
rect 2293 4602 2331 4635
rect 2181 4601 2331 4602
rect 2365 4601 2371 4635
rect 2181 4563 2371 4601
rect 2181 4529 2187 4563
rect 2221 4529 2259 4563
rect 2293 4562 2371 4563
rect 2293 4529 2331 4562
rect 2181 4528 2331 4529
rect 2365 4528 2371 4562
rect 2181 4490 2371 4528
rect 2181 4456 2187 4490
rect 2221 4456 2259 4490
rect 2293 4489 2371 4490
rect 2293 4456 2331 4489
rect 2181 4455 2331 4456
rect 2365 4455 2371 4489
rect 2181 4417 2371 4455
rect 2181 4383 2187 4417
rect 2221 4383 2259 4417
rect 2293 4416 2371 4417
rect 2293 4383 2331 4416
rect 2181 4382 2331 4383
rect 2365 4382 2371 4416
rect 2181 4344 2371 4382
rect 2181 4310 2187 4344
rect 2221 4310 2259 4344
rect 2293 4343 2371 4344
rect 2293 4310 2331 4343
rect 2181 4309 2331 4310
rect 2365 4309 2371 4343
rect 3189 4448 3759 4454
rect 3241 4396 3707 4448
rect 3189 4384 3759 4396
rect 3241 4332 3707 4384
rect 3189 4326 3759 4332
rect 2181 4271 2371 4309
rect 2181 4237 2187 4271
rect 2221 4237 2259 4271
rect 2293 4270 2371 4271
rect 2293 4237 2331 4270
rect 2181 4236 2331 4237
rect 2365 4236 2371 4270
rect 2181 4198 2371 4236
rect 2181 4164 2187 4198
rect 2221 4164 2259 4198
rect 2293 4197 2371 4198
rect 2293 4164 2331 4197
rect 2181 4163 2331 4164
rect 2365 4163 2371 4197
rect 2181 4125 2371 4163
rect 3859 4283 3911 4289
tri 4358 4240 4359 4241 se
rect 4359 4240 4401 4241
tri 4401 4240 4402 4241 sw
rect 3859 4219 3911 4231
tri 4343 4225 4358 4240 se
rect 4358 4225 4402 4240
tri 4402 4225 4417 4240 sw
tri 14055 4225 14070 4240 se
rect 14070 4225 14122 4240
tri 14122 4225 14137 4240 sw
tri 23768 4225 23783 4240 se
rect 23783 4225 23797 4240
tri 4329 4211 4343 4225 se
rect 4343 4211 4417 4225
tri 4417 4211 4431 4225 sw
tri 14041 4211 14055 4225 se
rect 14055 4211 14137 4225
tri 14137 4211 14151 4225 sw
tri 23754 4211 23768 4225 se
rect 23768 4211 23797 4225
tri 23752 4209 23754 4211 se
rect 23754 4209 23797 4211
rect 3859 4161 3911 4167
tri 14038 4161 14042 4165 ne
rect 14042 4161 14141 4165
tri 14042 4152 14051 4161 ne
rect 14051 4152 14141 4161
tri 14141 4152 14154 4165 nw
tri 14051 4133 14070 4152 ne
rect 14070 4133 14122 4152
tri 14122 4133 14141 4152 nw
rect 2181 4091 2187 4125
rect 2221 4091 2259 4125
rect 2293 4124 2371 4125
rect 2293 4091 2331 4124
rect 2181 4090 2331 4091
rect 2365 4090 2371 4124
rect 2181 4052 2371 4090
rect 2181 4018 2187 4052
rect 2221 4018 2259 4052
rect 2293 4051 2371 4052
rect 2293 4018 2331 4051
rect 2181 4017 2331 4018
rect 2365 4017 2371 4051
rect 2181 3979 2371 4017
rect 2181 3945 2187 3979
rect 2221 3945 2259 3979
rect 2293 3978 2371 3979
rect 2293 3945 2331 3978
rect 2181 3944 2331 3945
rect 2365 3944 2371 3978
rect 3707 4093 3759 4099
tri 3759 4086 3772 4099 sw
rect 3759 4041 3866 4086
rect 3707 4035 3866 4041
rect 3707 4034 3774 4035
tri 3774 4034 3775 4035 nw
tri 3859 4034 3860 4035 ne
rect 3860 4034 3866 4035
rect 3918 4034 3930 4086
rect 3982 4034 3988 4086
rect 3707 4029 3759 4034
tri 3759 4019 3774 4034 nw
rect 3707 3971 3759 3977
rect 2181 3906 2371 3944
rect 2181 3872 2187 3906
rect 2221 3872 2259 3906
rect 2293 3905 2371 3906
rect 2293 3872 2331 3905
rect 2181 3871 2331 3872
rect 2365 3871 2371 3905
rect 2181 3833 2371 3871
rect 2181 3799 2187 3833
rect 2221 3799 2259 3833
rect 2293 3832 2371 3833
rect 2293 3799 2331 3832
rect 2181 3798 2331 3799
rect 2365 3798 2371 3832
rect 24275 3946 24327 7164
rect 24371 5351 24423 7256
rect 27076 7291 27110 7325
rect 27144 7291 27182 7325
rect 27216 7291 27254 7325
rect 27288 7291 27294 7325
rect 27076 7252 27294 7291
rect 27076 7218 27110 7252
rect 27144 7218 27182 7252
rect 27216 7218 27254 7252
rect 27288 7218 27294 7252
rect 27076 7179 27294 7218
rect 27076 7145 27110 7179
rect 27144 7145 27182 7179
rect 27216 7145 27254 7179
rect 27288 7145 27294 7179
rect 27076 7106 27294 7145
rect 27076 7072 27110 7106
rect 27144 7072 27182 7106
rect 27216 7072 27254 7106
rect 27288 7072 27294 7106
rect 27076 7033 27294 7072
rect 27076 6999 27110 7033
rect 27144 6999 27182 7033
rect 27216 6999 27254 7033
rect 27288 6999 27294 7033
rect 27076 6960 27294 6999
rect 27076 6926 27110 6960
rect 27144 6926 27182 6960
rect 27216 6926 27254 6960
rect 27288 6926 27294 6960
rect 27076 6887 27294 6926
rect 27076 6853 27110 6887
rect 27144 6853 27182 6887
rect 27216 6853 27254 6887
rect 27288 6853 27294 6887
rect 27076 6814 27294 6853
rect 27076 6780 27110 6814
rect 27144 6780 27182 6814
rect 27216 6780 27254 6814
rect 27288 6780 27294 6814
rect 27076 6741 27294 6780
rect 27076 6707 27110 6741
rect 27144 6707 27182 6741
rect 27216 6707 27254 6741
rect 27288 6707 27294 6741
rect 27076 6668 27294 6707
rect 27076 6634 27110 6668
rect 27144 6634 27182 6668
rect 27216 6634 27254 6668
rect 27288 6634 27294 6668
rect 27076 6595 27294 6634
rect 27076 6561 27110 6595
rect 27144 6561 27182 6595
rect 27216 6561 27254 6595
rect 27288 6561 27294 6595
rect 27076 6522 27294 6561
rect 27076 6488 27110 6522
rect 27144 6488 27182 6522
rect 27216 6488 27254 6522
rect 27288 6488 27294 6522
rect 27076 6449 27294 6488
rect 27076 6415 27110 6449
rect 27144 6415 27182 6449
rect 27216 6415 27254 6449
rect 27288 6415 27294 6449
rect 27076 6376 27294 6415
rect 27076 6342 27110 6376
rect 27144 6342 27182 6376
rect 27216 6342 27254 6376
rect 27288 6342 27294 6376
rect 27076 6303 27294 6342
rect 27076 6269 27110 6303
rect 27144 6269 27182 6303
rect 27216 6269 27254 6303
rect 27288 6269 27294 6303
rect 27076 6230 27294 6269
rect 27076 6196 27110 6230
rect 27144 6196 27182 6230
rect 27216 6196 27254 6230
rect 27288 6196 27294 6230
rect 27076 6157 27294 6196
rect 27076 6123 27110 6157
rect 27144 6123 27182 6157
rect 27216 6123 27254 6157
rect 27288 6123 27294 6157
rect 27076 6084 27294 6123
rect 27076 6050 27110 6084
rect 27144 6050 27182 6084
rect 27216 6050 27254 6084
rect 27288 6050 27294 6084
rect 27076 6011 27294 6050
rect 27076 5977 27110 6011
rect 27144 5977 27182 6011
rect 27216 5977 27254 6011
rect 27288 5977 27294 6011
rect 27076 5938 27294 5977
rect 27076 5904 27110 5938
rect 27144 5904 27182 5938
rect 27216 5904 27254 5938
rect 27288 5904 27294 5938
rect 27076 5865 27294 5904
rect 27076 5831 27110 5865
rect 27144 5831 27182 5865
rect 27216 5831 27254 5865
rect 27288 5831 27294 5865
rect 27076 5792 27294 5831
rect 27076 5758 27110 5792
rect 27144 5758 27182 5792
rect 27216 5758 27254 5792
rect 27288 5758 27294 5792
rect 27076 5719 27294 5758
rect 27076 5685 27110 5719
rect 27144 5685 27182 5719
rect 27216 5685 27254 5719
rect 27288 5685 27294 5719
rect 27076 5646 27294 5685
rect 27076 5612 27110 5646
rect 27144 5612 27182 5646
rect 27216 5612 27254 5646
rect 27288 5612 27294 5646
rect 27076 5573 27294 5612
rect 27076 5539 27110 5573
rect 27144 5539 27182 5573
rect 27216 5539 27254 5573
rect 27288 5539 27294 5573
rect 27076 5500 27294 5539
rect 27076 5466 27110 5500
rect 27144 5466 27182 5500
rect 27216 5466 27254 5500
rect 27288 5466 27294 5500
rect 27076 5427 27294 5466
rect 27076 5393 27110 5427
rect 27144 5393 27182 5427
rect 27216 5393 27254 5427
rect 27288 5393 27294 5427
rect 24371 5282 24423 5299
rect 24371 5212 24423 5230
rect 24371 5154 24423 5160
tri 24667 5357 24670 5360 se
rect 24670 5357 24716 5360
tri 24716 5357 24719 5360 sw
rect 24667 5351 24719 5357
rect 27076 5354 27294 5393
rect 24667 5282 24719 5299
tri 24894 5330 24897 5333 se
rect 24897 5330 24903 5333
rect 24894 5284 24903 5330
tri 24894 5281 24897 5284 ne
rect 24897 5281 24903 5284
rect 24955 5281 24970 5333
rect 25022 5281 25037 5333
rect 25089 5281 25105 5333
rect 25157 5281 25173 5333
rect 25225 5281 25241 5333
rect 25293 5281 25309 5333
rect 25361 5281 25377 5333
rect 25429 5281 25445 5333
rect 25497 5281 25513 5333
rect 25565 5281 25581 5333
rect 25633 5281 25649 5333
rect 25701 5281 25717 5333
rect 25769 5330 25775 5333
tri 25775 5330 25778 5333 sw
rect 25769 5284 25778 5330
rect 25769 5281 25775 5284
tri 25775 5281 25778 5284 nw
rect 27076 5320 27110 5354
rect 27144 5320 27182 5354
rect 27216 5320 27254 5354
rect 27288 5320 27294 5354
rect 27076 5281 27294 5320
rect 24667 5212 24719 5230
rect 27076 5247 27110 5281
rect 27144 5247 27182 5281
rect 27216 5247 27254 5281
rect 27288 5247 27294 5281
rect 27076 5208 27294 5247
tri 24719 5174 24745 5200 sw
rect 27076 5174 27110 5208
rect 27144 5174 27182 5208
rect 27216 5174 27254 5208
rect 27288 5174 27294 5208
rect 24719 5160 24745 5174
rect 24667 5155 24745 5160
tri 24745 5155 24764 5174 sw
rect 24667 5154 24764 5155
tri 24667 5135 24686 5154 ne
rect 24686 5135 24764 5154
tri 24686 5103 24718 5135 ne
rect 24718 5103 24764 5135
rect 27076 5135 27294 5174
rect 27076 5101 27110 5135
rect 27144 5101 27182 5135
rect 27216 5101 27254 5135
rect 27288 5101 27294 5135
rect 27076 5062 27294 5101
rect 27076 5028 27110 5062
rect 27144 5028 27182 5062
rect 27216 5028 27254 5062
rect 27288 5028 27294 5062
rect 27076 4989 27294 5028
rect 27076 4955 27110 4989
rect 27144 4955 27182 4989
rect 27216 4955 27254 4989
rect 27288 4955 27294 4989
rect 27076 4916 27294 4955
rect 27076 4882 27110 4916
rect 27144 4882 27182 4916
rect 27216 4882 27254 4916
rect 27288 4882 27294 4916
rect 27076 4843 27294 4882
rect 27076 4809 27110 4843
rect 27144 4809 27182 4843
rect 27216 4809 27254 4843
rect 27288 4809 27294 4843
rect 27076 4770 27294 4809
rect 27076 4736 27110 4770
rect 27144 4736 27182 4770
rect 27216 4736 27254 4770
rect 27288 4736 27294 4770
rect 27076 4697 27294 4736
rect 27076 4663 27110 4697
rect 27144 4663 27182 4697
rect 27216 4663 27254 4697
rect 27288 4663 27294 4697
rect 27076 4624 27294 4663
rect 27076 4590 27110 4624
rect 27144 4590 27182 4624
rect 27216 4590 27254 4624
rect 27288 4590 27294 4624
tri 25823 4556 25829 4562 se
rect 25829 4556 25849 4562
rect 27076 4551 27294 4590
rect 27076 4517 27110 4551
rect 27144 4517 27182 4551
rect 27216 4517 27254 4551
rect 27288 4517 27294 4551
rect 27076 4478 27294 4517
rect 27076 4444 27110 4478
rect 27144 4444 27182 4478
rect 27216 4444 27254 4478
rect 27288 4444 27294 4478
rect 27076 4405 27294 4444
rect 27076 4371 27110 4405
rect 27144 4371 27182 4405
rect 27216 4371 27254 4405
rect 27288 4371 27294 4405
rect 27076 4332 27294 4371
rect 24603 4313 24655 4319
rect 24603 4249 24655 4261
rect 24603 4154 24655 4197
rect 27076 4298 27110 4332
rect 27144 4298 27182 4332
rect 27216 4298 27254 4332
rect 27288 4298 27294 4332
rect 27076 4259 27294 4298
rect 27076 4225 27110 4259
rect 27144 4225 27182 4259
rect 27216 4225 27254 4259
rect 27288 4225 27294 4259
rect 27076 4186 27294 4225
tri 24655 4154 24677 4176 sw
rect 24603 4152 24677 4154
tri 24677 4152 24679 4154 sw
tri 26926 4152 26928 4154 se
rect 26928 4152 26932 4154
rect 24603 4149 24679 4152
tri 24679 4149 24682 4152 sw
tri 26923 4149 26926 4152 se
rect 26926 4149 26932 4152
rect 24603 4069 26932 4149
rect 27076 4152 27110 4186
rect 27144 4152 27182 4186
rect 27216 4152 27254 4186
rect 27288 4152 27294 4186
rect 27076 4113 27294 4152
rect 27076 4079 27110 4113
rect 27144 4079 27182 4113
rect 27216 4079 27254 4113
rect 27288 4079 27294 4113
tri 26901 4041 26929 4069 ne
rect 24275 3882 24327 3894
rect 24275 3824 24327 3830
rect 27076 4040 27294 4079
rect 27076 4006 27110 4040
rect 27144 4006 27182 4040
rect 27216 4006 27254 4040
rect 27288 4006 27294 4040
rect 27076 3967 27294 4006
rect 27076 3933 27110 3967
rect 27144 3933 27182 3967
rect 27216 3933 27254 3967
rect 27288 3933 27294 3967
rect 27076 3894 27294 3933
rect 27076 3860 27110 3894
rect 27144 3860 27182 3894
rect 27216 3860 27254 3894
rect 27288 3860 27294 3894
rect 2181 3760 2371 3798
rect 2181 3726 2187 3760
rect 2221 3726 2259 3760
rect 2293 3759 2371 3760
rect 2293 3726 2331 3759
rect 2181 3725 2331 3726
rect 2365 3725 2371 3759
rect 2181 3687 2371 3725
rect 2181 3653 2187 3687
rect 2221 3653 2259 3687
rect 2293 3686 2371 3687
rect 2293 3653 2331 3686
rect 2181 3652 2331 3653
rect 2365 3652 2371 3686
rect 2181 3614 2371 3652
rect 2181 3580 2187 3614
rect 2221 3580 2259 3614
rect 2293 3613 2371 3614
rect 2293 3580 2331 3613
rect 2181 3579 2331 3580
rect 2365 3579 2371 3613
rect 27076 3821 27294 3860
rect 27076 3787 27110 3821
rect 27144 3787 27182 3821
rect 27216 3787 27254 3821
rect 27288 3787 27294 3821
rect 27076 3748 27294 3787
rect 27076 3714 27110 3748
rect 27144 3714 27182 3748
rect 27216 3714 27254 3748
rect 27288 3714 27294 3748
rect 27076 3675 27294 3714
rect 27076 3641 27110 3675
rect 27144 3641 27182 3675
rect 27216 3641 27254 3675
rect 27288 3641 27294 3675
rect 27076 3602 27294 3641
tri 24076 3596 24082 3602 se
rect 2181 3541 2371 3579
rect 24082 3550 24088 3602
rect 24140 3550 24152 3602
rect 24204 3550 24210 3602
rect 27076 3568 27110 3602
rect 27144 3568 27182 3602
rect 27216 3568 27254 3602
rect 27288 3568 27294 3602
rect 2181 3507 2187 3541
rect 2221 3507 2259 3541
rect 2293 3540 2371 3541
rect 2293 3507 2331 3540
rect 2181 3506 2331 3507
rect 2365 3506 2371 3540
rect 2181 3468 2371 3506
rect 27076 3529 27294 3568
rect 2181 3434 2187 3468
rect 2221 3434 2259 3468
rect 2293 3467 2371 3468
rect 2293 3434 2331 3467
rect 2181 3433 2331 3434
rect 2365 3433 2371 3467
rect 12574 3458 12881 3504
rect 27076 3495 27110 3529
rect 27144 3495 27182 3529
rect 27216 3495 27254 3529
rect 27288 3495 27294 3529
rect 23815 3458 23843 3473
tri 23843 3458 23858 3473 nw
rect 23815 3456 23841 3458
tri 23841 3456 23843 3458 nw
rect 27076 3456 27294 3495
rect 23815 3438 23823 3456
tri 23823 3438 23841 3456 nw
rect 2181 3395 2371 3433
rect 2181 3361 2187 3395
rect 2221 3361 2259 3395
rect 2293 3394 2371 3395
rect 2293 3361 2331 3394
rect 2181 3360 2331 3361
rect 2365 3360 2371 3394
rect 3707 3386 3713 3438
rect 3765 3386 3777 3438
rect 3829 3386 3835 3438
tri 23815 3430 23823 3438 nw
rect 27076 3422 27110 3456
rect 27144 3422 27182 3456
rect 27216 3422 27254 3456
rect 27288 3422 27294 3456
rect 2181 3322 2371 3360
rect 2181 3288 2187 3322
rect 2221 3288 2259 3322
rect 2293 3321 2371 3322
rect 2293 3288 2331 3321
rect 2181 3287 2331 3288
rect 2365 3287 2371 3321
rect 2181 3249 2371 3287
rect 2181 3215 2187 3249
rect 2221 3215 2259 3249
rect 2293 3248 2371 3249
rect 2293 3215 2331 3248
rect 2181 3214 2331 3215
rect 2365 3214 2371 3248
rect 2181 3176 2371 3214
rect 2181 3142 2187 3176
rect 2221 3142 2259 3176
rect 2293 3175 2371 3176
rect 2293 3142 2331 3175
rect 2181 3141 2331 3142
rect 2365 3141 2371 3175
rect 2181 3103 2371 3141
rect 2181 3069 2187 3103
rect 2221 3069 2259 3103
rect 2293 3102 2371 3103
rect 2293 3069 2331 3102
rect 2181 3068 2331 3069
rect 2365 3068 2371 3102
rect 2181 3030 2371 3068
rect 2181 2996 2187 3030
rect 2221 2996 2259 3030
rect 2293 3029 2371 3030
rect 2293 2996 2331 3029
rect 2181 2995 2331 2996
rect 2365 2995 2371 3029
rect 2181 2957 2371 2995
rect 2181 2923 2187 2957
rect 2221 2923 2259 2957
rect 2293 2956 2371 2957
rect 2293 2923 2331 2956
rect 2181 2922 2331 2923
rect 2365 2922 2371 2956
rect 2181 2884 2371 2922
rect 2181 2850 2187 2884
rect 2221 2850 2259 2884
rect 2293 2883 2371 2884
rect 2293 2850 2331 2883
rect 2181 2849 2331 2850
rect 2365 2849 2371 2883
rect 2181 2811 2371 2849
rect 2181 2777 2187 2811
rect 2221 2777 2259 2811
rect 2293 2810 2371 2811
rect 2293 2777 2331 2810
rect 2181 2776 2331 2777
rect 2365 2776 2371 2810
rect 2181 2738 2371 2776
rect 2181 2704 2187 2738
rect 2221 2704 2259 2738
rect 2293 2737 2371 2738
rect 2293 2704 2331 2737
rect 2181 2703 2331 2704
rect 2365 2703 2371 2737
rect 2181 2665 2371 2703
rect 27076 3383 27294 3422
rect 27076 3349 27110 3383
rect 27144 3349 27182 3383
rect 27216 3349 27254 3383
rect 27288 3349 27294 3383
rect 27076 3310 27294 3349
rect 27076 3276 27110 3310
rect 27144 3276 27182 3310
rect 27216 3276 27254 3310
rect 27288 3276 27294 3310
rect 27076 3237 27294 3276
rect 2181 2631 2187 2665
rect 2221 2631 2259 2665
rect 2293 2664 2371 2665
rect 2293 2631 2331 2664
rect 2181 2630 2331 2631
rect 2365 2630 2371 2664
rect 2181 2592 2371 2630
tri 3703 2666 3707 2670 se
rect 3707 2666 3713 2670
rect 3703 2622 3713 2666
tri 3703 2618 3707 2622 ne
rect 3707 2618 3713 2622
rect 3765 2618 3777 2670
rect 3829 2668 3837 2670
tri 3837 2668 3839 2670 sw
rect 3829 2622 3839 2668
rect 3829 2618 3835 2622
tri 3835 2618 3839 2622 nw
rect 2181 2558 2187 2592
rect 2221 2558 2259 2592
rect 2293 2591 2371 2592
rect 2293 2558 2331 2591
rect 2181 2557 2331 2558
rect 2365 2557 2371 2591
rect 2181 2519 2371 2557
rect 2181 2485 2187 2519
rect 2221 2485 2259 2519
rect 2293 2518 2371 2519
rect 2293 2485 2331 2518
rect 2181 2484 2331 2485
rect 2365 2484 2371 2518
rect 2181 2451 2371 2484
rect 27076 2451 27110 3237
rect 2181 2446 27110 2451
rect 2181 2412 2187 2446
rect 2221 2412 2259 2446
rect 2293 2445 4736 2446
rect 4788 2445 4802 2446
rect 4854 2445 4868 2446
rect 4920 2445 4934 2446
rect 4986 2445 4999 2446
rect 5051 2445 5064 2446
rect 5116 2445 10192 2446
rect 10244 2445 10258 2446
rect 10310 2445 10324 2446
rect 10376 2445 10390 2446
rect 10442 2445 10455 2446
rect 10507 2445 10520 2446
rect 10572 2445 11124 2446
rect 11176 2445 11190 2446
rect 11242 2445 11256 2446
rect 11308 2445 11322 2446
rect 11374 2445 11387 2446
rect 11439 2445 11452 2446
rect 11504 2445 16677 2446
rect 16729 2445 16743 2446
rect 16795 2445 16809 2446
rect 16861 2445 16875 2446
rect 16927 2445 16940 2446
rect 16992 2445 17005 2446
rect 17057 2445 17608 2446
rect 17660 2445 17674 2446
rect 17726 2445 17740 2446
rect 17792 2445 17806 2446
rect 17858 2445 17871 2446
rect 17923 2445 17936 2446
rect 17988 2445 23161 2446
rect 23213 2445 23227 2446
rect 23279 2445 23293 2446
rect 23345 2445 23359 2446
rect 23411 2445 23424 2446
rect 23476 2445 23489 2446
rect 23541 2445 27110 2446
rect 2293 2412 2331 2445
rect 2181 2373 2331 2412
rect 26341 2411 26380 2445
rect 26414 2411 26453 2445
rect 26487 2411 26526 2445
rect 26560 2411 26599 2445
rect 26633 2411 26672 2445
rect 26706 2411 26745 2445
rect 26779 2411 26818 2445
rect 26852 2411 26891 2445
rect 26925 2411 26964 2445
rect 26998 2411 27037 2445
rect 27071 2411 27110 2445
rect 2181 2339 2187 2373
rect 2221 2339 2259 2373
rect 2181 2267 2259 2339
rect 26341 2373 27182 2411
rect 26413 2339 26452 2373
rect 26486 2339 26525 2373
rect 26559 2339 26598 2373
rect 26632 2339 26671 2373
rect 26705 2339 26744 2373
rect 26778 2339 26817 2373
rect 26851 2339 26890 2373
rect 26924 2339 26963 2373
rect 26997 2339 27036 2373
rect 27070 2339 27109 2373
rect 27143 2339 27182 2373
rect 27288 2339 27294 3237
rect 26413 2301 27294 2339
rect 26413 2267 26452 2301
rect 26486 2267 26525 2301
rect 26559 2267 26598 2301
rect 26632 2267 26671 2301
rect 26705 2267 26744 2301
rect 26778 2267 26817 2301
rect 26851 2267 26890 2301
rect 26924 2267 26963 2301
rect 26997 2267 27036 2301
rect 27070 2267 27109 2301
rect 27143 2267 27182 2301
rect 27216 2267 27294 2301
rect 2181 2266 4736 2267
rect 4788 2266 4802 2267
rect 4854 2266 4868 2267
rect 4920 2266 4934 2267
rect 4986 2266 4999 2267
rect 5051 2266 5064 2267
rect 5116 2266 10192 2267
rect 10244 2266 10258 2267
rect 10310 2266 10324 2267
rect 10376 2266 10390 2267
rect 10442 2266 10455 2267
rect 10507 2266 10520 2267
rect 10572 2266 11124 2267
rect 11176 2266 11190 2267
rect 11242 2266 11256 2267
rect 11308 2266 11322 2267
rect 11374 2266 11387 2267
rect 11439 2266 11452 2267
rect 11504 2266 16677 2267
rect 16729 2266 16743 2267
rect 16795 2266 16809 2267
rect 16861 2266 16875 2267
rect 16927 2266 16940 2267
rect 16992 2266 17005 2267
rect 17057 2266 17608 2267
rect 17660 2266 17674 2267
rect 17726 2266 17740 2267
rect 17792 2266 17806 2267
rect 17858 2266 17871 2267
rect 17923 2266 17936 2267
rect 17988 2266 23161 2267
rect 23213 2266 23227 2267
rect 23279 2266 23293 2267
rect 23345 2266 23359 2267
rect 23411 2266 23424 2267
rect 23476 2266 23489 2267
rect 23541 2266 27294 2267
rect 2181 2261 27294 2266
rect 27502 8447 27508 8481
rect 27542 8479 27692 8481
rect 27542 8447 27580 8479
rect 27502 8445 27580 8447
rect 27614 8445 27652 8479
rect 27686 8445 27692 8479
rect 27502 8407 27692 8445
rect 27502 8373 27508 8407
rect 27542 8405 27692 8407
rect 27542 8373 27580 8405
rect 27502 8371 27580 8373
rect 27614 8371 27652 8405
rect 27686 8371 27692 8405
rect 27502 8333 27692 8371
rect 27502 8299 27508 8333
rect 27542 8332 27692 8333
rect 27542 8299 27580 8332
rect 27502 8298 27580 8299
rect 27614 8298 27652 8332
rect 27686 8298 27692 8332
rect 27502 8259 27692 8298
rect 27502 8225 27508 8259
rect 27542 8225 27580 8259
rect 27614 8225 27652 8259
rect 27686 8225 27692 8259
rect 27502 8149 27692 8225
rect 27502 8115 27508 8149
rect 27542 8115 27580 8149
rect 27614 8115 27652 8149
rect 27686 8115 27692 8149
rect 27502 8076 27692 8115
rect 27502 8042 27508 8076
rect 27542 8042 27580 8076
rect 27614 8042 27652 8076
rect 27686 8042 27692 8076
rect 27502 8003 27692 8042
rect 27502 7969 27508 8003
rect 27542 7969 27580 8003
rect 27614 7969 27652 8003
rect 27686 7969 27692 8003
rect 27502 7930 27692 7969
rect 27502 7896 27508 7930
rect 27542 7896 27580 7930
rect 27614 7896 27652 7930
rect 27686 7896 27692 7930
rect 27502 7857 27692 7896
rect 27502 7823 27508 7857
rect 27542 7823 27580 7857
rect 27614 7823 27652 7857
rect 27686 7823 27692 7857
rect 27502 7784 27692 7823
rect 1795 2218 1801 2252
rect 1835 2218 1873 2252
rect 1907 2251 1985 2252
rect 1907 2218 1945 2251
rect 1795 2217 1945 2218
rect 1979 2217 1985 2251
rect 1795 2179 1985 2217
rect 1795 2145 1801 2179
rect 1835 2145 1873 2179
rect 1907 2178 1985 2179
rect 1907 2145 1945 2178
rect 1795 2144 1945 2145
rect 1979 2144 1985 2178
rect 1795 2106 1985 2144
tri 25528 2113 25529 2114 se
rect 25529 2113 26102 2114
rect 1795 2072 1801 2106
rect 1835 2072 1873 2106
rect 1907 2105 1985 2106
rect 1907 2072 1945 2105
rect 1795 2071 1945 2072
rect 1979 2071 1985 2105
rect 1795 2033 1985 2071
rect 1795 1999 1801 2033
rect 1835 1999 1873 2033
rect 1907 2032 1985 2033
rect 1907 1999 1945 2032
rect 1795 1998 1945 1999
rect 1979 1998 1985 2032
rect 1795 1960 1985 1998
rect 2415 2111 26102 2113
rect 2415 2107 25877 2111
rect 2467 2055 2493 2107
rect 2545 2059 25877 2107
rect 25929 2059 25961 2111
rect 26013 2059 26044 2111
rect 26096 2059 26102 2111
rect 2545 2055 26102 2059
rect 2415 2040 26102 2055
rect 2467 1988 2493 2040
rect 2545 2035 26102 2040
rect 2545 1988 25877 2035
rect 2415 1983 25877 1988
rect 25929 1983 25961 2035
rect 26013 1983 26044 2035
rect 26096 1983 26102 2035
rect 2415 1982 26102 1983
rect 1795 1926 1801 1960
rect 1835 1926 1873 1960
rect 1907 1959 1985 1960
rect 1907 1926 1945 1959
rect 1795 1925 1945 1926
rect 1979 1925 1985 1959
rect 1795 1887 1985 1925
rect 1795 1853 1801 1887
rect 1835 1853 1873 1887
rect 1907 1886 1985 1887
rect 1907 1853 1945 1886
rect 1795 1852 1945 1853
rect 1979 1852 1985 1886
rect 1795 1814 1985 1852
rect 1795 1780 1801 1814
rect 1835 1780 1873 1814
rect 1907 1813 1985 1814
rect 1907 1780 1945 1813
rect 1795 1779 1945 1780
rect 1979 1779 1985 1813
rect 1795 1741 1985 1779
rect 1795 1707 1801 1741
rect 1835 1707 1873 1741
rect 1907 1740 1985 1741
rect 1907 1707 1945 1740
rect 1795 1706 1945 1707
rect 1979 1706 1985 1740
rect 1795 1668 1985 1706
rect 1795 1634 1801 1668
rect 1835 1634 1873 1668
rect 1907 1667 1985 1668
rect 1907 1634 1945 1667
rect 1795 1633 1945 1634
rect 1979 1633 1985 1667
rect 2042 1741 2054 1793
rect 2106 1741 2179 1793
rect 2231 1741 20490 1793
rect 2042 1715 20490 1741
rect 2042 1663 2054 1715
rect 2106 1663 2179 1715
rect 2231 1663 20490 1715
rect 2042 1662 20490 1663
rect 1795 1595 1985 1633
rect 1795 1561 1801 1595
rect 1835 1561 1873 1595
rect 1907 1594 1985 1595
rect 1907 1561 1945 1594
rect 1795 1560 1945 1561
rect 1979 1560 1985 1594
rect 1795 1522 1985 1560
rect 1795 1488 1801 1522
rect 1835 1488 1873 1522
rect 1907 1521 1985 1522
rect 1907 1488 1945 1521
rect 1795 1487 1945 1488
rect 1979 1487 1985 1521
rect 3543 1614 3595 1615
tri 3595 1614 3596 1615 sw
rect 3543 1609 9955 1614
rect 3595 1569 9955 1609
tri 9942 1562 9949 1569 ne
rect 9949 1562 9955 1569
rect 10007 1562 10019 1614
rect 10071 1562 10077 1614
rect 3543 1545 3595 1557
rect 3543 1487 3595 1493
rect 3641 1487 3647 1539
rect 3699 1487 3711 1539
rect 3763 1531 9895 1539
tri 9895 1531 9903 1539 sw
tri 10093 1531 10101 1539 se
rect 10101 1531 14352 1539
rect 3763 1487 14352 1531
rect 14404 1487 14416 1539
rect 14468 1487 14474 1539
rect 1795 1454 1985 1487
rect 27502 1454 27508 7784
rect 1795 1449 27508 1454
rect 1795 1415 1801 1449
rect 1835 1415 1873 1449
rect 1907 1448 27508 1449
rect 1907 1415 1945 1448
rect 1795 1376 1945 1415
rect 27323 1414 27362 1448
rect 27396 1414 27435 1448
rect 27469 1414 27508 1448
rect 27323 1376 27580 1414
rect 1795 1342 1801 1376
rect 1835 1342 1873 1376
rect 1795 1270 1873 1342
rect 27395 1342 27434 1376
rect 27468 1342 27507 1376
rect 27541 1342 27580 1376
rect 27686 1342 27692 7784
rect 27395 1304 27692 1342
rect 27395 1270 27434 1304
rect 27468 1270 27507 1304
rect 27541 1270 27580 1304
rect 27614 1270 27692 1304
rect 1795 1264 27692 1270
rect 27905 8841 27911 8875
rect 27945 8841 27983 8875
rect 28017 8841 28055 8875
rect 28089 8841 28095 8875
rect 27905 8796 28095 8841
rect 27905 8762 27911 8796
rect 27945 8762 27983 8796
rect 28017 8762 28055 8796
rect 28089 8762 28095 8796
rect 27905 8717 28095 8762
rect 27905 8683 27911 8717
rect 27945 8683 27983 8717
rect 28017 8683 28055 8717
rect 28089 8683 28095 8717
rect 27905 8638 28095 8683
rect 27905 8604 27911 8638
rect 27945 8604 27983 8638
rect 28017 8604 28055 8638
rect 28089 8604 28095 8638
rect 27905 8528 28095 8604
rect 27905 8494 27911 8528
rect 27945 8494 27983 8528
rect 28017 8494 28055 8528
rect 28089 8494 28095 8528
rect 27905 8455 28095 8494
rect 27905 8421 27911 8455
rect 27945 8421 27983 8455
rect 28017 8421 28055 8455
rect 28089 8421 28095 8455
rect 27905 8382 28095 8421
rect 27905 8348 27911 8382
rect 27945 8348 27983 8382
rect 28017 8348 28055 8382
rect 28089 8348 28095 8382
rect 27905 8309 28095 8348
rect 27905 8275 27911 8309
rect 27945 8275 27983 8309
rect 28017 8275 28055 8309
rect 28089 8275 28095 8309
rect 27905 8236 28095 8275
rect 1347 1223 1537 1261
rect 1347 1189 1353 1223
rect 1387 1189 1425 1223
rect 1459 1222 1537 1223
rect 1459 1189 1497 1222
rect 1347 1188 1497 1189
rect 1531 1188 1537 1222
rect 1347 1150 1537 1188
rect 1347 1116 1353 1150
rect 1387 1116 1425 1150
rect 1459 1149 1537 1150
rect 1459 1116 1497 1149
rect 1347 1115 1497 1116
rect 1531 1115 1537 1149
rect 1347 1082 1537 1115
rect 27905 1082 27911 8236
rect 1347 1077 27911 1082
rect 1347 1043 1353 1077
rect 1387 1043 1425 1077
rect 1459 1076 27911 1077
rect 1459 1043 1497 1076
rect 1347 1004 1497 1043
rect 23779 1042 23818 1076
rect 23852 1042 23891 1076
rect 23925 1042 23964 1076
rect 23998 1042 24037 1076
rect 24071 1042 24110 1076
rect 24144 1042 24183 1076
rect 24217 1042 24256 1076
rect 24290 1042 24329 1076
rect 24363 1042 24402 1076
rect 24436 1042 24475 1076
rect 24509 1042 24548 1076
rect 24582 1042 24621 1076
rect 24655 1042 24694 1076
rect 24728 1042 24767 1076
rect 24801 1042 24840 1076
rect 24874 1042 24913 1076
rect 24947 1042 24986 1076
rect 25020 1042 25059 1076
rect 25093 1042 25132 1076
rect 25166 1042 25205 1076
rect 25239 1042 25278 1076
rect 25312 1042 25351 1076
rect 25385 1042 25424 1076
rect 25458 1042 25497 1076
rect 25531 1042 25570 1076
rect 25604 1042 25643 1076
rect 25677 1042 25716 1076
rect 25750 1042 25789 1076
rect 25823 1042 25862 1076
rect 25896 1042 25935 1076
rect 25969 1042 26008 1076
rect 26042 1042 26081 1076
rect 26115 1042 26154 1076
rect 26188 1042 26227 1076
rect 26261 1042 26300 1076
rect 26334 1042 26373 1076
rect 26407 1042 26446 1076
rect 26480 1042 26519 1076
rect 26553 1042 26592 1076
rect 26626 1042 26665 1076
rect 26699 1042 26738 1076
rect 26772 1042 26811 1076
rect 26845 1042 26884 1076
rect 26918 1042 26957 1076
rect 26991 1042 27030 1076
rect 27064 1042 27103 1076
rect 27137 1042 27176 1076
rect 27210 1042 27249 1076
rect 27283 1042 27322 1076
rect 27356 1042 27395 1076
rect 27429 1042 27468 1076
rect 27502 1042 27541 1076
rect 27575 1042 27614 1076
rect 27648 1042 27687 1076
rect 27721 1042 27760 1076
rect 27794 1042 27833 1076
rect 27867 1042 27911 1076
rect 23779 1004 27911 1042
rect 1347 970 1353 1004
rect 1387 970 1425 1004
rect 1347 898 1425 970
rect 23779 970 23818 1004
rect 23852 970 23891 1004
rect 23925 970 23964 1004
rect 23998 970 24037 1004
rect 24071 970 24110 1004
rect 24144 970 24183 1004
rect 24217 970 24256 1004
rect 24290 970 24329 1004
rect 24363 970 24402 1004
rect 24436 970 24475 1004
rect 24509 970 24548 1004
rect 24582 970 24621 1004
rect 24655 970 24694 1004
rect 24728 970 24767 1004
rect 24801 970 24840 1004
rect 24874 970 24913 1004
rect 24947 970 24986 1004
rect 25020 970 25059 1004
rect 25093 970 25132 1004
rect 25166 970 25205 1004
rect 25239 970 25278 1004
rect 25312 970 25351 1004
rect 25385 970 25424 1004
rect 25458 970 25497 1004
rect 25531 970 25570 1004
rect 25604 970 25643 1004
rect 25677 970 25716 1004
rect 25750 970 25789 1004
rect 25823 970 25862 1004
rect 25896 970 25935 1004
rect 25969 970 26008 1004
rect 26042 970 26081 1004
rect 26115 970 26154 1004
rect 26188 970 26227 1004
rect 26261 970 26300 1004
rect 26334 970 26373 1004
rect 26407 970 26446 1004
rect 26480 970 26519 1004
rect 26553 970 26592 1004
rect 26626 970 26665 1004
rect 26699 970 26738 1004
rect 26772 970 26811 1004
rect 26845 970 26884 1004
rect 26918 970 26957 1004
rect 26991 970 27030 1004
rect 27064 970 27103 1004
rect 27137 970 27176 1004
rect 27210 970 27249 1004
rect 27283 970 27322 1004
rect 27356 970 27395 1004
rect 27429 970 27468 1004
rect 27502 970 27541 1004
rect 27575 970 27614 1004
rect 27648 970 27687 1004
rect 27721 970 27760 1004
rect 27794 970 27833 1004
rect 27867 970 27911 1004
rect 23779 932 27911 970
rect 23779 898 23818 932
rect 23852 898 23891 932
rect 23925 898 23964 932
rect 23998 898 24037 932
rect 24071 898 24110 932
rect 24144 898 24183 932
rect 24217 898 24256 932
rect 24290 898 24329 932
rect 24363 898 24402 932
rect 24436 898 24475 932
rect 24509 898 24548 932
rect 24582 898 24621 932
rect 24655 898 24694 932
rect 24728 898 24767 932
rect 24801 898 24840 932
rect 24874 898 24913 932
rect 24947 898 24986 932
rect 25020 898 25059 932
rect 25093 898 25132 932
rect 25166 898 25205 932
rect 25239 898 25278 932
rect 25312 898 25351 932
rect 25385 898 25424 932
rect 25458 898 25497 932
rect 25531 898 25570 932
rect 25604 898 25643 932
rect 25677 898 25716 932
rect 25750 898 25789 932
rect 25823 898 25862 932
rect 25896 898 25935 932
rect 25969 898 26008 932
rect 26042 898 26081 932
rect 26115 898 26154 932
rect 26188 898 26227 932
rect 26261 898 26300 932
rect 26334 898 26373 932
rect 26407 898 26446 932
rect 26480 898 26519 932
rect 26553 898 26592 932
rect 26626 898 26665 932
rect 26699 898 26738 932
rect 26772 898 26811 932
rect 26845 898 26884 932
rect 26918 898 26957 932
rect 26991 898 27030 932
rect 27064 898 27103 932
rect 27137 898 27176 932
rect 27210 898 27249 932
rect 27283 898 27322 932
rect 27356 898 27395 932
rect 27429 898 27468 932
rect 27502 898 27541 932
rect 27575 898 27614 932
rect 27648 898 27687 932
rect 27721 898 27760 932
rect 27794 898 27833 932
rect 27867 930 27911 932
rect 28089 930 28095 8236
rect 27867 898 28095 930
rect 1347 892 28095 898
rect 320 -1339 326 -1287
rect 378 -1339 411 -1287
rect 463 -1339 469 -1287
rect 320 -1367 469 -1339
tri 262 -1447 320 -1389 se
rect 320 -1419 326 -1367
rect 378 -1419 411 -1367
rect 463 -1419 469 -1367
rect 665 -1323 1057 -1307
rect 665 -1375 671 -1323
rect 723 -1375 753 -1323
rect 805 -1375 835 -1323
rect 887 -1375 917 -1323
rect 969 -1375 999 -1323
rect 1051 -1375 1057 -1323
rect 320 -1447 469 -1419
tri 469 -1447 527 -1389 sw
rect 665 -1391 1057 -1375
rect 153 -1453 326 -1447
rect 153 -1487 165 -1453
rect 199 -1487 253 -1453
rect 287 -1487 326 -1453
rect 153 -1499 326 -1487
rect 378 -1499 411 -1447
rect 463 -1453 560 -1447
rect 463 -1487 514 -1453
rect 548 -1487 560 -1453
rect 463 -1499 560 -1487
rect 153 -1527 560 -1499
rect 153 -1539 326 -1527
rect 153 -1573 165 -1539
rect 199 -1573 253 -1539
rect 287 -1573 326 -1539
rect 153 -1579 326 -1573
rect 378 -1579 411 -1527
rect 463 -1539 560 -1527
rect 463 -1573 514 -1539
rect 548 -1573 560 -1539
rect 463 -1579 560 -1573
<< via1 >>
rect 17189 21928 17241 21980
rect 17305 21928 17357 21980
rect 18081 21869 18133 21921
rect 18147 21869 18199 21921
rect 18081 21714 18133 21766
rect 18147 21714 18199 21766
rect 18368 21643 18420 21695
rect 17187 21573 17239 21625
rect 17254 21573 17306 21625
rect 17321 21573 17373 21625
rect 17388 21573 17440 21625
rect 17454 21573 17506 21625
rect 17520 21573 17572 21625
rect 17586 21573 17638 21625
rect 17652 21573 17704 21625
rect 17718 21573 17770 21625
rect 17784 21573 17836 21625
rect 17850 21573 17902 21625
rect 17916 21573 17968 21625
rect 17982 21573 18034 21625
rect 18368 21579 18420 21631
rect 18498 20147 18550 20199
rect 18498 20083 18550 20135
rect 3540 9876 3592 9928
rect 3604 9876 3656 9928
rect 18514 9870 18566 9922
rect 18514 9806 18566 9858
rect 8957 8188 9009 8240
rect 9021 8188 9073 8240
rect 12177 8188 12229 8240
rect 12241 8188 12293 8240
rect 15397 8188 15449 8240
rect 15461 8188 15513 8240
rect 18617 8188 18669 8240
rect 18681 8188 18733 8240
rect 21837 8188 21889 8240
rect 21901 8188 21953 8240
rect 25057 8188 25109 8240
rect 25121 8188 25173 8240
rect 26930 8184 26982 8236
rect 6990 8077 7042 8129
rect 7054 8077 7106 8129
rect 26930 8120 26982 8172
rect 26930 8056 26982 8108
rect 4436 8002 4488 8054
rect 4500 8002 4552 8054
rect 3304 7880 3356 7932
rect 3368 7880 3420 7932
rect 3621 7922 3673 7974
rect 3685 7922 3737 7974
rect 17133 7855 17185 7907
rect 17200 7855 17252 7907
rect 17267 7855 17319 7907
rect 17333 7855 17385 7907
rect 24216 7856 24332 7972
rect 25661 7904 25713 7956
rect 25725 7904 25777 7956
rect 3377 7793 3429 7845
rect 3441 7793 3493 7845
rect 7143 7656 7195 7708
rect 7207 7656 7259 7708
rect 8501 7656 8553 7708
rect 8565 7656 8617 7708
rect 8702 7578 8754 7630
rect 8771 7578 8823 7630
rect 8839 7578 8891 7630
rect 14313 7578 14365 7630
rect 14382 7578 14434 7630
rect 14450 7578 14502 7630
rect 17133 7578 17185 7630
rect 17200 7578 17252 7630
rect 17267 7578 17319 7630
rect 17333 7578 17385 7630
rect 20382 7578 20434 7630
rect 20451 7578 20503 7630
rect 20519 7578 20571 7630
rect 23776 7578 23828 7630
rect 23845 7578 23897 7630
rect 23913 7578 23965 7630
rect 3549 7424 3601 7476
rect 3613 7424 3665 7476
rect 3933 7344 3985 7396
rect 3997 7344 4049 7396
rect 23776 7264 23828 7316
rect 23845 7264 23897 7316
rect 23913 7264 23965 7316
rect 20382 7204 20434 7256
rect 20451 7204 20503 7256
rect 20519 7204 20571 7256
rect 3625 7138 3677 7190
rect 8702 7144 8754 7196
rect 8771 7144 8823 7196
rect 8839 7144 8891 7196
rect 8955 7144 9007 7196
rect 9019 7144 9071 7196
rect 9561 7144 9613 7196
rect 9625 7144 9677 7196
rect 12781 7144 12833 7196
rect 12845 7144 12897 7196
rect 14082 7144 14134 7196
rect 14146 7144 14198 7196
rect 14650 7144 14702 7196
rect 14714 7144 14766 7196
rect 16001 7144 16053 7196
rect 16065 7144 16117 7196
rect 19221 7144 19273 7196
rect 19285 7144 19337 7196
rect 20162 7144 20214 7196
rect 20226 7144 20278 7196
rect 20730 7144 20782 7196
rect 20794 7144 20846 7196
rect 22441 7144 22493 7196
rect 22505 7144 22557 7196
rect 23499 7144 23551 7196
rect 23563 7144 23615 7196
rect 3625 7074 3677 7126
rect 3863 7056 3915 7108
rect 14313 7082 14365 7134
rect 14382 7082 14434 7134
rect 14450 7082 14502 7134
rect 3863 6992 3915 7044
rect 3707 5108 3759 5160
rect 3858 5108 3910 5160
rect 3707 5044 3759 5096
rect 3858 5044 3910 5096
rect 3543 4909 3595 4961
rect 3543 4845 3595 4897
rect 3189 4396 3241 4448
rect 3707 4396 3759 4448
rect 3189 4332 3241 4384
rect 3707 4332 3759 4384
rect 3859 4231 3911 4283
rect 3859 4167 3911 4219
rect 3707 4041 3759 4093
rect 3866 4034 3918 4086
rect 3930 4034 3982 4086
rect 3707 3977 3759 4029
rect 24371 5299 24423 5351
rect 24371 5230 24423 5282
rect 24371 5160 24423 5212
rect 24667 5299 24719 5351
rect 24667 5230 24719 5282
rect 24903 5281 24955 5333
rect 24970 5281 25022 5333
rect 25037 5281 25089 5333
rect 25105 5281 25157 5333
rect 25173 5281 25225 5333
rect 25241 5281 25293 5333
rect 25309 5281 25361 5333
rect 25377 5281 25429 5333
rect 25445 5281 25497 5333
rect 25513 5281 25565 5333
rect 25581 5281 25633 5333
rect 25649 5281 25701 5333
rect 25717 5281 25769 5333
rect 24667 5160 24719 5212
rect 24603 4261 24655 4313
rect 24603 4197 24655 4249
rect 24275 3894 24327 3946
rect 24275 3830 24327 3882
rect 24088 3550 24140 3602
rect 24152 3550 24204 3602
rect 3713 3386 3765 3438
rect 3777 3386 3829 3438
rect 3713 2618 3765 2670
rect 3777 2618 3829 2670
rect 4736 2445 4788 2446
rect 4802 2445 4854 2446
rect 4868 2445 4920 2446
rect 4934 2445 4986 2446
rect 4999 2445 5051 2446
rect 5064 2445 5116 2446
rect 10192 2445 10244 2446
rect 10258 2445 10310 2446
rect 10324 2445 10376 2446
rect 10390 2445 10442 2446
rect 10455 2445 10507 2446
rect 10520 2445 10572 2446
rect 11124 2445 11176 2446
rect 11190 2445 11242 2446
rect 11256 2445 11308 2446
rect 11322 2445 11374 2446
rect 11387 2445 11439 2446
rect 11452 2445 11504 2446
rect 16677 2445 16729 2446
rect 16743 2445 16795 2446
rect 16809 2445 16861 2446
rect 16875 2445 16927 2446
rect 16940 2445 16992 2446
rect 17005 2445 17057 2446
rect 17608 2445 17660 2446
rect 17674 2445 17726 2446
rect 17740 2445 17792 2446
rect 17806 2445 17858 2446
rect 17871 2445 17923 2446
rect 17936 2445 17988 2446
rect 23161 2445 23213 2446
rect 23227 2445 23279 2446
rect 23293 2445 23345 2446
rect 23359 2445 23411 2446
rect 23424 2445 23476 2446
rect 23489 2445 23541 2446
rect 4736 2394 4788 2445
rect 4802 2394 4854 2445
rect 4868 2394 4920 2445
rect 4934 2394 4986 2445
rect 4999 2394 5051 2445
rect 5064 2394 5116 2445
rect 10192 2394 10244 2445
rect 10258 2394 10310 2445
rect 10324 2394 10376 2445
rect 10390 2394 10442 2445
rect 10455 2394 10507 2445
rect 10520 2394 10572 2445
rect 11124 2394 11176 2445
rect 11190 2394 11242 2445
rect 11256 2394 11308 2445
rect 11322 2394 11374 2445
rect 11387 2394 11439 2445
rect 11452 2394 11504 2445
rect 16677 2394 16729 2445
rect 16743 2394 16795 2445
rect 16809 2394 16861 2445
rect 16875 2394 16927 2445
rect 16940 2394 16992 2445
rect 17005 2394 17057 2445
rect 17608 2394 17660 2445
rect 17674 2394 17726 2445
rect 17740 2394 17792 2445
rect 17806 2394 17858 2445
rect 17871 2394 17923 2445
rect 17936 2394 17988 2445
rect 23161 2394 23213 2445
rect 23227 2394 23279 2445
rect 23293 2394 23345 2445
rect 23359 2394 23411 2445
rect 23424 2394 23476 2445
rect 23489 2394 23541 2445
rect 4736 2330 4788 2382
rect 4802 2330 4854 2382
rect 4868 2330 4920 2382
rect 4934 2330 4986 2382
rect 4999 2330 5051 2382
rect 5064 2330 5116 2382
rect 10192 2330 10244 2382
rect 10258 2330 10310 2382
rect 10324 2330 10376 2382
rect 10390 2330 10442 2382
rect 10455 2330 10507 2382
rect 10520 2330 10572 2382
rect 11124 2330 11176 2382
rect 11190 2330 11242 2382
rect 11256 2330 11308 2382
rect 11322 2330 11374 2382
rect 11387 2330 11439 2382
rect 11452 2330 11504 2382
rect 16677 2330 16729 2382
rect 16743 2330 16795 2382
rect 16809 2330 16861 2382
rect 16875 2330 16927 2382
rect 16940 2330 16992 2382
rect 17005 2330 17057 2382
rect 17608 2330 17660 2382
rect 17674 2330 17726 2382
rect 17740 2330 17792 2382
rect 17806 2330 17858 2382
rect 17871 2330 17923 2382
rect 17936 2330 17988 2382
rect 23161 2330 23213 2382
rect 23227 2330 23279 2382
rect 23293 2330 23345 2382
rect 23359 2330 23411 2382
rect 23424 2330 23476 2382
rect 23489 2330 23541 2382
rect 4736 2267 4788 2318
rect 4802 2267 4854 2318
rect 4868 2267 4920 2318
rect 4934 2267 4986 2318
rect 4999 2267 5051 2318
rect 5064 2267 5116 2318
rect 10192 2267 10244 2318
rect 10258 2267 10310 2318
rect 10324 2267 10376 2318
rect 10390 2267 10442 2318
rect 10455 2267 10507 2318
rect 10520 2267 10572 2318
rect 11124 2267 11176 2318
rect 11190 2267 11242 2318
rect 11256 2267 11308 2318
rect 11322 2267 11374 2318
rect 11387 2267 11439 2318
rect 11452 2267 11504 2318
rect 16677 2267 16729 2318
rect 16743 2267 16795 2318
rect 16809 2267 16861 2318
rect 16875 2267 16927 2318
rect 16940 2267 16992 2318
rect 17005 2267 17057 2318
rect 17608 2267 17660 2318
rect 17674 2267 17726 2318
rect 17740 2267 17792 2318
rect 17806 2267 17858 2318
rect 17871 2267 17923 2318
rect 17936 2267 17988 2318
rect 23161 2267 23213 2318
rect 23227 2267 23279 2318
rect 23293 2267 23345 2318
rect 23359 2267 23411 2318
rect 23424 2267 23476 2318
rect 23489 2267 23541 2318
rect 4736 2266 4788 2267
rect 4802 2266 4854 2267
rect 4868 2266 4920 2267
rect 4934 2266 4986 2267
rect 4999 2266 5051 2267
rect 5064 2266 5116 2267
rect 10192 2266 10244 2267
rect 10258 2266 10310 2267
rect 10324 2266 10376 2267
rect 10390 2266 10442 2267
rect 10455 2266 10507 2267
rect 10520 2266 10572 2267
rect 11124 2266 11176 2267
rect 11190 2266 11242 2267
rect 11256 2266 11308 2267
rect 11322 2266 11374 2267
rect 11387 2266 11439 2267
rect 11452 2266 11504 2267
rect 16677 2266 16729 2267
rect 16743 2266 16795 2267
rect 16809 2266 16861 2267
rect 16875 2266 16927 2267
rect 16940 2266 16992 2267
rect 17005 2266 17057 2267
rect 17608 2266 17660 2267
rect 17674 2266 17726 2267
rect 17740 2266 17792 2267
rect 17806 2266 17858 2267
rect 17871 2266 17923 2267
rect 17936 2266 17988 2267
rect 23161 2266 23213 2267
rect 23227 2266 23279 2267
rect 23293 2266 23345 2267
rect 23359 2266 23411 2267
rect 23424 2266 23476 2267
rect 23489 2266 23541 2267
rect 2415 2055 2467 2107
rect 2493 2055 2545 2107
rect 25877 2059 25929 2111
rect 25961 2059 26013 2111
rect 26044 2059 26096 2111
rect 2415 1988 2467 2040
rect 2493 1988 2545 2040
rect 25877 1983 25929 2035
rect 25961 1983 26013 2035
rect 26044 1983 26096 2035
rect 2054 1741 2106 1793
rect 2179 1741 2231 1793
rect 2054 1663 2106 1715
rect 2179 1663 2231 1715
rect 3543 1557 3595 1609
rect 9955 1562 10007 1614
rect 10019 1562 10071 1614
rect 3543 1493 3595 1545
rect 3647 1487 3699 1539
rect 3711 1487 3763 1539
rect 14352 1487 14404 1539
rect 14416 1487 14468 1539
rect 326 -1339 378 -1287
rect 411 -1339 463 -1287
rect 326 -1419 378 -1367
rect 411 -1419 463 -1367
rect 671 -1375 723 -1323
rect 753 -1375 805 -1323
rect 835 -1375 887 -1323
rect 917 -1375 969 -1323
rect 999 -1375 1051 -1323
rect 326 -1453 378 -1447
rect 326 -1487 340 -1453
rect 340 -1487 374 -1453
rect 374 -1487 378 -1453
rect 326 -1499 378 -1487
rect 411 -1453 463 -1447
rect 411 -1487 427 -1453
rect 427 -1487 461 -1453
rect 461 -1487 463 -1453
rect 411 -1499 463 -1487
rect 326 -1539 378 -1527
rect 326 -1573 340 -1539
rect 340 -1573 374 -1539
rect 374 -1573 378 -1539
rect 326 -1579 378 -1573
rect 411 -1539 463 -1527
rect 411 -1573 427 -1539
rect 427 -1573 461 -1539
rect 461 -1573 463 -1539
rect 411 -1579 463 -1573
<< metal2 >>
rect 17183 21928 17189 21980
rect 17241 21928 17305 21980
rect 17357 21928 17363 21980
rect 17183 21766 17363 21928
rect 18080 21921 18430 21927
rect 18080 21869 18081 21921
rect 18133 21869 18147 21921
rect 18199 21871 18430 21921
tri 18430 21871 18486 21927 sw
rect 18199 21869 18486 21871
tri 17363 21766 17368 21771 sw
rect 18080 21766 18486 21869
rect 17183 21714 17368 21766
tri 17368 21714 17420 21766 sw
rect 18080 21714 18081 21766
rect 18133 21714 18147 21766
rect 18199 21744 18486 21766
rect 18199 21714 18277 21744
rect 17183 21695 17420 21714
tri 17420 21695 17439 21714 sw
rect 18080 21701 18277 21714
tri 18277 21701 18320 21744 nw
rect 18368 21695 18420 21701
rect 17183 21643 17439 21695
tri 17439 21643 17491 21695 sw
tri 18353 21643 18368 21658 se
rect 17183 21631 17491 21643
tri 17491 21631 17503 21643 sw
tri 18341 21631 18353 21643 se
rect 18353 21631 18420 21643
rect 17183 21625 17503 21631
tri 17503 21625 17509 21631 sw
tri 18335 21625 18341 21631 se
rect 18341 21625 18368 21631
rect 17181 21573 17187 21625
rect 17239 21573 17254 21625
rect 17306 21573 17321 21625
rect 17373 21573 17388 21625
rect 17440 21573 17454 21625
rect 17506 21573 17520 21625
rect 17572 21573 17586 21625
rect 17638 21573 17652 21625
rect 17704 21573 17718 21625
rect 17770 21573 17784 21625
rect 17836 21573 17850 21625
rect 17902 21573 17916 21625
rect 17968 21573 17982 21625
rect 18034 21579 18368 21625
rect 18034 21573 18420 21579
rect 18498 20199 18550 20205
rect 18498 20135 18550 20147
rect 18498 18946 18550 20083
tri 18498 18937 18507 18946 ne
rect 18507 18937 18550 18946
tri 18550 18937 18591 18978 sw
tri 18507 18894 18550 18937 ne
rect 18550 18894 18591 18937
tri 18550 18853 18591 18894 ne
tri 18591 18853 18675 18937 sw
tri 18591 18769 18675 18853 ne
tri 18675 18769 18759 18853 sw
tri 18675 18737 18707 18769 ne
tri 18623 18274 18707 18358 se
rect 18707 18326 18759 18769
tri 18707 18274 18759 18326 nw
tri 18539 18190 18623 18274 se
tri 18623 18190 18707 18274 nw
tri 18514 18165 18539 18190 se
rect 18539 18165 18598 18190
tri 18598 18165 18623 18190 nw
tri 2943 14360 2997 14414 ne
tri 2851 14036 2905 14090 ne
tri 2759 12896 2813 12950 ne
rect 1630 11412 1660 11416
tri 1660 11412 1664 11416 nw
tri 1630 11382 1660 11412 nw
tri 1797 11382 1827 11412 se
tri 1793 11378 1797 11382 se
rect 1797 11378 1827 11382
rect 1719 11303 1730 11326
tri 1730 11303 1753 11326 nw
tri 1719 11292 1730 11303 nw
tri 1900 11292 1911 11303 se
tri 1877 11269 1900 11292 se
rect 1900 11269 1911 11292
tri 1803 11183 1837 11217 nw
rect 3534 9876 3540 9928
rect 3592 9876 3604 9928
rect 3656 9876 3662 9928
rect 18514 9922 18566 18165
tri 18566 18133 18598 18165 nw
rect 3534 9870 3610 9876
tri 3610 9870 3616 9876 nw
rect 3534 9858 3598 9870
tri 3598 9858 3610 9870 nw
rect 18514 9858 18566 9870
tri 2957 8936 2993 8972 sw
rect 2957 8884 2993 8936
tri 2957 8848 2993 8884 nw
tri 3141 8549 3177 8585 sw
rect 3141 8497 3177 8549
tri 3141 8461 3177 8497 nw
rect 3534 8077 3586 9858
tri 3586 9846 3598 9858 nw
rect 18514 9800 18566 9806
tri 13787 9219 13790 9222 sw
rect 13787 9055 13790 9219
rect 13787 9054 13789 9055
tri 13789 9054 13790 9055 nw
rect 8951 8240 9079 8242
rect 8951 8188 8957 8240
rect 9009 8188 9021 8240
rect 9073 8188 9079 8240
rect 8951 8184 9075 8188
tri 9075 8184 9079 8188 nw
rect 12171 8240 12299 8242
rect 12171 8188 12177 8240
rect 12229 8188 12241 8240
rect 12293 8188 12299 8240
rect 12171 8184 12295 8188
tri 12295 8184 12299 8188 nw
rect 15391 8240 15519 8242
rect 15391 8188 15397 8240
rect 15449 8188 15461 8240
rect 15513 8188 15519 8240
rect 15391 8184 15515 8188
tri 15515 8184 15519 8188 nw
rect 18611 8240 18739 8242
rect 18611 8188 18617 8240
rect 18669 8188 18681 8240
rect 18733 8188 18739 8240
rect 18611 8184 18735 8188
tri 18735 8184 18739 8188 nw
rect 21831 8240 21959 8242
rect 21831 8188 21837 8240
rect 21889 8188 21901 8240
rect 21953 8188 21959 8240
rect 21831 8184 21955 8188
tri 21955 8184 21959 8188 nw
rect 25051 8240 25179 8242
rect 25051 8188 25057 8240
rect 25109 8188 25121 8240
rect 25173 8188 25179 8240
rect 25051 8184 25175 8188
tri 25175 8184 25179 8188 nw
rect 26914 8236 26998 8242
rect 26914 8184 26930 8236
rect 26982 8184 26998 8236
tri 3586 8077 3588 8079 sw
rect 6984 8077 6990 8129
rect 7042 8077 7054 8129
rect 7106 8077 7112 8129
rect 3534 8056 3588 8077
tri 3588 8056 3609 8077 sw
rect 3534 8054 3609 8056
tri 3609 8054 3611 8056 sw
rect 3534 8010 3773 8054
rect 3534 8002 3603 8010
tri 3603 8002 3611 8010 nw
tri 3765 8002 3773 8010 ne
rect 4430 8002 4436 8054
rect 4488 8002 4500 8054
rect 4552 8002 4558 8054
rect 3298 7880 3304 7932
rect 3356 7880 3368 7932
rect 3420 7880 3426 7932
rect 3298 7855 3341 7880
tri 3341 7855 3366 7880 nw
tri 2309 7476 2339 7506 sw
rect 2309 7472 2339 7476
tri 2339 7472 2343 7476 sw
tri 2403 7396 2427 7420 ne
rect 2427 7396 2437 7420
tri 2427 7386 2437 7396 ne
tri 2225 7316 2228 7319 sw
rect 2225 7285 2228 7316
tri 2228 7285 2259 7316 sw
tri 2402 7204 2431 7233 ne
rect 2431 7204 2436 7233
tri 2431 7199 2436 7204 ne
tri 2135 6742 2169 6776 sw
tri 2402 6676 2416 6690 ne
rect 2416 6676 2436 6690
tri 2416 6656 2436 6676 ne
tri 3297 6675 3298 6676 se
rect 3298 6675 3338 7855
tri 3338 7852 3341 7855 nw
rect 3371 7793 3377 7845
rect 3429 7793 3441 7845
rect 3493 7793 3499 7845
tri 3413 7759 3447 7793 ne
rect 3447 7680 3499 7793
rect 3534 7760 3586 8002
tri 3586 7985 3603 8002 nw
tri 4437 7985 4454 8002 ne
rect 4454 7985 4517 8002
tri 4454 7974 4465 7985 ne
rect 3615 7922 3621 7974
rect 3673 7922 3685 7974
rect 3737 7972 3813 7974
tri 3813 7972 3815 7974 sw
rect 3737 7958 3815 7972
tri 3815 7958 3829 7972 sw
rect 3737 7922 3829 7958
tri 3774 7907 3789 7922 ne
tri 3586 7760 3621 7795 sw
rect 3662 7708 3759 7760
tri 3680 7692 3696 7708 ne
rect 3696 7692 3759 7708
tri 3499 7680 3511 7692 sw
tri 3696 7681 3707 7692 ne
rect 3447 7660 3511 7680
tri 3447 7656 3451 7660 ne
rect 3451 7656 3511 7660
tri 3451 7648 3459 7656 ne
tri 3338 6675 3349 6686 sw
rect 3297 6572 3338 6675
tri 2051 6497 2085 6531 sw
tri 2417 6411 2451 6445 ne
tri 1803 5873 1837 5907 sw
tri 2403 5873 2437 5907 se
tri 2434 5818 2437 5821 ne
tri 1719 5771 1753 5805 sw
tri 2417 5685 2451 5719 ne
tri 1635 5108 1648 5121 sw
rect 1635 5096 1648 5108
tri 1648 5096 1660 5108 sw
rect 1635 5087 1660 5096
tri 1660 5087 1669 5096 sw
tri 2417 5001 2451 5035 ne
rect 3459 4799 3511 7656
rect 3543 7424 3549 7476
rect 3601 7424 3613 7476
rect 3665 7424 3671 7476
rect 3543 7396 3601 7424
tri 3601 7396 3629 7424 nw
rect 3543 4961 3595 7396
tri 3595 7390 3601 7396 nw
rect 3543 4897 3595 4909
rect 3543 4839 3595 4845
rect 3625 7190 3677 7196
rect 3625 7126 3677 7138
tri 3459 4795 3463 4799 ne
rect 3463 4795 3511 4799
tri 3511 4795 3529 4813 sw
tri 3463 4747 3511 4795 ne
rect 3511 4747 3529 4795
tri 3511 4729 3529 4747 ne
tri 3529 4729 3595 4795 sw
tri 3529 4715 3543 4729 ne
rect 3189 4448 3241 4454
rect 3189 4384 3241 4396
rect 3189 4326 3241 4332
rect 1257 2714 2501 2758
tri 2501 2714 2545 2758 sw
rect 1257 2551 2545 2714
tri 2360 2496 2415 2551 ne
rect 1244 2394 2125 2427
tri 2125 2394 2158 2427 sw
rect 1244 2382 2158 2394
tri 2158 2382 2170 2394 sw
rect 1244 2330 2170 2382
tri 2170 2330 2222 2382 sw
rect 1244 2318 2222 2330
tri 2222 2318 2234 2330 sw
rect 1244 2314 2234 2318
tri 2234 2314 2238 2318 sw
rect 1244 2170 2238 2314
tri 1999 2123 2046 2170 ne
rect 2046 1793 2238 2170
rect 2415 2107 2545 2551
rect 2467 2055 2493 2107
rect 2415 2040 2545 2055
rect 2467 1988 2493 2040
rect 2415 1982 2545 1988
rect 2046 1741 2054 1793
rect 2106 1741 2179 1793
rect 2231 1741 2238 1793
rect 2046 1715 2238 1741
rect 2046 1663 2054 1715
rect 2106 1663 2179 1715
rect 2231 1663 2238 1715
rect 2046 1662 2238 1663
rect 3543 1609 3595 4729
rect 3543 1545 3595 1557
rect 3543 1487 3595 1493
rect 3625 1562 3677 7074
rect 3707 5284 3759 7692
rect 3707 5160 3759 5166
rect 3707 5096 3759 5108
rect 3707 4448 3759 5044
rect 3707 4384 3759 4396
rect 3707 4326 3759 4332
rect 3707 4093 3759 4099
rect 3707 4029 3759 4041
rect 3707 3468 3759 3977
rect 3789 3526 3829 7922
rect 3927 7396 3936 7398
rect 3992 7396 4016 7398
rect 3927 7344 3933 7396
rect 3992 7344 3997 7396
rect 3927 7342 3936 7344
rect 3992 7342 4016 7344
rect 4072 7342 4081 7398
rect 3863 7108 3915 7114
rect 3863 7044 3915 7056
rect 3863 6986 3915 6992
rect 3863 6430 3903 6986
tri 3903 6974 3915 6986 nw
tri 3903 6558 3915 6570 sw
rect 3858 5160 3910 6055
rect 3858 5096 3910 5108
rect 3858 5038 3910 5044
rect 3859 4283 3911 4289
rect 3859 4219 3911 4231
rect 3859 4088 3911 4167
tri 3911 4088 3950 4127 sw
tri 4430 4088 4465 4123 se
rect 4465 4088 4517 7985
tri 4517 7974 4545 8002 nw
tri 6974 7907 6984 7917 se
rect 6984 7907 7112 8077
tri 6952 7885 6974 7907 se
rect 6974 7885 7112 7907
tri 6342 7867 6360 7885 se
rect 6360 7867 7112 7885
tri 6330 7855 6342 7867 se
rect 6342 7855 7112 7867
tri 7112 7855 7124 7867 sw
tri 6329 7854 6330 7855 se
rect 6330 7854 7124 7855
rect 6329 7832 7124 7854
tri 7124 7832 7147 7855 sw
rect 6329 7810 7243 7832
tri 7243 7810 7265 7832 sw
rect 6329 7806 7265 7810
tri 6312 7656 6329 7673 se
rect 6329 7656 6481 7806
tri 6481 7780 6507 7806 nw
tri 7039 7780 7065 7806 ne
rect 7065 7780 7265 7806
tri 7065 7708 7137 7780 ne
rect 7137 7708 7265 7780
rect 8951 7708 9065 8184
tri 9065 8174 9075 8184 nw
tri 9065 7708 9111 7754 sw
rect 12171 7708 12285 8184
tri 12285 8174 12295 8184 nw
tri 14153 7754 14156 7757 se
rect 14156 7754 14686 7757
tri 14686 7754 14689 7757 sw
tri 12285 7708 12331 7754 sw
tri 14107 7708 14153 7754 se
rect 14153 7708 14689 7754
tri 14689 7708 14735 7754 sw
rect 15391 7708 15505 8184
tri 15505 8174 15515 8184 nw
rect 17127 7855 17133 7907
rect 17185 7855 17200 7907
rect 17252 7855 17267 7907
rect 17319 7855 17333 7907
rect 17385 7855 17391 7907
tri 15505 7708 15551 7754 sw
rect 7137 7656 7143 7708
rect 7195 7656 7207 7708
rect 7259 7656 7265 7708
rect 8495 7656 8501 7708
rect 8553 7656 8565 7708
rect 8617 7695 8643 7708
tri 8643 7695 8656 7708 sw
rect 8617 7656 8656 7695
tri 6286 7630 6312 7656 se
rect 6312 7630 6481 7656
tri 8568 7655 8569 7656 ne
rect 8569 7655 8656 7656
tri 6481 7630 6506 7655 sw
tri 8569 7630 8594 7655 ne
rect 8594 7630 8656 7655
tri 14076 7677 14107 7708 se
rect 14107 7677 14735 7708
rect 14076 7673 14735 7677
tri 14735 7673 14770 7708 sw
rect 14076 7630 14212 7673
tri 14212 7630 14255 7673 nw
tri 14585 7630 14628 7673 ne
rect 14628 7671 14770 7673
tri 14770 7671 14772 7673 sw
rect 14628 7630 14772 7671
tri 8594 7628 8596 7630 ne
rect 8596 7114 8656 7630
rect 8696 7578 8702 7630
rect 8754 7578 8771 7630
rect 8823 7578 8839 7630
rect 8891 7578 8897 7630
rect 8696 7196 8897 7578
rect 9555 7196 9683 7482
rect 8696 7144 8702 7196
rect 8754 7144 8771 7196
rect 8823 7144 8839 7196
rect 8891 7144 8897 7196
rect 8949 7144 8955 7196
rect 9007 7144 9019 7196
rect 9071 7144 9077 7196
rect 9555 7144 9561 7196
rect 9613 7144 9625 7196
rect 9677 7144 9683 7196
rect 12775 7196 12903 7482
rect 12775 7144 12781 7196
rect 12833 7144 12845 7196
rect 12897 7144 12903 7196
rect 14076 7196 14204 7630
tri 14204 7622 14212 7630 nw
rect 14076 7144 14082 7196
rect 14134 7144 14146 7196
rect 14198 7144 14204 7196
rect 14307 7578 14313 7630
rect 14365 7578 14382 7630
rect 14434 7578 14450 7630
rect 14502 7578 14508 7630
tri 14628 7614 14644 7630 ne
rect 8949 7134 9022 7144
tri 9022 7134 9032 7144 nw
rect 14307 7134 14508 7578
rect 14644 7196 14772 7630
rect 17127 7630 17391 7855
rect 18611 7708 18725 8184
tri 18725 8174 18735 8184 nw
tri 20233 7754 20236 7757 se
rect 20236 7754 20766 7757
tri 20766 7754 20769 7757 sw
tri 18725 7708 18771 7754 sw
tri 20187 7708 20233 7754 se
rect 20233 7708 20769 7754
tri 20769 7708 20815 7754 sw
rect 21831 7708 21945 8184
tri 21945 8174 21955 8184 nw
rect 24210 7856 24216 7972
rect 24332 7856 24338 7972
tri 24151 7757 24210 7816 se
rect 24210 7759 24338 7856
rect 24210 7757 24336 7759
tri 24336 7757 24338 7759 nw
tri 23570 7754 23573 7757 se
rect 23573 7754 24287 7757
tri 21945 7708 21991 7754 sw
tri 23524 7708 23570 7754 se
rect 23570 7708 24287 7754
tri 24287 7708 24336 7757 nw
rect 25051 7708 25165 8184
tri 25165 8174 25175 8184 nw
rect 26914 8172 26998 8184
rect 26914 8120 26930 8172
rect 26982 8120 26998 8172
rect 26914 8108 26998 8120
rect 26914 8056 26930 8108
rect 26982 8056 26998 8108
rect 26914 8050 26998 8056
tri 26914 8027 26937 8050 ne
rect 25655 7956 25783 7972
rect 25655 7904 25661 7956
rect 25713 7904 25725 7956
rect 25777 7904 25783 7956
tri 25165 7708 25211 7754 sw
rect 25655 7708 25783 7904
rect 17127 7578 17133 7630
rect 17185 7578 17200 7630
rect 17252 7578 17267 7630
rect 17319 7578 17333 7630
rect 17385 7578 17391 7630
tri 20156 7677 20187 7708 se
rect 20187 7677 20815 7708
rect 20156 7673 20815 7677
tri 20815 7673 20850 7708 sw
tri 23493 7677 23524 7708 se
rect 23524 7677 24256 7708
tri 24256 7677 24287 7708 nw
rect 23493 7673 24252 7677
tri 24252 7673 24256 7677 nw
rect 20156 7630 20292 7673
tri 20292 7630 20335 7673 nw
tri 20665 7630 20708 7673 ne
rect 20708 7671 20850 7673
tri 20850 7671 20852 7673 sw
rect 20708 7630 20852 7671
rect 14644 7144 14650 7196
rect 14702 7144 14714 7196
rect 14766 7144 14772 7196
rect 15995 7196 16123 7482
rect 15995 7144 16001 7196
rect 16053 7144 16065 7196
rect 16117 7144 16123 7196
rect 19215 7196 19343 7482
rect 19215 7144 19221 7196
rect 19273 7144 19285 7196
rect 19337 7144 19343 7196
rect 20156 7196 20284 7630
tri 20284 7622 20292 7630 nw
rect 20376 7578 20382 7630
rect 20434 7578 20451 7630
rect 20503 7578 20519 7630
rect 20571 7578 20577 7630
tri 20708 7614 20724 7630 ne
rect 20376 7256 20577 7578
rect 20376 7204 20382 7256
rect 20434 7204 20451 7256
rect 20503 7204 20519 7256
rect 20571 7204 20577 7256
rect 20156 7144 20162 7196
rect 20214 7144 20226 7196
rect 20278 7144 20284 7196
rect 20724 7196 20852 7630
rect 23493 7630 23629 7673
tri 23629 7630 23672 7673 nw
rect 20724 7144 20730 7196
rect 20782 7144 20794 7196
rect 20846 7144 20852 7196
rect 22435 7196 22563 7482
rect 22435 7144 22441 7196
rect 22493 7144 22505 7196
rect 22557 7144 22563 7196
rect 23493 7196 23621 7630
tri 23621 7622 23629 7630 nw
rect 23770 7578 23776 7630
rect 23828 7578 23845 7630
rect 23897 7578 23913 7630
rect 23965 7578 23971 7630
rect 23770 7316 23971 7578
tri 26866 7437 26937 7508 se
rect 26937 7482 26982 8050
tri 26982 8034 26998 8050 nw
tri 26937 7437 26982 7482 nw
rect 23770 7264 23776 7316
rect 23828 7264 23845 7316
rect 23897 7264 23913 7316
rect 23965 7264 23971 7316
tri 26849 7420 26866 7437 se
rect 26866 7420 26920 7437
tri 26920 7420 26937 7437 nw
rect 23493 7144 23499 7196
rect 23551 7144 23563 7196
rect 23615 7144 23621 7196
rect 26849 7151 26901 7420
tri 26901 7401 26920 7420 nw
rect 8949 7130 9018 7134
tri 9018 7130 9022 7134 nw
tri 8944 7125 8949 7130 se
rect 8949 7125 8978 7130
tri 8656 7114 8667 7125 sw
tri 8933 7114 8944 7125 se
rect 8944 7114 8978 7125
rect 8596 7090 8667 7114
tri 8667 7090 8691 7114 sw
tri 8909 7090 8933 7114 se
rect 8933 7090 8978 7114
tri 8978 7090 9018 7130 nw
rect 8596 7082 8970 7090
tri 8970 7082 8978 7090 nw
rect 14307 7082 14313 7134
rect 14365 7082 14382 7134
rect 14434 7082 14450 7134
rect 14502 7082 14508 7134
rect 8596 7081 8969 7082
tri 8969 7081 8970 7082 nw
tri 8596 7043 8634 7081 ne
rect 8634 7043 8931 7081
tri 8931 7043 8969 7081 nw
rect 24371 5351 24719 5357
rect 24423 5299 24667 5351
rect 24371 5282 24719 5299
rect 24423 5230 24667 5282
rect 24897 5281 24903 5333
rect 24955 5281 24970 5333
rect 25022 5281 25037 5333
rect 25089 5281 25105 5333
rect 25157 5281 25173 5333
rect 25225 5281 25241 5333
rect 25293 5281 25309 5333
rect 25361 5281 25377 5333
rect 25429 5281 25445 5333
rect 25497 5281 25513 5333
rect 25565 5281 25581 5333
rect 25633 5281 25649 5333
rect 25701 5281 25717 5333
rect 25769 5281 25775 5333
rect 24371 5212 24719 5230
rect 24423 5160 24667 5212
rect 24371 5154 24719 5160
tri 24762 4953 24897 5088 se
rect 21843 4755 24897 4953
tri 24797 4752 24800 4755 ne
rect 24800 4752 24897 4755
tri 24800 4655 24897 4752 ne
rect 25875 4743 26095 4752
rect 25931 4687 25957 4743
rect 26013 4687 26039 4743
rect 25875 4663 26095 4687
rect 25931 4607 25957 4663
rect 26013 4607 26039 4663
rect 25875 4583 26095 4607
rect 25931 4527 25957 4583
rect 26013 4527 26039 4583
rect 25875 4503 26095 4527
rect 25931 4447 25957 4503
rect 26013 4447 26039 4503
rect 25875 4423 26095 4447
rect 25931 4367 25957 4423
rect 26013 4367 26039 4423
rect 24603 4313 24655 4319
rect 24603 4249 24655 4261
tri 24579 4162 24603 4186 se
rect 24603 4162 24655 4197
rect 3859 4086 4517 4088
rect 3859 4034 3866 4086
rect 3918 4034 3930 4086
rect 3982 4034 4517 4086
rect 24231 4125 24655 4162
rect 24231 4099 24245 4125
tri 24245 4099 24271 4125 nw
tri 24577 4099 24603 4125 ne
rect 24603 4099 24655 4125
rect 24231 4088 24234 4099
tri 24234 4088 24245 4099 nw
tri 24231 4085 24234 4088 nw
rect 3859 4031 4517 4034
rect 24275 3949 24327 3952
tri 24327 3949 24330 3952 sw
rect 24275 3946 24330 3949
rect 24327 3894 24330 3946
rect 24275 3882 24330 3894
rect 24327 3830 24330 3882
rect 16967 3676 17272 3685
tri 3829 3526 3846 3543 sw
rect 3789 3525 3846 3526
tri 3789 3474 3840 3525 ne
rect 3840 3474 3846 3525
tri 3759 3468 3765 3474 sw
tri 3840 3468 3846 3474 ne
tri 3846 3468 3904 3526 sw
rect 3707 3450 3765 3468
tri 3765 3450 3783 3468 sw
tri 3846 3450 3864 3468 ne
rect 3707 3438 3783 3450
tri 3783 3438 3795 3450 sw
rect 3707 3386 3713 3438
rect 3765 3386 3777 3438
rect 3829 3386 3835 3438
rect 3707 2674 3759 3386
tri 3759 3350 3795 3386 nw
tri 3841 3275 3864 3298 se
rect 3864 3275 3904 3468
rect 9382 3520 9391 3576
rect 9447 3520 9481 3576
rect 9537 3520 9571 3576
rect 9627 3520 9660 3576
rect 9716 3520 9749 3576
rect 9805 3520 9814 3576
rect 9382 3496 9814 3520
rect 9382 3440 9391 3496
rect 9447 3440 9481 3496
rect 9537 3440 9571 3496
rect 9627 3440 9660 3496
rect 9716 3440 9749 3496
rect 9805 3440 9814 3496
tri 8432 3399 8473 3440 se
rect 8473 3399 8680 3440
tri 3829 3263 3841 3275 se
rect 3841 3263 3892 3275
tri 3892 3263 3904 3275 nw
rect 7863 3390 8680 3399
tri 3789 3223 3829 3263 se
rect 3789 2900 3829 3223
tri 3829 3200 3892 3263 nw
rect 7999 3287 8680 3390
rect 9382 3416 9814 3440
rect 9382 3360 9391 3416
rect 9447 3360 9481 3416
rect 9537 3360 9571 3416
rect 9627 3360 9660 3416
rect 9716 3360 9749 3416
rect 9805 3360 9814 3416
rect 14029 3520 14038 3576
rect 14094 3520 14128 3576
rect 14184 3520 14218 3576
rect 14274 3520 14307 3576
rect 14363 3520 14396 3576
rect 14452 3520 14666 3576
rect 14029 3496 14666 3520
rect 14029 3440 14038 3496
rect 14094 3440 14128 3496
rect 14184 3440 14218 3496
rect 14274 3440 14307 3496
rect 14363 3440 14396 3496
rect 14452 3440 14666 3496
rect 14029 3416 14666 3440
rect 14029 3360 14038 3416
rect 14094 3360 14128 3416
rect 14184 3360 14218 3416
rect 14274 3360 14307 3416
rect 14363 3360 14396 3416
rect 14452 3360 14666 3416
rect 15558 3520 15567 3576
rect 15623 3520 15655 3576
rect 15711 3520 15743 3576
rect 15799 3520 15831 3576
rect 15887 3520 15918 3576
rect 15974 3520 15983 3576
rect 15558 3496 15983 3520
rect 15558 3440 15567 3496
rect 15623 3440 15655 3496
rect 15711 3440 15743 3496
rect 15799 3440 15831 3496
rect 15887 3440 15918 3496
rect 15974 3440 15983 3496
rect 16967 3460 17134 3676
rect 17270 3460 17272 3676
tri 20176 3680 20178 3682 se
rect 20178 3680 20494 3682
tri 20494 3680 20496 3682 sw
rect 20176 3628 20496 3680
tri 20176 3626 20178 3628 ne
rect 20178 3626 20494 3628
tri 20494 3626 20496 3628 nw
tri 24252 3626 24275 3649 se
rect 24275 3626 24330 3830
tri 24228 3602 24252 3626 se
rect 24252 3602 24330 3626
rect 24082 3550 24088 3602
rect 24140 3550 24152 3602
rect 24204 3550 24330 3602
rect 16967 3451 17272 3460
rect 15558 3416 15983 3440
rect 15558 3360 15567 3416
rect 15623 3360 15655 3416
rect 15711 3360 15743 3416
rect 15799 3360 15831 3416
rect 15887 3360 15918 3416
rect 15974 3360 15983 3416
tri 20176 3362 20178 3364 se
rect 20178 3362 20494 3364
tri 20494 3362 20496 3364 sw
tri 10437 3308 10459 3330 se
tri 10432 3303 10437 3308 se
rect 10437 3306 10459 3308
rect 10437 3303 10589 3306
rect 7999 3174 8558 3287
rect 7863 3165 8558 3174
tri 8558 3165 8680 3287 nw
tri 9986 3267 10022 3303 se
rect 10022 3278 10589 3303
rect 14029 3284 14666 3360
rect 20176 3310 20496 3362
tri 20176 3308 20178 3310 ne
rect 20178 3308 20494 3310
tri 20494 3308 20496 3310 nw
rect 10022 3267 10578 3278
tri 10578 3267 10589 3278 nw
rect 9986 3263 10574 3267
tri 10574 3263 10578 3267 nw
rect 9986 3237 10548 3263
tri 10548 3237 10574 3263 nw
tri 3789 2893 3796 2900 ne
rect 3796 2893 3829 2900
tri 3829 2893 3850 2914 sw
tri 3796 2860 3829 2893 ne
rect 3829 2860 3850 2893
tri 3829 2839 3850 2860 ne
tri 3850 2839 3904 2893 sw
tri 3850 2785 3904 2839 ne
tri 3904 2785 3958 2839 sw
tri 3904 2771 3918 2785 ne
tri 3759 2674 3835 2750 sw
rect 3707 2670 3835 2674
rect 3707 2618 3713 2670
rect 3765 2618 3777 2670
rect 3829 2618 3835 2670
rect 3918 1639 3958 2785
rect 4730 2446 4824 2448
rect 4880 2446 4943 2448
rect 4999 2446 5061 2448
rect 4730 2394 4736 2446
rect 4788 2394 4802 2446
rect 4920 2394 4934 2446
rect 5051 2394 5061 2446
rect 4730 2392 4824 2394
rect 4880 2392 4943 2394
rect 4999 2392 5061 2394
rect 5117 2392 5126 2448
rect 4730 2382 5126 2392
rect 4730 2330 4736 2382
rect 4788 2330 4802 2382
rect 4854 2368 4868 2382
rect 4920 2330 4934 2382
rect 4986 2368 4999 2382
rect 5051 2368 5064 2382
rect 5116 2368 5126 2382
rect 5051 2330 5061 2368
rect 4730 2318 4824 2330
rect 4880 2318 4943 2330
rect 4999 2318 5061 2330
rect 4730 2266 4736 2318
rect 4788 2266 4802 2318
rect 4854 2266 4868 2312
rect 4920 2266 4934 2318
rect 4986 2266 4999 2312
rect 5051 2312 5061 2318
rect 5117 2312 5126 2368
rect 5051 2266 5064 2312
rect 5116 2266 5122 2312
tri 3958 1639 3979 1660 sw
rect 9986 1651 10036 3237
tri 10036 3208 10065 3237 nw
tri 14824 3168 14851 3195 se
rect 14851 3168 14981 3280
tri 14399 3144 14423 3168 se
rect 14423 3160 14981 3168
rect 14423 3144 14965 3160
tri 14965 3144 14981 3160 nw
rect 14399 3102 14923 3144
tri 14923 3102 14965 3144 nw
rect 10184 2446 10583 2451
rect 10184 2394 10192 2446
rect 10244 2424 10258 2446
rect 10310 2424 10324 2446
rect 10251 2394 10258 2424
rect 10376 2394 10390 2446
rect 10442 2424 10455 2446
rect 10507 2424 10520 2446
rect 10507 2394 10513 2424
rect 10572 2394 10583 2446
rect 10184 2382 10195 2394
rect 10251 2382 10301 2394
rect 10357 2382 10407 2394
rect 10463 2382 10513 2394
rect 10569 2382 10583 2394
rect 10184 2330 10192 2382
rect 10251 2368 10258 2382
rect 10244 2344 10258 2368
rect 10310 2344 10324 2368
rect 10251 2330 10258 2344
rect 10376 2330 10390 2382
rect 10507 2368 10513 2382
rect 10442 2344 10455 2368
rect 10507 2344 10520 2368
rect 10507 2330 10513 2344
rect 10572 2330 10583 2382
rect 10184 2318 10195 2330
rect 10251 2318 10301 2330
rect 10357 2318 10407 2330
rect 10463 2318 10513 2330
rect 10569 2318 10583 2330
rect 10184 2266 10192 2318
rect 10251 2288 10258 2318
rect 10244 2266 10258 2288
rect 10310 2266 10324 2288
rect 10376 2266 10390 2318
rect 10507 2288 10513 2318
rect 10442 2266 10455 2288
rect 10507 2266 10520 2288
rect 10572 2266 10583 2318
rect 10184 2261 10583 2266
rect 11116 2446 11515 2451
rect 11116 2394 11124 2446
rect 11176 2424 11190 2446
rect 11242 2424 11256 2446
rect 11183 2394 11190 2424
rect 11308 2394 11322 2446
rect 11374 2424 11387 2446
rect 11439 2424 11452 2446
rect 11439 2394 11445 2424
rect 11504 2394 11515 2446
rect 11116 2382 11127 2394
rect 11183 2382 11233 2394
rect 11289 2382 11339 2394
rect 11395 2382 11445 2394
rect 11501 2382 11515 2394
rect 11116 2330 11124 2382
rect 11183 2368 11190 2382
rect 11176 2344 11190 2368
rect 11242 2344 11256 2368
rect 11183 2330 11190 2344
rect 11308 2330 11322 2382
rect 11439 2368 11445 2382
rect 11374 2344 11387 2368
rect 11439 2344 11452 2368
rect 11439 2330 11445 2344
rect 11504 2330 11515 2382
rect 11116 2318 11127 2330
rect 11183 2318 11233 2330
rect 11289 2318 11339 2330
rect 11395 2318 11445 2330
rect 11501 2318 11515 2330
rect 11116 2266 11124 2318
rect 11183 2288 11190 2318
rect 11176 2266 11190 2288
rect 11242 2266 11256 2288
rect 11308 2266 11322 2318
rect 11439 2288 11445 2318
rect 11374 2266 11387 2288
rect 11439 2266 11452 2288
rect 11504 2266 11515 2318
rect 11116 2261 11515 2266
tri 10036 1651 10040 1655 sw
tri 9974 1639 9986 1651 se
rect 9986 1639 10040 1651
rect 3918 1630 3983 1639
tri 3677 1562 3699 1584 sw
rect 3918 1574 3927 1630
rect 3625 1539 3699 1562
tri 3699 1539 3722 1562 sw
rect 3918 1550 3983 1574
tri 9949 1614 9974 1639 se
rect 9974 1614 10040 1639
tri 10040 1614 10077 1651 sw
rect 9949 1562 9955 1614
rect 10007 1562 10019 1614
rect 10071 1562 10077 1614
tri 14396 1562 14399 1565 se
rect 14399 1562 14449 3102
tri 14449 3085 14466 3102 nw
rect 24897 2582 25775 4351
rect 25875 4343 26095 4367
rect 25931 4287 25957 4343
rect 26013 4287 26039 4343
rect 25875 4263 26095 4287
rect 25931 4207 25957 4263
rect 26013 4207 26039 4263
rect 25875 4198 26095 4207
rect 16669 2446 17068 2451
rect 16669 2394 16677 2446
rect 16729 2424 16743 2446
rect 16795 2424 16809 2446
rect 16861 2424 16875 2446
rect 16927 2424 16940 2446
rect 16992 2424 17005 2446
rect 17057 2424 17068 2446
rect 16736 2394 16743 2424
rect 16669 2382 16680 2394
rect 16736 2382 16761 2394
rect 16817 2382 16842 2394
rect 16669 2330 16677 2382
rect 16736 2368 16743 2382
rect 16729 2344 16743 2368
rect 16795 2344 16809 2368
rect 16736 2330 16743 2344
rect 16669 2318 16680 2330
rect 16736 2318 16761 2330
rect 16817 2318 16842 2330
rect 16669 2266 16677 2318
rect 16736 2288 16743 2318
rect 17058 2288 17068 2424
rect 16729 2266 16743 2288
rect 16795 2266 16809 2288
rect 16861 2266 16875 2288
rect 16927 2266 16940 2288
rect 16992 2266 17005 2288
rect 17057 2266 17068 2288
rect 16669 2261 17068 2266
rect 17600 2446 17999 2451
rect 17600 2394 17608 2446
rect 17660 2424 17674 2446
rect 17726 2424 17740 2446
rect 17792 2424 17806 2446
rect 17858 2424 17871 2446
rect 17923 2424 17936 2446
rect 17988 2424 17999 2446
rect 17667 2394 17674 2424
rect 17600 2382 17611 2394
rect 17667 2382 17692 2394
rect 17748 2382 17773 2394
rect 17600 2330 17608 2382
rect 17667 2368 17674 2382
rect 17660 2344 17674 2368
rect 17726 2344 17740 2368
rect 17667 2330 17674 2344
rect 17600 2318 17611 2330
rect 17667 2318 17692 2330
rect 17748 2318 17773 2330
rect 17600 2266 17608 2318
rect 17667 2288 17674 2318
rect 17989 2288 17999 2424
rect 17660 2266 17674 2288
rect 17726 2266 17740 2288
rect 17792 2266 17806 2288
rect 17858 2266 17871 2288
rect 17923 2266 17936 2288
rect 17988 2266 17999 2288
rect 17600 2261 17999 2266
rect 23153 2446 23552 2451
rect 23153 2394 23161 2446
rect 23213 2394 23227 2446
rect 23279 2424 23293 2446
rect 23345 2424 23359 2446
rect 23411 2424 23424 2446
rect 23476 2424 23489 2446
rect 23541 2424 23552 2446
rect 23476 2394 23486 2424
rect 23153 2382 23243 2394
rect 23299 2382 23324 2394
rect 23380 2382 23405 2394
rect 23461 2382 23486 2394
rect 23153 2330 23161 2382
rect 23213 2330 23227 2382
rect 23476 2368 23486 2382
rect 23542 2368 23552 2424
rect 23279 2344 23293 2368
rect 23345 2344 23359 2368
rect 23411 2344 23424 2368
rect 23476 2344 23489 2368
rect 23541 2344 23552 2368
rect 23476 2330 23486 2344
rect 23153 2318 23243 2330
rect 23299 2318 23324 2330
rect 23380 2318 23405 2330
rect 23461 2318 23486 2330
rect 23153 2266 23161 2318
rect 23213 2266 23227 2318
rect 23476 2288 23486 2318
rect 23542 2288 23552 2344
rect 23279 2266 23293 2288
rect 23345 2266 23359 2288
rect 23411 2266 23424 2288
rect 23476 2266 23489 2288
rect 23541 2266 23552 2288
rect 23153 2261 23552 2266
rect 25871 2111 25880 2116
rect 25936 2111 26037 2116
rect 26093 2111 26102 2116
rect 25871 2059 25877 2111
rect 25936 2060 25961 2111
rect 25929 2059 25961 2060
rect 26013 2060 26037 2111
rect 26013 2059 26044 2060
rect 26096 2059 26102 2111
rect 25871 2036 26102 2059
rect 25871 2035 25880 2036
rect 25936 2035 26037 2036
rect 26093 2035 26102 2036
rect 25871 1983 25877 2035
rect 25936 1983 25961 2035
rect 26013 1983 26037 2035
rect 26096 1983 26102 2035
rect 25871 1980 25880 1983
rect 25936 1980 26037 1983
rect 26093 1980 26102 1983
rect 3625 1487 3647 1539
rect 3699 1487 3711 1539
rect 3763 1487 3769 1539
rect 3918 1494 3927 1550
tri 14373 1539 14396 1562 se
rect 14396 1539 14449 1562
tri 14449 1539 14473 1563 sw
rect 3918 1485 3983 1494
rect 14346 1487 14352 1539
rect 14404 1487 14416 1539
rect 14468 1487 14474 1539
rect 387 1399 9390 1455
rect 9446 1399 9480 1455
rect 9536 1399 9570 1455
rect 9626 1399 9659 1455
rect 9715 1399 9748 1455
rect 9804 1399 15563 1455
rect 15619 1399 15653 1455
rect 15709 1399 15743 1455
rect 15799 1399 15832 1455
rect 15888 1399 15921 1455
rect 15977 1399 15986 1455
rect 387 1375 15986 1399
rect 387 1319 9390 1375
rect 9446 1319 9480 1375
rect 9536 1319 9570 1375
rect 9626 1319 9659 1375
rect 9715 1319 9748 1375
rect 9804 1319 15563 1375
rect 15619 1319 15653 1375
rect 15709 1319 15743 1375
rect 15799 1319 15832 1375
rect 15888 1319 15921 1375
rect 15977 1319 15986 1375
rect 17129 1349 18356 1358
tri 320 -1285 387 -1218 se
rect 387 -1285 507 1319
tri 507 1284 542 1319 nw
rect 17185 1293 17219 1349
rect 17275 1302 18356 1349
rect 18412 1302 18439 1358
rect 18495 1302 18522 1358
rect 18578 1302 18587 1358
rect 17275 1293 18587 1302
rect 320 -1287 507 -1285
rect 320 -1339 326 -1287
rect 378 -1339 411 -1287
rect 463 -1339 507 -1287
rect 320 -1367 507 -1339
rect 320 -1419 326 -1367
rect 378 -1419 411 -1367
rect 463 -1419 507 -1367
rect 550 1252 14461 1284
rect 550 1196 14038 1252
rect 14094 1196 14128 1252
rect 14184 1196 14218 1252
rect 14274 1196 14307 1252
rect 14363 1196 14396 1252
rect 14452 1196 14461 1252
rect 550 1165 14461 1196
rect 17129 1224 18587 1293
rect 17185 1168 17219 1224
rect 17275 1216 18587 1224
rect 17275 1168 18356 1216
rect 550 1159 717 1165
tri 717 1159 723 1165 nw
rect 17129 1160 18356 1168
rect 18412 1160 18439 1216
rect 18495 1160 18522 1216
rect 18578 1160 18587 1216
rect 17129 1159 18587 1160
rect 550 -1296 671 1159
tri 671 1113 717 1159 nw
tri 671 -1296 759 -1208 sw
rect 550 -1323 1057 -1296
rect 550 -1360 671 -1323
tri 550 -1375 565 -1360 ne
rect 565 -1375 671 -1360
rect 723 -1375 753 -1323
rect 805 -1375 835 -1323
rect 887 -1375 917 -1323
rect 969 -1375 999 -1323
rect 1051 -1375 1057 -1323
tri 565 -1391 581 -1375 ne
rect 581 -1391 1057 -1375
tri 581 -1393 583 -1391 ne
rect 583 -1393 1057 -1391
rect 320 -1447 507 -1419
rect 320 -1499 326 -1447
rect 378 -1499 411 -1447
rect 463 -1466 507 -1447
rect 463 -1499 469 -1466
rect 320 -1527 469 -1499
tri 469 -1504 507 -1466 nw
rect 320 -1579 326 -1527
rect 378 -1579 411 -1527
rect 463 -1579 469 -1527
<< via2 >>
rect 3936 7396 3992 7398
rect 4016 7396 4072 7398
rect 3936 7344 3985 7396
rect 3985 7344 3992 7396
rect 4016 7344 4049 7396
rect 4049 7344 4072 7396
rect 3936 7342 3992 7344
rect 4016 7342 4072 7344
rect 25875 4687 25931 4743
rect 25957 4687 26013 4743
rect 26039 4687 26095 4743
rect 25875 4607 25931 4663
rect 25957 4607 26013 4663
rect 26039 4607 26095 4663
rect 25875 4527 25931 4583
rect 25957 4527 26013 4583
rect 26039 4527 26095 4583
rect 25875 4447 25931 4503
rect 25957 4447 26013 4503
rect 26039 4447 26095 4503
rect 25875 4367 25931 4423
rect 25957 4367 26013 4423
rect 26039 4367 26095 4423
rect 9391 3520 9447 3576
rect 9481 3520 9537 3576
rect 9571 3520 9627 3576
rect 9660 3520 9716 3576
rect 9749 3520 9805 3576
rect 9391 3440 9447 3496
rect 9481 3440 9537 3496
rect 9571 3440 9627 3496
rect 9660 3440 9716 3496
rect 9749 3440 9805 3496
rect 7863 3174 7999 3390
rect 9391 3360 9447 3416
rect 9481 3360 9537 3416
rect 9571 3360 9627 3416
rect 9660 3360 9716 3416
rect 9749 3360 9805 3416
rect 14038 3520 14094 3576
rect 14128 3520 14184 3576
rect 14218 3520 14274 3576
rect 14307 3520 14363 3576
rect 14396 3520 14452 3576
rect 14038 3440 14094 3496
rect 14128 3440 14184 3496
rect 14218 3440 14274 3496
rect 14307 3440 14363 3496
rect 14396 3440 14452 3496
rect 14038 3360 14094 3416
rect 14128 3360 14184 3416
rect 14218 3360 14274 3416
rect 14307 3360 14363 3416
rect 14396 3360 14452 3416
rect 15567 3520 15623 3576
rect 15655 3520 15711 3576
rect 15743 3520 15799 3576
rect 15831 3520 15887 3576
rect 15918 3520 15974 3576
rect 15567 3440 15623 3496
rect 15655 3440 15711 3496
rect 15743 3440 15799 3496
rect 15831 3440 15887 3496
rect 15918 3440 15974 3496
rect 17134 3460 17270 3676
rect 15567 3360 15623 3416
rect 15655 3360 15711 3416
rect 15743 3360 15799 3416
rect 15831 3360 15887 3416
rect 15918 3360 15974 3416
rect 4824 2446 4880 2448
rect 4943 2446 4999 2448
rect 5061 2446 5117 2448
rect 4824 2394 4854 2446
rect 4854 2394 4868 2446
rect 4868 2394 4880 2446
rect 4943 2394 4986 2446
rect 4986 2394 4999 2446
rect 5061 2394 5064 2446
rect 5064 2394 5116 2446
rect 5116 2394 5117 2446
rect 4824 2392 4880 2394
rect 4943 2392 4999 2394
rect 5061 2392 5117 2394
rect 4824 2330 4854 2368
rect 4854 2330 4868 2368
rect 4868 2330 4880 2368
rect 4943 2330 4986 2368
rect 4986 2330 4999 2368
rect 5061 2330 5064 2368
rect 5064 2330 5116 2368
rect 5116 2330 5117 2368
rect 4824 2318 4880 2330
rect 4943 2318 4999 2330
rect 5061 2318 5117 2330
rect 4824 2312 4854 2318
rect 4854 2312 4868 2318
rect 4868 2312 4880 2318
rect 4943 2312 4986 2318
rect 4986 2312 4999 2318
rect 5061 2312 5064 2318
rect 5064 2312 5116 2318
rect 5116 2312 5117 2318
rect 10195 2394 10244 2424
rect 10244 2394 10251 2424
rect 10301 2394 10310 2424
rect 10310 2394 10324 2424
rect 10324 2394 10357 2424
rect 10407 2394 10442 2424
rect 10442 2394 10455 2424
rect 10455 2394 10463 2424
rect 10513 2394 10520 2424
rect 10520 2394 10569 2424
rect 10195 2382 10251 2394
rect 10301 2382 10357 2394
rect 10407 2382 10463 2394
rect 10513 2382 10569 2394
rect 10195 2368 10244 2382
rect 10244 2368 10251 2382
rect 10301 2368 10310 2382
rect 10310 2368 10324 2382
rect 10324 2368 10357 2382
rect 10195 2330 10244 2344
rect 10244 2330 10251 2344
rect 10301 2330 10310 2344
rect 10310 2330 10324 2344
rect 10324 2330 10357 2344
rect 10407 2368 10442 2382
rect 10442 2368 10455 2382
rect 10455 2368 10463 2382
rect 10513 2368 10520 2382
rect 10520 2368 10569 2382
rect 10407 2330 10442 2344
rect 10442 2330 10455 2344
rect 10455 2330 10463 2344
rect 10513 2330 10520 2344
rect 10520 2330 10569 2344
rect 10195 2318 10251 2330
rect 10301 2318 10357 2330
rect 10407 2318 10463 2330
rect 10513 2318 10569 2330
rect 10195 2288 10244 2318
rect 10244 2288 10251 2318
rect 10301 2288 10310 2318
rect 10310 2288 10324 2318
rect 10324 2288 10357 2318
rect 10407 2288 10442 2318
rect 10442 2288 10455 2318
rect 10455 2288 10463 2318
rect 10513 2288 10520 2318
rect 10520 2288 10569 2318
rect 11127 2394 11176 2424
rect 11176 2394 11183 2424
rect 11233 2394 11242 2424
rect 11242 2394 11256 2424
rect 11256 2394 11289 2424
rect 11339 2394 11374 2424
rect 11374 2394 11387 2424
rect 11387 2394 11395 2424
rect 11445 2394 11452 2424
rect 11452 2394 11501 2424
rect 11127 2382 11183 2394
rect 11233 2382 11289 2394
rect 11339 2382 11395 2394
rect 11445 2382 11501 2394
rect 11127 2368 11176 2382
rect 11176 2368 11183 2382
rect 11233 2368 11242 2382
rect 11242 2368 11256 2382
rect 11256 2368 11289 2382
rect 11127 2330 11176 2344
rect 11176 2330 11183 2344
rect 11233 2330 11242 2344
rect 11242 2330 11256 2344
rect 11256 2330 11289 2344
rect 11339 2368 11374 2382
rect 11374 2368 11387 2382
rect 11387 2368 11395 2382
rect 11445 2368 11452 2382
rect 11452 2368 11501 2382
rect 11339 2330 11374 2344
rect 11374 2330 11387 2344
rect 11387 2330 11395 2344
rect 11445 2330 11452 2344
rect 11452 2330 11501 2344
rect 11127 2318 11183 2330
rect 11233 2318 11289 2330
rect 11339 2318 11395 2330
rect 11445 2318 11501 2330
rect 11127 2288 11176 2318
rect 11176 2288 11183 2318
rect 11233 2288 11242 2318
rect 11242 2288 11256 2318
rect 11256 2288 11289 2318
rect 11339 2288 11374 2318
rect 11374 2288 11387 2318
rect 11387 2288 11395 2318
rect 11445 2288 11452 2318
rect 11452 2288 11501 2318
rect 3927 1574 3983 1630
rect 25875 4287 25931 4343
rect 25957 4287 26013 4343
rect 26039 4287 26095 4343
rect 25875 4207 25931 4263
rect 25957 4207 26013 4263
rect 26039 4207 26095 4263
rect 16680 2394 16729 2424
rect 16729 2394 16736 2424
rect 16761 2394 16795 2424
rect 16795 2394 16809 2424
rect 16809 2394 16817 2424
rect 16842 2394 16861 2424
rect 16861 2394 16875 2424
rect 16875 2394 16927 2424
rect 16927 2394 16940 2424
rect 16940 2394 16992 2424
rect 16992 2394 17005 2424
rect 17005 2394 17057 2424
rect 17057 2394 17058 2424
rect 16680 2382 16736 2394
rect 16761 2382 16817 2394
rect 16842 2382 17058 2394
rect 16680 2368 16729 2382
rect 16729 2368 16736 2382
rect 16761 2368 16795 2382
rect 16795 2368 16809 2382
rect 16809 2368 16817 2382
rect 16680 2330 16729 2344
rect 16729 2330 16736 2344
rect 16761 2330 16795 2344
rect 16795 2330 16809 2344
rect 16809 2330 16817 2344
rect 16842 2330 16861 2382
rect 16861 2330 16875 2382
rect 16875 2330 16927 2382
rect 16927 2330 16940 2382
rect 16940 2330 16992 2382
rect 16992 2330 17005 2382
rect 17005 2330 17057 2382
rect 17057 2330 17058 2382
rect 16680 2318 16736 2330
rect 16761 2318 16817 2330
rect 16842 2318 17058 2330
rect 16680 2288 16729 2318
rect 16729 2288 16736 2318
rect 16761 2288 16795 2318
rect 16795 2288 16809 2318
rect 16809 2288 16817 2318
rect 16842 2288 16861 2318
rect 16861 2288 16875 2318
rect 16875 2288 16927 2318
rect 16927 2288 16940 2318
rect 16940 2288 16992 2318
rect 16992 2288 17005 2318
rect 17005 2288 17057 2318
rect 17057 2288 17058 2318
rect 17611 2394 17660 2424
rect 17660 2394 17667 2424
rect 17692 2394 17726 2424
rect 17726 2394 17740 2424
rect 17740 2394 17748 2424
rect 17773 2394 17792 2424
rect 17792 2394 17806 2424
rect 17806 2394 17858 2424
rect 17858 2394 17871 2424
rect 17871 2394 17923 2424
rect 17923 2394 17936 2424
rect 17936 2394 17988 2424
rect 17988 2394 17989 2424
rect 17611 2382 17667 2394
rect 17692 2382 17748 2394
rect 17773 2382 17989 2394
rect 17611 2368 17660 2382
rect 17660 2368 17667 2382
rect 17692 2368 17726 2382
rect 17726 2368 17740 2382
rect 17740 2368 17748 2382
rect 17611 2330 17660 2344
rect 17660 2330 17667 2344
rect 17692 2330 17726 2344
rect 17726 2330 17740 2344
rect 17740 2330 17748 2344
rect 17773 2330 17792 2382
rect 17792 2330 17806 2382
rect 17806 2330 17858 2382
rect 17858 2330 17871 2382
rect 17871 2330 17923 2382
rect 17923 2330 17936 2382
rect 17936 2330 17988 2382
rect 17988 2330 17989 2382
rect 17611 2318 17667 2330
rect 17692 2318 17748 2330
rect 17773 2318 17989 2330
rect 17611 2288 17660 2318
rect 17660 2288 17667 2318
rect 17692 2288 17726 2318
rect 17726 2288 17740 2318
rect 17740 2288 17748 2318
rect 17773 2288 17792 2318
rect 17792 2288 17806 2318
rect 17806 2288 17858 2318
rect 17858 2288 17871 2318
rect 17871 2288 17923 2318
rect 17923 2288 17936 2318
rect 17936 2288 17988 2318
rect 17988 2288 17989 2318
rect 23243 2394 23279 2424
rect 23279 2394 23293 2424
rect 23293 2394 23299 2424
rect 23324 2394 23345 2424
rect 23345 2394 23359 2424
rect 23359 2394 23380 2424
rect 23405 2394 23411 2424
rect 23411 2394 23424 2424
rect 23424 2394 23461 2424
rect 23486 2394 23489 2424
rect 23489 2394 23541 2424
rect 23541 2394 23542 2424
rect 23243 2382 23299 2394
rect 23324 2382 23380 2394
rect 23405 2382 23461 2394
rect 23486 2382 23542 2394
rect 23243 2368 23279 2382
rect 23279 2368 23293 2382
rect 23293 2368 23299 2382
rect 23324 2368 23345 2382
rect 23345 2368 23359 2382
rect 23359 2368 23380 2382
rect 23405 2368 23411 2382
rect 23411 2368 23424 2382
rect 23424 2368 23461 2382
rect 23486 2368 23489 2382
rect 23489 2368 23541 2382
rect 23541 2368 23542 2382
rect 23243 2330 23279 2344
rect 23279 2330 23293 2344
rect 23293 2330 23299 2344
rect 23324 2330 23345 2344
rect 23345 2330 23359 2344
rect 23359 2330 23380 2344
rect 23405 2330 23411 2344
rect 23411 2330 23424 2344
rect 23424 2330 23461 2344
rect 23486 2330 23489 2344
rect 23489 2330 23541 2344
rect 23541 2330 23542 2344
rect 23243 2318 23299 2330
rect 23324 2318 23380 2330
rect 23405 2318 23461 2330
rect 23486 2318 23542 2330
rect 23243 2288 23279 2318
rect 23279 2288 23293 2318
rect 23293 2288 23299 2318
rect 23324 2288 23345 2318
rect 23345 2288 23359 2318
rect 23359 2288 23380 2318
rect 23405 2288 23411 2318
rect 23411 2288 23424 2318
rect 23424 2288 23461 2318
rect 23486 2288 23489 2318
rect 23489 2288 23541 2318
rect 23541 2288 23542 2318
rect 25880 2111 25936 2116
rect 26037 2111 26093 2116
rect 25880 2060 25929 2111
rect 25929 2060 25936 2111
rect 26037 2060 26044 2111
rect 26044 2060 26093 2111
rect 25880 2035 25936 2036
rect 26037 2035 26093 2036
rect 25880 1983 25929 2035
rect 25929 1983 25936 2035
rect 26037 1983 26044 2035
rect 26044 1983 26093 2035
rect 25880 1980 25936 1983
rect 26037 1980 26093 1983
rect 3927 1494 3983 1550
rect 9390 1399 9446 1455
rect 9480 1399 9536 1455
rect 9570 1399 9626 1455
rect 9659 1399 9715 1455
rect 9748 1399 9804 1455
rect 15563 1399 15619 1455
rect 15653 1399 15709 1455
rect 15743 1399 15799 1455
rect 15832 1399 15888 1455
rect 15921 1399 15977 1455
rect 9390 1319 9446 1375
rect 9480 1319 9536 1375
rect 9570 1319 9626 1375
rect 9659 1319 9715 1375
rect 9748 1319 9804 1375
rect 15563 1319 15619 1375
rect 15653 1319 15709 1375
rect 15743 1319 15799 1375
rect 15832 1319 15888 1375
rect 15921 1319 15977 1375
rect 17129 1293 17185 1349
rect 17219 1293 17275 1349
rect 18356 1302 18412 1358
rect 18439 1302 18495 1358
rect 18522 1302 18578 1358
rect 14038 1196 14094 1252
rect 14128 1196 14184 1252
rect 14218 1196 14274 1252
rect 14307 1196 14363 1252
rect 14396 1196 14452 1252
rect 17129 1168 17185 1224
rect 17219 1168 17275 1224
rect 18356 1160 18412 1216
rect 18439 1160 18495 1216
rect 18522 1160 18578 1216
<< metal3 >>
rect 2308 24975 2548 25028
rect 18174 9317 19056 9349
tri 19056 9317 19057 9318 sw
rect 3931 7398 4077 7403
rect 3931 7342 3936 7398
rect 3992 7342 4016 7398
rect 4072 7342 4077 7398
rect 3931 7337 4077 7342
rect 3931 1980 4017 7337
tri 4017 7277 4077 7337 nw
rect 5206 6842 6088 8947
rect 8877 8423 10010 8954
tri 8877 8172 9128 8423 ne
rect 9128 6842 10010 8423
rect 11690 8947 12572 8953
tri 12572 8947 12578 8953 sw
rect 11690 8423 13037 8947
rect 11690 6842 12572 8423
tri 12572 8105 12890 8423 nw
rect 15612 6842 16494 8954
rect 18174 8453 19057 9317
rect 18174 6842 19056 8453
tri 19056 8452 19057 8453 nw
rect 22096 6842 22978 9349
rect 25869 4743 26102 4753
rect 25869 4687 25875 4743
rect 25931 4687 25957 4743
rect 26013 4687 26039 4743
rect 26095 4687 26102 4743
rect 25869 4663 26102 4687
rect 25869 4607 25875 4663
rect 25931 4607 25957 4663
rect 26013 4607 26039 4663
rect 26095 4607 26102 4663
rect 25869 4583 26102 4607
rect 25869 4527 25875 4583
rect 25931 4527 25957 4583
rect 26013 4527 26039 4583
rect 26095 4527 26102 4583
rect 25869 4503 26102 4527
rect 25869 4447 25875 4503
rect 25931 4447 25957 4503
rect 26013 4447 26039 4503
rect 26095 4447 26102 4503
rect 25869 4423 26102 4447
rect 25869 4367 25875 4423
rect 25931 4367 25957 4423
rect 26013 4367 26039 4423
rect 26095 4367 26102 4423
rect 25869 4343 26102 4367
rect 25869 4287 25875 4343
rect 25931 4287 25957 4343
rect 26013 4287 26039 4343
rect 26095 4287 26102 4343
rect 25869 4263 26102 4287
rect 25869 4207 25875 4263
rect 25931 4207 25957 4263
rect 26013 4207 26039 4263
rect 26095 4207 26102 4263
rect 17129 3676 17275 3681
rect 9385 3576 9810 3581
rect 9385 3520 9391 3576
rect 9447 3520 9481 3576
rect 9537 3520 9571 3576
rect 9627 3520 9660 3576
rect 9716 3520 9749 3576
rect 9805 3520 9810 3576
rect 9385 3496 9810 3520
rect 9385 3440 9391 3496
rect 9447 3440 9481 3496
rect 9537 3440 9571 3496
rect 9627 3440 9660 3496
rect 9716 3440 9749 3496
rect 9805 3440 9810 3496
rect 9385 3416 9810 3440
rect 7858 3390 8004 3395
rect 7858 3174 7863 3390
rect 7999 3174 8004 3390
rect 4819 2448 5122 2453
rect 4819 2392 4824 2448
rect 4880 2392 4943 2448
rect 4999 2392 5061 2448
rect 5117 2392 5122 2448
rect 4819 2368 5122 2392
rect 4819 2312 4824 2368
rect 4880 2312 4943 2368
rect 4999 2312 5061 2368
rect 5117 2312 5122 2368
rect 4819 2307 5122 2312
tri 4017 1980 4044 2007 sw
rect 3931 1956 4044 1980
tri 3931 1910 3977 1956 ne
rect 3977 1910 4044 1956
tri 4044 1910 4114 1980 sw
tri 3977 1870 4017 1910 ne
rect 4017 1870 4114 1910
tri 4017 1773 4114 1870 ne
tri 4114 1773 4251 1910 sw
tri 4114 1722 4165 1773 ne
rect 3922 1630 3996 1635
rect 3922 1574 3927 1630
rect 3983 1574 3996 1630
rect 3922 1550 3996 1574
rect 3922 1494 3927 1550
rect 3983 1494 3996 1550
rect 3922 1457 3996 1494
tri 3922 1455 3924 1457 ne
rect 3924 1455 3996 1457
tri 3996 1455 4038 1497 sw
tri 3924 1399 3980 1455 ne
rect 3980 1399 4038 1455
tri 4038 1399 4094 1455 sw
tri 3980 1390 3989 1399 ne
rect 3989 1390 4094 1399
tri 4094 1390 4103 1399 sw
tri 3989 1383 3996 1390 ne
rect 3996 1383 4103 1390
tri 3996 1375 4004 1383 ne
rect 4004 1375 4103 1383
tri 4004 1362 4017 1375 ne
rect 4017 822 4103 1375
rect 4165 822 4251 1773
rect 7858 877 8004 3174
rect 9385 3360 9391 3416
rect 9447 3360 9481 3416
rect 9537 3360 9571 3416
rect 9627 3360 9660 3416
rect 9716 3360 9749 3416
rect 9805 3360 9810 3416
rect 9385 1455 9810 3360
rect 14033 3576 14457 3581
rect 14033 3520 14038 3576
rect 14094 3520 14128 3576
rect 14184 3520 14218 3576
rect 14274 3520 14307 3576
rect 14363 3520 14396 3576
rect 14452 3520 14457 3576
rect 14033 3496 14457 3520
rect 14033 3440 14038 3496
rect 14094 3440 14128 3496
rect 14184 3440 14218 3496
rect 14274 3440 14307 3496
rect 14363 3440 14396 3496
rect 14452 3440 14457 3496
rect 14033 3416 14457 3440
rect 14033 3360 14038 3416
rect 14094 3360 14128 3416
rect 14184 3360 14218 3416
rect 14274 3360 14307 3416
rect 14363 3360 14396 3416
rect 14452 3360 14457 3416
rect 10190 2424 10574 2429
rect 10190 2368 10195 2424
rect 10251 2368 10301 2424
rect 10357 2368 10407 2424
rect 10463 2368 10513 2424
rect 10569 2368 10574 2424
rect 10190 2344 10574 2368
rect 10190 2288 10195 2344
rect 10251 2288 10301 2344
rect 10357 2288 10407 2344
rect 10463 2288 10513 2344
rect 10569 2288 10574 2344
rect 10190 2283 10574 2288
rect 11122 2424 11506 2429
rect 11122 2368 11127 2424
rect 11183 2368 11233 2424
rect 11289 2368 11339 2424
rect 11395 2368 11445 2424
rect 11501 2368 11506 2424
rect 11122 2344 11506 2368
rect 11122 2288 11127 2344
rect 11183 2288 11233 2344
rect 11289 2288 11339 2344
rect 11395 2288 11445 2344
rect 11501 2288 11506 2344
rect 11122 2283 11506 2288
rect 9385 1399 9390 1455
rect 9446 1399 9480 1455
rect 9536 1399 9570 1455
rect 9626 1399 9659 1455
rect 9715 1399 9748 1455
rect 9804 1399 9810 1455
rect 9385 1375 9810 1399
rect 9385 1319 9390 1375
rect 9446 1319 9480 1375
rect 9536 1319 9570 1375
rect 9626 1319 9659 1375
rect 9715 1319 9748 1375
rect 9804 1319 9810 1375
rect 9385 1314 9810 1319
rect 14033 1252 14457 3360
rect 15558 3576 15983 3581
rect 15558 3520 15567 3576
rect 15623 3520 15655 3576
rect 15711 3520 15743 3576
rect 15799 3520 15831 3576
rect 15887 3520 15918 3576
rect 15974 3520 15983 3576
rect 15558 3496 15983 3520
rect 15558 3440 15567 3496
rect 15623 3440 15655 3496
rect 15711 3440 15743 3496
rect 15799 3440 15831 3496
rect 15887 3440 15918 3496
rect 15974 3440 15983 3496
rect 15558 3416 15983 3440
rect 15558 3360 15567 3416
rect 15623 3360 15655 3416
rect 15711 3360 15743 3416
rect 15799 3360 15831 3416
rect 15887 3360 15918 3416
rect 15974 3360 15983 3416
rect 15558 1455 15983 3360
rect 17129 3460 17134 3676
rect 17270 3460 17275 3676
rect 16675 2424 17063 2429
rect 16675 2368 16680 2424
rect 16736 2368 16761 2424
rect 16817 2368 16842 2424
rect 16675 2344 16842 2368
rect 16675 2288 16680 2344
rect 16736 2288 16761 2344
rect 16817 2288 16842 2344
rect 17058 2288 17063 2424
rect 16675 2283 17063 2288
rect 15558 1399 15563 1455
rect 15619 1399 15653 1455
rect 15709 1399 15743 1455
rect 15799 1399 15832 1455
rect 15888 1399 15921 1455
rect 15977 1399 15983 1455
rect 15558 1375 15983 1399
rect 15558 1319 15563 1375
rect 15619 1319 15653 1375
rect 15709 1319 15743 1375
rect 15799 1319 15832 1375
rect 15888 1319 15921 1375
rect 15977 1319 15983 1375
rect 15558 1314 15983 1319
tri 17124 1358 17129 1363 se
rect 17129 1358 17275 3460
rect 17606 2424 17994 2429
rect 17606 2368 17611 2424
rect 17667 2368 17692 2424
rect 17748 2368 17773 2424
rect 17606 2344 17773 2368
rect 17606 2288 17611 2344
rect 17667 2288 17692 2344
rect 17748 2288 17773 2344
rect 17989 2288 17994 2424
rect 17606 2283 17994 2288
rect 23238 2424 23547 2429
rect 23238 2368 23243 2424
rect 23299 2368 23324 2424
rect 23380 2368 23405 2424
rect 23461 2368 23486 2424
rect 23542 2368 23547 2424
rect 23238 2344 23547 2368
rect 23238 2288 23243 2344
rect 23299 2288 23324 2344
rect 23380 2288 23405 2344
rect 23461 2288 23486 2344
rect 23542 2288 23547 2344
rect 23238 2283 23547 2288
rect 25869 2116 26102 4207
rect 25869 2060 25880 2116
rect 25936 2060 26037 2116
rect 26093 2060 26102 2116
rect 25869 2036 26102 2060
rect 25869 1980 25880 2036
rect 25936 1980 26037 2036
rect 26093 1980 26102 2036
rect 25869 1975 26102 1980
tri 17275 1358 17280 1363 sw
rect 17124 1349 17280 1358
rect 14033 1196 14038 1252
rect 14094 1196 14128 1252
rect 14184 1196 14218 1252
rect 14274 1196 14307 1252
rect 14363 1196 14396 1252
rect 14452 1196 14457 1252
rect 14033 1160 14457 1196
rect 17124 1293 17129 1349
rect 17185 1293 17219 1349
rect 17275 1293 17280 1349
rect 17124 1224 17280 1293
rect 17124 1168 17129 1224
rect 17185 1168 17219 1224
rect 17275 1168 17280 1224
rect 17124 1159 17280 1168
rect 18347 1358 18587 1363
rect 18347 1302 18356 1358
rect 18412 1302 18439 1358
rect 18495 1302 18522 1358
rect 18578 1302 18587 1358
rect 18347 1216 18587 1302
rect 18347 1160 18356 1216
rect 18412 1160 18439 1216
rect 18495 1160 18522 1216
rect 18578 1160 18587 1216
tri 8004 877 8189 1062 sw
rect 7858 868 8189 877
tri 7858 822 7904 868 ne
rect 7904 822 8189 868
tri 7904 742 7984 822 ne
rect 7984 742 8189 822
rect 18347 717 18587 1160
use sky130_fd_io__gpio_ovtv2_pudrvr_strong  sky130_fd_io__gpio_ovtv2_pudrvr_strong_0
timestamp 1666464484
transform 1 0 4173 0 1 4091
box -2942 -3816 24038 16959
use sky130_fd_io__gpio_ovtv2_pudrvr_strong_slow  sky130_fd_io__gpio_ovtv2_pudrvr_strong_slow_0
timestamp 1666464484
transform -1 0 24145 0 -1 3742
box -4066 -17308 22914 3000
use sky130_fd_io__gpio_ovtv2_pudrvr_weak_1  sky130_fd_io__gpio_ovtv2_pudrvr_weak_1_0
timestamp 1666464484
transform 1 0 25741 0 1 4130
box -24510 -3388 2470 16920
use sky130_fd_io__gpio_ovtv2_vpbdrvr_tswitch  sky130_fd_io__gpio_ovtv2_vpbdrvr_tswitch_0
timestamp 1666464484
transform 1 0 -2712 0 1 7443
box 4295 -5902 26973 17585
<< labels >>
flabel comment s 4118 3395 4118 3395 0 FreeSans 1000 0 0 0 ------>
flabel comment s 4118 4014 4118 4014 0 FreeSans 1000 0 0 0 ------>
flabel comment s 4118 4614 4118 4614 0 FreeSans 1000 0 0 0 ------>
flabel comment s 3564 1657 3564 1657 0 FreeSans 400 90 0 0 PUG<0>
flabel comment s 3652 1657 3652 1657 0 FreeSans 400 90 0 0 PUG<1>
flabel comment s 26392 7935 26392 7935 0 FreeSans 400 0 0 0 TIE_HI
flabel comment s 26271 4109 26271 4109 0 FreeSans 400 0 0 0 TIE_HI_VPBDRVR
flabel comment s 4199 1178 4199 1178 0 FreeSans 800 90 0 0 PADLO
flabel comment s 3997 1178 3997 1178 0 FreeSans 800 90 0 0 PGHS_H_LATCH
<< properties >>
string GDS_END 38948156
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 37632632
<< end >>
