magic
tech sky130A
magscale 1 2
timestamp 1666199351
<< nwell >>
rect -38 261 2890 582
<< pwell >>
rect 1411 157 1769 201
rect 2190 157 2850 203
rect 1 21 2850 157
rect 29 -17 63 21
<< locali >>
rect 17 153 68 335
rect 210 153 267 335
rect 581 323 620 394
rect 581 211 713 323
rect 581 145 620 211
rect 2292 51 2371 493
rect 2682 299 2748 490
rect 2703 165 2748 299
rect 2682 55 2748 165
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2852 561
rect 17 415 69 493
rect 103 455 169 527
rect 203 451 421 493
rect 203 415 237 451
rect 455 417 507 493
rect 541 428 620 527
rect 17 369 237 415
rect 271 369 339 417
rect 108 255 164 335
rect 108 221 121 255
rect 155 221 164 255
rect 108 153 164 221
rect 301 144 339 369
rect 300 141 339 144
rect 396 352 507 417
rect 654 400 695 465
rect 729 455 795 527
rect 829 427 888 493
rect 396 181 447 352
rect 654 366 799 400
rect 481 255 547 318
rect 481 221 489 255
rect 523 221 547 255
rect 481 215 547 221
rect 396 143 506 181
rect 747 177 799 366
rect 299 129 339 141
rect 299 119 334 129
rect 17 17 140 119
rect 174 51 334 119
rect 368 17 418 109
rect 452 51 506 143
rect 654 143 799 177
rect 833 284 888 427
rect 933 323 978 493
rect 1012 427 1161 493
rect 1200 455 1266 527
rect 933 318 994 323
rect 943 289 994 318
rect 1041 315 1093 391
rect 833 218 898 284
rect 540 17 620 111
rect 654 51 694 143
rect 833 117 867 218
rect 943 184 977 289
rect 1127 279 1161 427
rect 1321 421 1364 490
rect 1412 425 1603 527
rect 1637 425 1798 492
rect 1832 447 1898 527
rect 1195 387 1364 421
rect 1764 413 1798 425
rect 1932 413 1986 490
rect 2020 447 2086 527
rect 1195 315 1229 387
rect 1328 289 1413 353
rect 1477 341 1611 391
rect 1028 255 1295 279
rect 1471 255 1541 265
rect 728 17 788 109
rect 822 51 867 117
rect 901 51 977 184
rect 1011 245 1541 255
rect 1011 51 1090 245
rect 1124 161 1203 203
rect 1261 195 1541 245
rect 1577 179 1611 341
rect 1684 215 1730 381
rect 1764 379 2086 413
rect 1776 323 1987 345
rect 1776 289 1788 323
rect 1822 305 1987 323
rect 2021 305 2086 379
rect 1822 289 1823 305
rect 1776 287 1823 289
rect 2120 271 2169 493
rect 2216 297 2258 527
rect 1766 179 1817 253
rect 1124 127 1310 161
rect 1133 17 1233 93
rect 1267 51 1310 127
rect 1344 17 1541 161
rect 1577 139 1817 179
rect 1857 237 2182 271
rect 1857 171 1903 237
rect 1937 169 2112 203
rect 1937 103 1971 169
rect 2146 117 2182 237
rect 1693 55 1971 103
rect 2007 17 2057 109
rect 2093 51 2182 117
rect 2224 17 2258 177
rect 2405 297 2463 527
rect 2506 265 2543 493
rect 2577 327 2648 527
rect 2506 199 2669 265
rect 2405 17 2463 177
rect 2506 51 2543 199
rect 2782 297 2835 527
rect 2577 17 2648 165
rect 2782 17 2835 177
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2852 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 2605 527 2639 561
rect 2697 527 2731 561
rect 2789 527 2823 561
rect 121 221 155 255
rect 489 221 523 255
rect 1788 289 1822 323
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
rect 2697 -17 2731 17
rect 2789 -17 2823 17
<< metal1 >>
rect 0 561 2852 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2852 561
rect 0 496 2852 527
rect 1316 320 1374 329
rect 1776 323 1834 329
rect 1776 320 1788 323
rect 1316 292 1788 320
rect 1316 283 1374 292
rect 1776 289 1788 292
rect 1822 289 1834 323
rect 1776 283 1834 289
rect 109 255 167 261
rect 109 221 121 255
rect 155 252 167 255
rect 477 255 535 261
rect 477 252 489 255
rect 155 224 489 252
rect 155 221 167 224
rect 109 215 167 221
rect 477 221 489 224
rect 523 221 535 255
rect 477 215 535 221
rect 0 17 2852 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2852 17
rect 0 -48 2852 -17
<< obsm1 >>
rect 753 388 811 397
rect 1040 388 1098 397
rect 1500 388 1558 397
rect 753 360 1558 388
rect 753 351 811 360
rect 1040 351 1098 360
rect 1500 351 1558 360
rect 293 320 351 329
rect 948 320 1006 329
rect 293 292 1006 320
rect 293 283 351 292
rect 948 283 1006 292
rect 845 252 903 261
rect 1684 252 1742 261
rect 845 224 1742 252
rect 845 215 903 224
rect 1684 215 1742 224
<< labels >>
rlabel locali s 581 145 620 211 6 CLK
port 1 nsew clock input
rlabel locali s 581 211 713 323 6 CLK
port 1 nsew clock input
rlabel locali s 581 323 620 394 6 CLK
port 1 nsew clock input
rlabel locali s 210 153 267 335 6 D
port 2 nsew signal input
rlabel locali s 17 153 68 335 6 SCD
port 3 nsew signal input
rlabel metal1 s 477 215 535 224 6 SCE
port 4 nsew signal input
rlabel metal1 s 109 215 167 224 6 SCE
port 4 nsew signal input
rlabel metal1 s 109 224 535 252 6 SCE
port 4 nsew signal input
rlabel metal1 s 477 252 535 261 6 SCE
port 4 nsew signal input
rlabel metal1 s 109 252 167 261 6 SCE
port 4 nsew signal input
rlabel metal1 s 1776 283 1834 292 6 SET_B
port 5 nsew signal input
rlabel metal1 s 1316 283 1374 292 6 SET_B
port 5 nsew signal input
rlabel metal1 s 1316 292 1834 320 6 SET_B
port 5 nsew signal input
rlabel metal1 s 1776 320 1834 329 6 SET_B
port 5 nsew signal input
rlabel metal1 s 1316 320 1374 329 6 SET_B
port 5 nsew signal input
rlabel metal1 s 0 -48 2852 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 1 21 2850 157 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 2190 157 2850 203 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 1411 157 1769 201 6 VNB
port 7 nsew ground bidirectional
rlabel nwell s -38 261 2890 582 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 496 2852 592 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 2682 55 2748 165 6 Q
port 10 nsew signal output
rlabel locali s 2703 165 2748 299 6 Q
port 10 nsew signal output
rlabel locali s 2682 299 2748 490 6 Q
port 10 nsew signal output
rlabel locali s 2292 51 2371 493 6 Q_N
port 11 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2852 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 264324
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 241692
<< end >>
