magic
tech sky130A
magscale 1 2
timestamp 1666464484
<< nwell >>
rect 2931 1501 5929 2209
rect 2931 1500 4697 1501
<< pwell >>
rect 2971 1203 5892 1395
<< mvnmos >>
rect 3050 1229 3170 1369
rect 3226 1229 3346 1369
rect 3402 1229 3522 1369
rect 3578 1229 3698 1369
rect 3754 1229 3874 1369
rect 3930 1229 4050 1369
rect 4106 1229 4226 1369
rect 4282 1229 4402 1369
rect 4458 1229 4578 1369
rect 4634 1229 4754 1369
rect 4810 1229 4930 1369
rect 4986 1229 5106 1369
rect 5162 1229 5282 1369
rect 5338 1229 5458 1369
rect 5514 1229 5634 1369
rect 5690 1229 5810 1369
<< mvpmos >>
rect 3050 1835 3170 2035
rect 3226 1835 3346 2035
rect 3402 1835 3522 2035
rect 3578 1835 3698 2035
rect 3754 1835 3874 2035
rect 3930 1835 4050 2035
rect 4106 1835 4226 2035
rect 4282 1835 4402 2035
rect 4458 1835 4578 2035
rect 4634 1835 4754 2035
rect 4810 1835 4930 2035
rect 4986 1835 5106 2035
rect 5162 1835 5282 2035
rect 5338 1835 5458 2035
rect 5514 1835 5634 2035
rect 5690 1835 5810 2035
rect 3050 1567 3170 1767
rect 3226 1567 3346 1767
rect 3402 1567 3522 1767
rect 3578 1567 3698 1767
rect 3754 1567 3874 1767
rect 3930 1567 4050 1767
rect 4106 1567 4226 1767
rect 4282 1567 4402 1767
rect 4458 1567 4578 1767
rect 4634 1567 4754 1767
rect 4810 1567 4930 1767
rect 4986 1567 5106 1767
rect 5162 1567 5282 1767
rect 5338 1567 5458 1767
rect 5514 1567 5634 1767
rect 5690 1567 5810 1767
<< mvndiff >>
rect 2997 1357 3050 1369
rect 2997 1323 3005 1357
rect 3039 1323 3050 1357
rect 2997 1289 3050 1323
rect 2997 1255 3005 1289
rect 3039 1255 3050 1289
rect 2997 1229 3050 1255
rect 3170 1357 3226 1369
rect 3170 1323 3181 1357
rect 3215 1323 3226 1357
rect 3170 1289 3226 1323
rect 3170 1255 3181 1289
rect 3215 1255 3226 1289
rect 3170 1229 3226 1255
rect 3346 1357 3402 1369
rect 3346 1323 3357 1357
rect 3391 1323 3402 1357
rect 3346 1289 3402 1323
rect 3346 1255 3357 1289
rect 3391 1255 3402 1289
rect 3346 1229 3402 1255
rect 3522 1357 3578 1369
rect 3522 1323 3533 1357
rect 3567 1323 3578 1357
rect 3522 1289 3578 1323
rect 3522 1255 3533 1289
rect 3567 1255 3578 1289
rect 3522 1229 3578 1255
rect 3698 1357 3754 1369
rect 3698 1323 3709 1357
rect 3743 1323 3754 1357
rect 3698 1289 3754 1323
rect 3698 1255 3709 1289
rect 3743 1255 3754 1289
rect 3698 1229 3754 1255
rect 3874 1357 3930 1369
rect 3874 1323 3885 1357
rect 3919 1323 3930 1357
rect 3874 1289 3930 1323
rect 3874 1255 3885 1289
rect 3919 1255 3930 1289
rect 3874 1229 3930 1255
rect 4050 1357 4106 1369
rect 4050 1323 4061 1357
rect 4095 1323 4106 1357
rect 4050 1289 4106 1323
rect 4050 1255 4061 1289
rect 4095 1255 4106 1289
rect 4050 1229 4106 1255
rect 4226 1357 4282 1369
rect 4226 1323 4237 1357
rect 4271 1323 4282 1357
rect 4226 1289 4282 1323
rect 4226 1255 4237 1289
rect 4271 1255 4282 1289
rect 4226 1229 4282 1255
rect 4402 1357 4458 1369
rect 4402 1323 4413 1357
rect 4447 1323 4458 1357
rect 4402 1289 4458 1323
rect 4402 1255 4413 1289
rect 4447 1255 4458 1289
rect 4402 1229 4458 1255
rect 4578 1357 4634 1369
rect 4578 1323 4589 1357
rect 4623 1323 4634 1357
rect 4578 1289 4634 1323
rect 4578 1255 4589 1289
rect 4623 1255 4634 1289
rect 4578 1229 4634 1255
rect 4754 1357 4810 1369
rect 4754 1323 4765 1357
rect 4799 1323 4810 1357
rect 4754 1289 4810 1323
rect 4754 1255 4765 1289
rect 4799 1255 4810 1289
rect 4754 1229 4810 1255
rect 4930 1357 4986 1369
rect 4930 1323 4941 1357
rect 4975 1323 4986 1357
rect 4930 1289 4986 1323
rect 4930 1255 4941 1289
rect 4975 1255 4986 1289
rect 4930 1229 4986 1255
rect 5106 1357 5162 1369
rect 5106 1323 5117 1357
rect 5151 1323 5162 1357
rect 5106 1289 5162 1323
rect 5106 1255 5117 1289
rect 5151 1255 5162 1289
rect 5106 1229 5162 1255
rect 5282 1357 5338 1369
rect 5282 1323 5293 1357
rect 5327 1323 5338 1357
rect 5282 1289 5338 1323
rect 5282 1255 5293 1289
rect 5327 1255 5338 1289
rect 5282 1229 5338 1255
rect 5458 1357 5514 1369
rect 5458 1323 5469 1357
rect 5503 1323 5514 1357
rect 5458 1289 5514 1323
rect 5458 1255 5469 1289
rect 5503 1255 5514 1289
rect 5458 1229 5514 1255
rect 5634 1357 5690 1369
rect 5634 1323 5645 1357
rect 5679 1323 5690 1357
rect 5634 1289 5690 1323
rect 5634 1255 5645 1289
rect 5679 1255 5690 1289
rect 5634 1229 5690 1255
rect 5810 1357 5866 1369
rect 5810 1323 5821 1357
rect 5855 1323 5866 1357
rect 5810 1289 5866 1323
rect 5810 1255 5821 1289
rect 5855 1255 5866 1289
rect 5810 1229 5866 1255
<< mvpdiff >>
rect 2997 2017 3050 2035
rect 2997 1983 3005 2017
rect 3039 1983 3050 2017
rect 2997 1949 3050 1983
rect 2997 1915 3005 1949
rect 3039 1915 3050 1949
rect 2997 1881 3050 1915
rect 2997 1847 3005 1881
rect 3039 1847 3050 1881
rect 2997 1835 3050 1847
rect 3170 2017 3226 2035
rect 3170 1983 3181 2017
rect 3215 1983 3226 2017
rect 3170 1949 3226 1983
rect 3170 1915 3181 1949
rect 3215 1915 3226 1949
rect 3170 1881 3226 1915
rect 3170 1847 3181 1881
rect 3215 1847 3226 1881
rect 3170 1835 3226 1847
rect 3346 2017 3402 2035
rect 3346 1983 3357 2017
rect 3391 1983 3402 2017
rect 3346 1949 3402 1983
rect 3346 1915 3357 1949
rect 3391 1915 3402 1949
rect 3346 1881 3402 1915
rect 3346 1847 3357 1881
rect 3391 1847 3402 1881
rect 3346 1835 3402 1847
rect 3522 2017 3578 2035
rect 3522 1983 3533 2017
rect 3567 1983 3578 2017
rect 3522 1949 3578 1983
rect 3522 1915 3533 1949
rect 3567 1915 3578 1949
rect 3522 1881 3578 1915
rect 3522 1847 3533 1881
rect 3567 1847 3578 1881
rect 3522 1835 3578 1847
rect 3698 2017 3754 2035
rect 3698 1983 3709 2017
rect 3743 1983 3754 2017
rect 3698 1949 3754 1983
rect 3698 1915 3709 1949
rect 3743 1915 3754 1949
rect 3698 1881 3754 1915
rect 3698 1847 3709 1881
rect 3743 1847 3754 1881
rect 3698 1835 3754 1847
rect 3874 2017 3930 2035
rect 3874 1983 3885 2017
rect 3919 1983 3930 2017
rect 3874 1949 3930 1983
rect 3874 1915 3885 1949
rect 3919 1915 3930 1949
rect 3874 1881 3930 1915
rect 3874 1847 3885 1881
rect 3919 1847 3930 1881
rect 3874 1835 3930 1847
rect 4050 2017 4106 2035
rect 4050 1983 4061 2017
rect 4095 1983 4106 2017
rect 4050 1949 4106 1983
rect 4050 1915 4061 1949
rect 4095 1915 4106 1949
rect 4050 1881 4106 1915
rect 4050 1847 4061 1881
rect 4095 1847 4106 1881
rect 4050 1835 4106 1847
rect 4226 2017 4282 2035
rect 4226 1983 4237 2017
rect 4271 1983 4282 2017
rect 4226 1949 4282 1983
rect 4226 1915 4237 1949
rect 4271 1915 4282 1949
rect 4226 1881 4282 1915
rect 4226 1847 4237 1881
rect 4271 1847 4282 1881
rect 4226 1835 4282 1847
rect 4402 2017 4458 2035
rect 4402 1983 4413 2017
rect 4447 1983 4458 2017
rect 4402 1949 4458 1983
rect 4402 1915 4413 1949
rect 4447 1915 4458 1949
rect 4402 1881 4458 1915
rect 4402 1847 4413 1881
rect 4447 1847 4458 1881
rect 4402 1835 4458 1847
rect 4578 2017 4634 2035
rect 4578 1983 4589 2017
rect 4623 1983 4634 2017
rect 4578 1949 4634 1983
rect 4578 1915 4589 1949
rect 4623 1915 4634 1949
rect 4578 1881 4634 1915
rect 4578 1847 4589 1881
rect 4623 1847 4634 1881
rect 4578 1835 4634 1847
rect 4754 2017 4810 2035
rect 4754 1983 4765 2017
rect 4799 1983 4810 2017
rect 4754 1949 4810 1983
rect 4754 1915 4765 1949
rect 4799 1915 4810 1949
rect 4754 1881 4810 1915
rect 4754 1847 4765 1881
rect 4799 1847 4810 1881
rect 4754 1835 4810 1847
rect 4930 2017 4986 2035
rect 4930 1983 4941 2017
rect 4975 1983 4986 2017
rect 4930 1949 4986 1983
rect 4930 1915 4941 1949
rect 4975 1915 4986 1949
rect 4930 1881 4986 1915
rect 4930 1847 4941 1881
rect 4975 1847 4986 1881
rect 4930 1835 4986 1847
rect 5106 2017 5162 2035
rect 5106 1983 5117 2017
rect 5151 1983 5162 2017
rect 5106 1949 5162 1983
rect 5106 1915 5117 1949
rect 5151 1915 5162 1949
rect 5106 1881 5162 1915
rect 5106 1847 5117 1881
rect 5151 1847 5162 1881
rect 5106 1835 5162 1847
rect 5282 2017 5338 2035
rect 5282 1983 5293 2017
rect 5327 1983 5338 2017
rect 5282 1949 5338 1983
rect 5282 1915 5293 1949
rect 5327 1915 5338 1949
rect 5282 1881 5338 1915
rect 5282 1847 5293 1881
rect 5327 1847 5338 1881
rect 5282 1835 5338 1847
rect 5458 2017 5514 2035
rect 5458 1983 5469 2017
rect 5503 1983 5514 2017
rect 5458 1949 5514 1983
rect 5458 1915 5469 1949
rect 5503 1915 5514 1949
rect 5458 1881 5514 1915
rect 5458 1847 5469 1881
rect 5503 1847 5514 1881
rect 5458 1835 5514 1847
rect 5634 2017 5690 2035
rect 5634 1983 5645 2017
rect 5679 1983 5690 2017
rect 5634 1949 5690 1983
rect 5634 1915 5645 1949
rect 5679 1915 5690 1949
rect 5634 1881 5690 1915
rect 5634 1847 5645 1881
rect 5679 1847 5690 1881
rect 5634 1835 5690 1847
rect 5810 2017 5863 2035
rect 5810 1983 5821 2017
rect 5855 1983 5863 2017
rect 5810 1949 5863 1983
rect 5810 1915 5821 1949
rect 5855 1915 5863 1949
rect 5810 1881 5863 1915
rect 5810 1847 5821 1881
rect 5855 1847 5863 1881
rect 5810 1835 5863 1847
rect 2997 1749 3050 1767
rect 2997 1715 3005 1749
rect 3039 1715 3050 1749
rect 2997 1681 3050 1715
rect 2997 1647 3005 1681
rect 3039 1647 3050 1681
rect 2997 1613 3050 1647
rect 2997 1579 3005 1613
rect 3039 1579 3050 1613
rect 2997 1567 3050 1579
rect 3170 1749 3226 1767
rect 3170 1715 3181 1749
rect 3215 1715 3226 1749
rect 3170 1681 3226 1715
rect 3170 1647 3181 1681
rect 3215 1647 3226 1681
rect 3170 1613 3226 1647
rect 3170 1579 3181 1613
rect 3215 1579 3226 1613
rect 3170 1567 3226 1579
rect 3346 1749 3402 1767
rect 3346 1715 3357 1749
rect 3391 1715 3402 1749
rect 3346 1681 3402 1715
rect 3346 1647 3357 1681
rect 3391 1647 3402 1681
rect 3346 1613 3402 1647
rect 3346 1579 3357 1613
rect 3391 1579 3402 1613
rect 3346 1567 3402 1579
rect 3522 1749 3578 1767
rect 3522 1715 3533 1749
rect 3567 1715 3578 1749
rect 3522 1681 3578 1715
rect 3522 1647 3533 1681
rect 3567 1647 3578 1681
rect 3522 1613 3578 1647
rect 3522 1579 3533 1613
rect 3567 1579 3578 1613
rect 3522 1567 3578 1579
rect 3698 1749 3754 1767
rect 3698 1715 3709 1749
rect 3743 1715 3754 1749
rect 3698 1681 3754 1715
rect 3698 1647 3709 1681
rect 3743 1647 3754 1681
rect 3698 1613 3754 1647
rect 3698 1579 3709 1613
rect 3743 1579 3754 1613
rect 3698 1567 3754 1579
rect 3874 1749 3930 1767
rect 3874 1715 3885 1749
rect 3919 1715 3930 1749
rect 3874 1681 3930 1715
rect 3874 1647 3885 1681
rect 3919 1647 3930 1681
rect 3874 1613 3930 1647
rect 3874 1579 3885 1613
rect 3919 1579 3930 1613
rect 3874 1567 3930 1579
rect 4050 1749 4106 1767
rect 4050 1715 4061 1749
rect 4095 1715 4106 1749
rect 4050 1681 4106 1715
rect 4050 1647 4061 1681
rect 4095 1647 4106 1681
rect 4050 1613 4106 1647
rect 4050 1579 4061 1613
rect 4095 1579 4106 1613
rect 4050 1567 4106 1579
rect 4226 1749 4282 1767
rect 4226 1715 4237 1749
rect 4271 1715 4282 1749
rect 4226 1681 4282 1715
rect 4226 1647 4237 1681
rect 4271 1647 4282 1681
rect 4226 1613 4282 1647
rect 4226 1579 4237 1613
rect 4271 1579 4282 1613
rect 4226 1567 4282 1579
rect 4402 1749 4458 1767
rect 4402 1715 4413 1749
rect 4447 1715 4458 1749
rect 4402 1681 4458 1715
rect 4402 1647 4413 1681
rect 4447 1647 4458 1681
rect 4402 1613 4458 1647
rect 4402 1579 4413 1613
rect 4447 1579 4458 1613
rect 4402 1567 4458 1579
rect 4578 1749 4634 1767
rect 4578 1715 4589 1749
rect 4623 1715 4634 1749
rect 4578 1681 4634 1715
rect 4578 1647 4589 1681
rect 4623 1647 4634 1681
rect 4578 1613 4634 1647
rect 4578 1579 4589 1613
rect 4623 1579 4634 1613
rect 4578 1567 4634 1579
rect 4754 1749 4810 1767
rect 4754 1715 4765 1749
rect 4799 1715 4810 1749
rect 4754 1681 4810 1715
rect 4754 1647 4765 1681
rect 4799 1647 4810 1681
rect 4754 1613 4810 1647
rect 4754 1579 4765 1613
rect 4799 1579 4810 1613
rect 4754 1567 4810 1579
rect 4930 1749 4986 1767
rect 4930 1715 4941 1749
rect 4975 1715 4986 1749
rect 4930 1681 4986 1715
rect 4930 1647 4941 1681
rect 4975 1647 4986 1681
rect 4930 1613 4986 1647
rect 4930 1579 4941 1613
rect 4975 1579 4986 1613
rect 4930 1567 4986 1579
rect 5106 1749 5162 1767
rect 5106 1715 5117 1749
rect 5151 1715 5162 1749
rect 5106 1681 5162 1715
rect 5106 1647 5117 1681
rect 5151 1647 5162 1681
rect 5106 1613 5162 1647
rect 5106 1579 5117 1613
rect 5151 1579 5162 1613
rect 5106 1567 5162 1579
rect 5282 1749 5338 1767
rect 5282 1715 5293 1749
rect 5327 1715 5338 1749
rect 5282 1681 5338 1715
rect 5282 1647 5293 1681
rect 5327 1647 5338 1681
rect 5282 1613 5338 1647
rect 5282 1579 5293 1613
rect 5327 1579 5338 1613
rect 5282 1567 5338 1579
rect 5458 1749 5514 1767
rect 5458 1715 5469 1749
rect 5503 1715 5514 1749
rect 5458 1681 5514 1715
rect 5458 1647 5469 1681
rect 5503 1647 5514 1681
rect 5458 1613 5514 1647
rect 5458 1579 5469 1613
rect 5503 1579 5514 1613
rect 5458 1567 5514 1579
rect 5634 1749 5690 1767
rect 5634 1715 5645 1749
rect 5679 1715 5690 1749
rect 5634 1681 5690 1715
rect 5634 1647 5645 1681
rect 5679 1647 5690 1681
rect 5634 1613 5690 1647
rect 5634 1579 5645 1613
rect 5679 1579 5690 1613
rect 5634 1567 5690 1579
rect 5810 1749 5863 1767
rect 5810 1715 5821 1749
rect 5855 1715 5863 1749
rect 5810 1681 5863 1715
rect 5810 1647 5821 1681
rect 5855 1647 5863 1681
rect 5810 1613 5863 1647
rect 5810 1579 5821 1613
rect 5855 1579 5863 1613
rect 5810 1567 5863 1579
<< mvndiffc >>
rect 3005 1323 3039 1357
rect 3005 1255 3039 1289
rect 3181 1323 3215 1357
rect 3181 1255 3215 1289
rect 3357 1323 3391 1357
rect 3357 1255 3391 1289
rect 3533 1323 3567 1357
rect 3533 1255 3567 1289
rect 3709 1323 3743 1357
rect 3709 1255 3743 1289
rect 3885 1323 3919 1357
rect 3885 1255 3919 1289
rect 4061 1323 4095 1357
rect 4061 1255 4095 1289
rect 4237 1323 4271 1357
rect 4237 1255 4271 1289
rect 4413 1323 4447 1357
rect 4413 1255 4447 1289
rect 4589 1323 4623 1357
rect 4589 1255 4623 1289
rect 4765 1323 4799 1357
rect 4765 1255 4799 1289
rect 4941 1323 4975 1357
rect 4941 1255 4975 1289
rect 5117 1323 5151 1357
rect 5117 1255 5151 1289
rect 5293 1323 5327 1357
rect 5293 1255 5327 1289
rect 5469 1323 5503 1357
rect 5469 1255 5503 1289
rect 5645 1323 5679 1357
rect 5645 1255 5679 1289
rect 5821 1323 5855 1357
rect 5821 1255 5855 1289
<< mvpdiffc >>
rect 3005 1983 3039 2017
rect 3005 1915 3039 1949
rect 3005 1847 3039 1881
rect 3181 1983 3215 2017
rect 3181 1915 3215 1949
rect 3181 1847 3215 1881
rect 3357 1983 3391 2017
rect 3357 1915 3391 1949
rect 3357 1847 3391 1881
rect 3533 1983 3567 2017
rect 3533 1915 3567 1949
rect 3533 1847 3567 1881
rect 3709 1983 3743 2017
rect 3709 1915 3743 1949
rect 3709 1847 3743 1881
rect 3885 1983 3919 2017
rect 3885 1915 3919 1949
rect 3885 1847 3919 1881
rect 4061 1983 4095 2017
rect 4061 1915 4095 1949
rect 4061 1847 4095 1881
rect 4237 1983 4271 2017
rect 4237 1915 4271 1949
rect 4237 1847 4271 1881
rect 4413 1983 4447 2017
rect 4413 1915 4447 1949
rect 4413 1847 4447 1881
rect 4589 1983 4623 2017
rect 4589 1915 4623 1949
rect 4589 1847 4623 1881
rect 4765 1983 4799 2017
rect 4765 1915 4799 1949
rect 4765 1847 4799 1881
rect 4941 1983 4975 2017
rect 4941 1915 4975 1949
rect 4941 1847 4975 1881
rect 5117 1983 5151 2017
rect 5117 1915 5151 1949
rect 5117 1847 5151 1881
rect 5293 1983 5327 2017
rect 5293 1915 5327 1949
rect 5293 1847 5327 1881
rect 5469 1983 5503 2017
rect 5469 1915 5503 1949
rect 5469 1847 5503 1881
rect 5645 1983 5679 2017
rect 5645 1915 5679 1949
rect 5645 1847 5679 1881
rect 5821 1983 5855 2017
rect 5821 1915 5855 1949
rect 5821 1847 5855 1881
rect 3005 1715 3039 1749
rect 3005 1647 3039 1681
rect 3005 1579 3039 1613
rect 3181 1715 3215 1749
rect 3181 1647 3215 1681
rect 3181 1579 3215 1613
rect 3357 1715 3391 1749
rect 3357 1647 3391 1681
rect 3357 1579 3391 1613
rect 3533 1715 3567 1749
rect 3533 1647 3567 1681
rect 3533 1579 3567 1613
rect 3709 1715 3743 1749
rect 3709 1647 3743 1681
rect 3709 1579 3743 1613
rect 3885 1715 3919 1749
rect 3885 1647 3919 1681
rect 3885 1579 3919 1613
rect 4061 1715 4095 1749
rect 4061 1647 4095 1681
rect 4061 1579 4095 1613
rect 4237 1715 4271 1749
rect 4237 1647 4271 1681
rect 4237 1579 4271 1613
rect 4413 1715 4447 1749
rect 4413 1647 4447 1681
rect 4413 1579 4447 1613
rect 4589 1715 4623 1749
rect 4589 1647 4623 1681
rect 4589 1579 4623 1613
rect 4765 1715 4799 1749
rect 4765 1647 4799 1681
rect 4765 1579 4799 1613
rect 4941 1715 4975 1749
rect 4941 1647 4975 1681
rect 4941 1579 4975 1613
rect 5117 1715 5151 1749
rect 5117 1647 5151 1681
rect 5117 1579 5151 1613
rect 5293 1715 5327 1749
rect 5293 1647 5327 1681
rect 5293 1579 5327 1613
rect 5469 1715 5503 1749
rect 5469 1647 5503 1681
rect 5469 1579 5503 1613
rect 5645 1715 5679 1749
rect 5645 1647 5679 1681
rect 5645 1579 5679 1613
rect 5821 1715 5855 1749
rect 5821 1647 5855 1681
rect 5821 1579 5855 1613
<< mvnsubdiff >>
rect 2997 2109 3021 2143
rect 3055 2109 3090 2143
rect 3124 2109 3159 2143
rect 3193 2109 3228 2143
rect 3262 2109 3297 2143
rect 3331 2109 3366 2143
rect 3400 2109 3435 2143
rect 3469 2109 3504 2143
rect 3538 2109 3573 2143
rect 3607 2109 3642 2143
rect 3676 2109 3711 2143
rect 3745 2109 3780 2143
rect 3814 2109 3849 2143
rect 3883 2109 3918 2143
rect 3952 2109 3987 2143
rect 4021 2109 4056 2143
rect 4090 2109 4125 2143
rect 4159 2109 4195 2143
rect 4229 2109 4265 2143
rect 4299 2109 4335 2143
rect 4369 2109 4405 2143
rect 4439 2109 4475 2143
rect 4509 2109 4545 2143
rect 4579 2109 4615 2143
rect 4649 2109 4685 2143
rect 4719 2109 4755 2143
rect 4789 2109 4825 2143
rect 4859 2109 4895 2143
rect 4929 2109 4965 2143
rect 4999 2109 5035 2143
rect 5069 2109 5105 2143
rect 5139 2109 5175 2143
rect 5209 2109 5245 2143
rect 5279 2109 5315 2143
rect 5349 2109 5385 2143
rect 5419 2109 5455 2143
rect 5489 2109 5525 2143
rect 5559 2109 5595 2143
rect 5629 2109 5665 2143
rect 5699 2109 5735 2143
rect 5769 2109 5805 2143
rect 5839 2109 5863 2143
<< mvnsubdiffcont >>
rect 3021 2109 3055 2143
rect 3090 2109 3124 2143
rect 3159 2109 3193 2143
rect 3228 2109 3262 2143
rect 3297 2109 3331 2143
rect 3366 2109 3400 2143
rect 3435 2109 3469 2143
rect 3504 2109 3538 2143
rect 3573 2109 3607 2143
rect 3642 2109 3676 2143
rect 3711 2109 3745 2143
rect 3780 2109 3814 2143
rect 3849 2109 3883 2143
rect 3918 2109 3952 2143
rect 3987 2109 4021 2143
rect 4056 2109 4090 2143
rect 4125 2109 4159 2143
rect 4195 2109 4229 2143
rect 4265 2109 4299 2143
rect 4335 2109 4369 2143
rect 4405 2109 4439 2143
rect 4475 2109 4509 2143
rect 4545 2109 4579 2143
rect 4615 2109 4649 2143
rect 4685 2109 4719 2143
rect 4755 2109 4789 2143
rect 4825 2109 4859 2143
rect 4895 2109 4929 2143
rect 4965 2109 4999 2143
rect 5035 2109 5069 2143
rect 5105 2109 5139 2143
rect 5175 2109 5209 2143
rect 5245 2109 5279 2143
rect 5315 2109 5349 2143
rect 5385 2109 5419 2143
rect 5455 2109 5489 2143
rect 5525 2109 5559 2143
rect 5595 2109 5629 2143
rect 5665 2109 5699 2143
rect 5735 2109 5769 2143
rect 5805 2109 5839 2143
<< poly >>
rect 3050 2035 3170 2061
rect 3226 2035 3346 2061
rect 3402 2035 3522 2061
rect 3578 2035 3698 2061
rect 3754 2035 3874 2061
rect 3930 2035 4050 2061
rect 4106 2035 4226 2061
rect 4282 2035 4402 2061
rect 4458 2035 4578 2061
rect 4634 2035 4754 2061
rect 4810 2035 4930 2061
rect 4986 2035 5106 2061
rect 5162 2035 5282 2061
rect 5338 2035 5458 2061
rect 5514 2035 5634 2061
rect 5690 2035 5810 2061
rect 3050 1767 3170 1835
rect 3226 1767 3346 1835
rect 3402 1767 3522 1835
rect 3578 1767 3698 1835
rect 3754 1767 3874 1835
rect 3930 1767 4050 1835
rect 4106 1767 4226 1835
rect 4282 1767 4402 1835
rect 4458 1767 4578 1835
rect 4634 1767 4754 1835
rect 4810 1767 4930 1835
rect 4986 1767 5106 1835
rect 5162 1767 5282 1835
rect 5338 1767 5458 1835
rect 5514 1767 5634 1835
rect 5690 1767 5810 1835
rect 3050 1541 3170 1567
rect 3226 1541 3346 1567
rect 3402 1541 3522 1567
rect 3578 1541 3698 1567
rect 3754 1541 3874 1567
rect 3930 1541 4050 1567
rect 4106 1541 4226 1567
rect 4282 1541 4402 1567
rect 3050 1486 4402 1541
rect 3050 1452 3084 1486
rect 3118 1452 3153 1486
rect 3187 1452 3222 1486
rect 3256 1452 3291 1486
rect 3325 1452 3360 1486
rect 3394 1452 3429 1486
rect 3463 1452 3498 1486
rect 3532 1452 3567 1486
rect 3601 1452 3636 1486
rect 3670 1452 3705 1486
rect 3739 1452 3774 1486
rect 3808 1452 3843 1486
rect 3877 1452 3912 1486
rect 3946 1452 3981 1486
rect 4015 1452 4050 1486
rect 4084 1452 4120 1486
rect 4154 1452 4190 1486
rect 4224 1452 4260 1486
rect 4294 1452 4330 1486
rect 4364 1452 4402 1486
rect 3050 1395 4402 1452
rect 3050 1369 3170 1395
rect 3226 1369 3346 1395
rect 3402 1369 3522 1395
rect 3578 1369 3698 1395
rect 3754 1369 3874 1395
rect 3930 1369 4050 1395
rect 4106 1369 4226 1395
rect 4282 1369 4402 1395
rect 4458 1541 4578 1567
rect 4634 1541 4754 1567
rect 4810 1541 4930 1567
rect 4986 1541 5106 1567
rect 5162 1541 5282 1567
rect 5338 1541 5458 1567
rect 5514 1541 5634 1567
rect 5690 1541 5810 1567
rect 4458 1486 5810 1541
rect 4458 1452 4582 1486
rect 4616 1452 4651 1486
rect 4685 1452 4720 1486
rect 4754 1452 4789 1486
rect 4823 1452 4858 1486
rect 4892 1452 4926 1486
rect 4960 1452 4994 1486
rect 5028 1452 5062 1486
rect 5096 1452 5130 1486
rect 5164 1452 5198 1486
rect 5232 1452 5266 1486
rect 5300 1452 5334 1486
rect 5368 1452 5402 1486
rect 5436 1452 5470 1486
rect 5504 1452 5538 1486
rect 5572 1452 5606 1486
rect 5640 1452 5674 1486
rect 5708 1452 5742 1486
rect 5776 1452 5810 1486
rect 4458 1395 5810 1452
rect 4458 1369 4578 1395
rect 4634 1369 4754 1395
rect 4810 1369 4930 1395
rect 4986 1369 5106 1395
rect 5162 1369 5282 1395
rect 5338 1369 5458 1395
rect 5514 1369 5634 1395
rect 5690 1369 5810 1395
rect 3050 1203 3170 1229
rect 3226 1203 3346 1229
rect 3402 1203 3522 1229
rect 3578 1203 3698 1229
rect 3754 1203 3874 1229
rect 3930 1203 4050 1229
rect 4106 1203 4226 1229
rect 4282 1203 4402 1229
rect 4458 1203 4578 1229
rect 4634 1203 4754 1229
rect 4810 1203 4930 1229
rect 4986 1203 5106 1229
rect 5162 1203 5282 1229
rect 5338 1203 5458 1229
rect 5514 1203 5634 1229
rect 5690 1203 5810 1229
<< polycont >>
rect 3084 1452 3118 1486
rect 3153 1452 3187 1486
rect 3222 1452 3256 1486
rect 3291 1452 3325 1486
rect 3360 1452 3394 1486
rect 3429 1452 3463 1486
rect 3498 1452 3532 1486
rect 3567 1452 3601 1486
rect 3636 1452 3670 1486
rect 3705 1452 3739 1486
rect 3774 1452 3808 1486
rect 3843 1452 3877 1486
rect 3912 1452 3946 1486
rect 3981 1452 4015 1486
rect 4050 1452 4084 1486
rect 4120 1452 4154 1486
rect 4190 1452 4224 1486
rect 4260 1452 4294 1486
rect 4330 1452 4364 1486
rect 4582 1452 4616 1486
rect 4651 1452 4685 1486
rect 4720 1452 4754 1486
rect 4789 1452 4823 1486
rect 4858 1452 4892 1486
rect 4926 1452 4960 1486
rect 4994 1452 5028 1486
rect 5062 1452 5096 1486
rect 5130 1452 5164 1486
rect 5198 1452 5232 1486
rect 5266 1452 5300 1486
rect 5334 1452 5368 1486
rect 5402 1452 5436 1486
rect 5470 1452 5504 1486
rect 5538 1452 5572 1486
rect 5606 1452 5640 1486
rect 5674 1452 5708 1486
rect 5742 1452 5776 1486
<< locali >>
rect 2997 2109 3021 2143
rect 3055 2109 3090 2143
rect 3124 2109 3155 2143
rect 3193 2109 3228 2143
rect 3262 2109 3297 2143
rect 3335 2109 3366 2143
rect 3408 2109 3435 2143
rect 3481 2109 3504 2143
rect 3554 2109 3573 2143
rect 3627 2109 3642 2143
rect 3700 2109 3711 2143
rect 3773 2109 3780 2143
rect 3846 2109 3849 2143
rect 3883 2109 3885 2143
rect 3952 2109 3958 2143
rect 4021 2109 4031 2143
rect 4090 2109 4104 2143
rect 4159 2109 4177 2143
rect 4229 2109 4250 2143
rect 4299 2109 4324 2143
rect 4369 2109 4398 2143
rect 4439 2109 4472 2143
rect 4509 2109 4545 2143
rect 4580 2109 4615 2143
rect 4654 2109 4685 2143
rect 4728 2109 4755 2143
rect 4802 2109 4825 2143
rect 4876 2109 4895 2143
rect 4950 2109 4965 2143
rect 5024 2109 5035 2143
rect 5098 2109 5105 2143
rect 5172 2109 5175 2143
rect 5209 2109 5212 2143
rect 5279 2109 5286 2143
rect 5349 2109 5360 2143
rect 5419 2109 5434 2143
rect 5489 2109 5508 2143
rect 5559 2109 5582 2143
rect 5629 2109 5656 2143
rect 5699 2109 5730 2143
rect 5769 2109 5804 2143
rect 5839 2109 5863 2143
rect 3005 2017 3039 2033
rect 3005 1949 3039 1983
rect 3005 1895 3039 1915
rect 3181 2017 3215 2029
rect 3181 1949 3215 1957
rect 3005 1881 3006 1895
rect 3040 1861 3078 1895
rect 3181 1881 3215 1915
rect 3357 2017 3391 2033
rect 3357 1949 3391 1983
rect 3357 1895 3391 1915
rect 3533 2017 3567 2029
rect 3533 1949 3567 1957
rect 3005 1749 3039 1847
rect 3005 1681 3039 1715
rect 3005 1613 3039 1647
rect 3005 1563 3039 1579
rect 3355 1881 3393 1895
rect 3355 1861 3357 1881
rect 3181 1749 3215 1847
rect 3181 1681 3215 1715
rect 3181 1613 3215 1647
rect 3181 1563 3215 1579
rect 3391 1861 3393 1881
rect 3533 1881 3567 1915
rect 3709 2017 3743 2033
rect 3709 1949 3743 1983
rect 3709 1895 3743 1915
rect 3885 2017 3919 2029
rect 3885 1949 3919 1957
rect 3357 1749 3391 1847
rect 3357 1681 3391 1715
rect 3357 1613 3391 1647
rect 3357 1563 3391 1579
rect 3707 1881 3745 1895
rect 3707 1861 3709 1881
rect 3533 1749 3567 1847
rect 3533 1681 3567 1715
rect 3533 1613 3567 1647
rect 3533 1563 3567 1579
rect 3743 1861 3745 1881
rect 3885 1881 3919 1915
rect 4061 2017 4095 2033
rect 4061 1949 4095 1983
rect 4061 1895 4095 1915
rect 4237 2017 4271 2029
rect 4237 1949 4271 1957
rect 3709 1749 3743 1847
rect 3709 1681 3743 1715
rect 3709 1613 3743 1647
rect 3709 1563 3743 1579
rect 4059 1881 4097 1895
rect 4059 1861 4061 1881
rect 3885 1749 3919 1847
rect 3885 1681 3919 1715
rect 3885 1613 3919 1647
rect 3885 1563 3919 1579
rect 4095 1861 4097 1881
rect 4237 1881 4271 1915
rect 4413 2017 4447 2033
rect 4413 1949 4447 1983
rect 4413 1895 4447 1915
rect 4589 2017 4623 2063
rect 4589 1949 4623 1983
rect 4061 1749 4095 1847
rect 4061 1681 4095 1715
rect 4061 1613 4095 1647
rect 4061 1563 4095 1579
rect 4411 1881 4449 1895
rect 4411 1861 4413 1881
rect 4237 1749 4271 1847
rect 4237 1681 4271 1715
rect 4237 1613 4271 1647
rect 4237 1563 4271 1579
rect 4447 1861 4449 1881
rect 4589 1881 4623 1915
rect 4765 2017 4799 2033
rect 4765 1949 4799 1983
rect 4765 1895 4799 1915
rect 4941 2017 4975 2033
rect 4941 1949 4975 1983
rect 4413 1749 4447 1847
rect 4763 1881 4801 1895
rect 4763 1861 4765 1881
rect 4589 1749 4623 1847
rect 4413 1681 4447 1715
rect 4587 1715 4589 1744
rect 4799 1861 4801 1881
rect 4941 1881 4975 1915
rect 5117 2017 5151 2033
rect 5117 1949 5151 1983
rect 5117 1895 5151 1915
rect 5293 2017 5327 2033
rect 5293 1949 5327 1983
rect 4765 1749 4799 1847
rect 4623 1715 4625 1744
rect 4587 1710 4625 1715
rect 5115 1881 5153 1895
rect 5115 1861 5117 1881
rect 4941 1749 4975 1847
rect 4413 1613 4447 1647
rect 4413 1563 4447 1579
rect 4589 1681 4623 1710
rect 4589 1613 4623 1647
rect 4589 1563 4623 1579
rect 4765 1681 4799 1715
rect 4939 1715 4941 1744
rect 5151 1861 5153 1881
rect 5293 1881 5327 1915
rect 5469 2017 5503 2033
rect 5469 1949 5503 1983
rect 5469 1895 5503 1915
rect 5645 2017 5679 2033
rect 5645 1949 5679 1983
rect 5117 1749 5151 1847
rect 4975 1715 4977 1744
rect 4939 1710 4977 1715
rect 5467 1881 5505 1895
rect 5467 1861 5469 1881
rect 5293 1749 5327 1847
rect 4765 1613 4799 1647
rect 4765 1563 4799 1579
rect 4941 1681 4975 1710
rect 4941 1613 4975 1647
rect 4941 1563 4975 1579
rect 5117 1681 5151 1715
rect 5291 1715 5293 1744
rect 5503 1861 5505 1881
rect 5645 1881 5679 1915
rect 5821 2017 5855 2033
rect 5821 1949 5855 1983
rect 5821 1895 5855 1915
rect 5469 1749 5503 1847
rect 5327 1715 5329 1744
rect 5291 1710 5329 1715
rect 5783 1861 5821 1895
rect 5645 1749 5679 1847
rect 5117 1613 5151 1647
rect 5117 1563 5151 1579
rect 5293 1681 5327 1710
rect 5293 1613 5327 1647
rect 5293 1563 5327 1579
rect 5469 1681 5503 1715
rect 5607 1710 5645 1744
rect 5469 1613 5503 1647
rect 5469 1563 5503 1579
rect 5645 1681 5679 1710
rect 5645 1613 5679 1647
rect 5645 1563 5679 1579
rect 5821 1749 5855 1847
rect 5821 1681 5855 1715
rect 5821 1613 5855 1647
rect 5821 1563 5855 1579
rect 3068 1452 3084 1486
rect 3123 1452 3153 1486
rect 3197 1452 3222 1486
rect 3271 1452 3291 1486
rect 3344 1452 3360 1486
rect 3417 1452 3429 1486
rect 3490 1452 3498 1486
rect 3563 1452 3567 1486
rect 3601 1452 3602 1486
rect 3670 1452 3675 1486
rect 3739 1452 3748 1486
rect 3808 1452 3821 1486
rect 3877 1452 3894 1486
rect 3946 1452 3967 1486
rect 4015 1452 4040 1486
rect 4084 1452 4113 1486
rect 4154 1452 4186 1486
rect 4224 1452 4259 1486
rect 4294 1452 4330 1486
rect 4366 1452 4380 1486
rect 4566 1452 4582 1486
rect 4616 1452 4651 1486
rect 4691 1452 4720 1486
rect 4763 1452 4789 1486
rect 4823 1452 4858 1486
rect 4892 1452 4926 1486
rect 4960 1452 4994 1486
rect 5028 1452 5062 1486
rect 5128 1452 5130 1486
rect 5164 1452 5167 1486
rect 5232 1452 5240 1486
rect 5300 1452 5313 1486
rect 5368 1452 5386 1486
rect 5436 1452 5459 1486
rect 5504 1452 5531 1486
rect 5572 1452 5603 1486
rect 5640 1452 5674 1486
rect 5709 1452 5742 1486
rect 5781 1452 5792 1486
rect 3005 1357 3039 1373
rect 3179 1358 3217 1392
rect 3005 1312 3039 1323
rect 3005 1240 3039 1255
rect 3181 1357 3215 1358
rect 3181 1289 3215 1323
rect 3181 1239 3215 1255
rect 3357 1357 3391 1373
rect 3531 1358 3569 1392
rect 3357 1312 3391 1323
rect 3357 1240 3391 1255
rect 3533 1357 3567 1358
rect 3533 1289 3567 1323
rect 3533 1239 3567 1255
rect 3709 1357 3743 1373
rect 3883 1358 3921 1392
rect 3709 1312 3743 1323
rect 3709 1240 3743 1255
rect 3885 1357 3919 1358
rect 3885 1289 3919 1323
rect 3885 1239 3919 1255
rect 4061 1357 4095 1373
rect 4235 1358 4273 1392
rect 4061 1312 4095 1323
rect 4061 1240 4095 1255
rect 4237 1357 4271 1358
rect 4237 1289 4271 1323
rect 4237 1239 4271 1255
rect 4413 1357 4447 1373
rect 4587 1358 4625 1392
rect 4413 1312 4447 1323
rect 4413 1240 4447 1255
rect 4589 1357 4623 1358
rect 4589 1289 4623 1323
rect 4589 1239 4623 1255
rect 4765 1357 4799 1373
rect 4939 1358 4977 1392
rect 4765 1312 4799 1323
rect 4765 1240 4799 1255
rect 4941 1357 4975 1358
rect 4941 1289 4975 1323
rect 4941 1239 4975 1255
rect 5117 1357 5151 1373
rect 5291 1358 5329 1392
rect 5117 1312 5151 1323
rect 5117 1240 5151 1255
rect 5293 1357 5327 1358
rect 5293 1289 5327 1323
rect 5293 1239 5327 1255
rect 5469 1357 5503 1373
rect 5643 1358 5681 1392
rect 5469 1312 5503 1323
rect 5469 1240 5503 1255
rect 5645 1357 5679 1358
rect 5645 1289 5679 1323
rect 5645 1239 5679 1255
rect 5821 1357 5855 1373
rect 5821 1312 5855 1323
rect 5821 1240 5855 1255
<< viali >>
rect 3155 2109 3159 2143
rect 3159 2109 3189 2143
rect 3228 2109 3262 2143
rect 3301 2109 3331 2143
rect 3331 2109 3335 2143
rect 3374 2109 3400 2143
rect 3400 2109 3408 2143
rect 3447 2109 3469 2143
rect 3469 2109 3481 2143
rect 3520 2109 3538 2143
rect 3538 2109 3554 2143
rect 3593 2109 3607 2143
rect 3607 2109 3627 2143
rect 3666 2109 3676 2143
rect 3676 2109 3700 2143
rect 3739 2109 3745 2143
rect 3745 2109 3773 2143
rect 3812 2109 3814 2143
rect 3814 2109 3846 2143
rect 3885 2109 3918 2143
rect 3918 2109 3919 2143
rect 3958 2109 3987 2143
rect 3987 2109 3992 2143
rect 4031 2109 4056 2143
rect 4056 2109 4065 2143
rect 4104 2109 4125 2143
rect 4125 2109 4138 2143
rect 4177 2109 4195 2143
rect 4195 2109 4211 2143
rect 4250 2109 4265 2143
rect 4265 2109 4284 2143
rect 4324 2109 4335 2143
rect 4335 2109 4358 2143
rect 4398 2109 4405 2143
rect 4405 2109 4432 2143
rect 4472 2109 4475 2143
rect 4475 2109 4506 2143
rect 4546 2109 4579 2143
rect 4579 2109 4580 2143
rect 4620 2109 4649 2143
rect 4649 2109 4654 2143
rect 4694 2109 4719 2143
rect 4719 2109 4728 2143
rect 4768 2109 4789 2143
rect 4789 2109 4802 2143
rect 4842 2109 4859 2143
rect 4859 2109 4876 2143
rect 4916 2109 4929 2143
rect 4929 2109 4950 2143
rect 4990 2109 4999 2143
rect 4999 2109 5024 2143
rect 5064 2109 5069 2143
rect 5069 2109 5098 2143
rect 5138 2109 5139 2143
rect 5139 2109 5172 2143
rect 5212 2109 5245 2143
rect 5245 2109 5246 2143
rect 5286 2109 5315 2143
rect 5315 2109 5320 2143
rect 5360 2109 5385 2143
rect 5385 2109 5394 2143
rect 5434 2109 5455 2143
rect 5455 2109 5468 2143
rect 5508 2109 5525 2143
rect 5525 2109 5542 2143
rect 5582 2109 5595 2143
rect 5595 2109 5616 2143
rect 5656 2109 5665 2143
rect 5665 2109 5690 2143
rect 5730 2109 5735 2143
rect 5735 2109 5764 2143
rect 5804 2109 5805 2143
rect 5805 2109 5838 2143
rect 3181 2029 3215 2063
rect 3181 1983 3215 1991
rect 3181 1957 3215 1983
rect 3006 1881 3040 1895
rect 3006 1861 3039 1881
rect 3039 1861 3040 1881
rect 3078 1861 3112 1895
rect 3533 2029 3567 2063
rect 3533 1983 3567 1991
rect 3533 1957 3567 1983
rect 3321 1861 3355 1895
rect 3393 1861 3427 1895
rect 3885 2029 3919 2063
rect 3885 1983 3919 1991
rect 3885 1957 3919 1983
rect 3673 1861 3707 1895
rect 3745 1861 3779 1895
rect 4237 2029 4271 2063
rect 4237 1983 4271 1991
rect 4237 1957 4271 1983
rect 4025 1861 4059 1895
rect 4097 1861 4131 1895
rect 4377 1861 4411 1895
rect 4449 1861 4483 1895
rect 4729 1861 4763 1895
rect 4553 1710 4587 1744
rect 4801 1861 4835 1895
rect 4625 1710 4659 1744
rect 5081 1861 5115 1895
rect 4905 1710 4939 1744
rect 5153 1861 5187 1895
rect 4977 1710 5011 1744
rect 5433 1861 5467 1895
rect 5257 1710 5291 1744
rect 5505 1861 5539 1895
rect 5329 1710 5363 1744
rect 5749 1861 5783 1895
rect 5821 1881 5855 1895
rect 5821 1861 5855 1881
rect 5573 1710 5607 1744
rect 5645 1715 5679 1744
rect 5645 1710 5679 1715
rect 3089 1452 3118 1486
rect 3118 1452 3123 1486
rect 3163 1452 3187 1486
rect 3187 1452 3197 1486
rect 3237 1452 3256 1486
rect 3256 1452 3271 1486
rect 3310 1452 3325 1486
rect 3325 1452 3344 1486
rect 3383 1452 3394 1486
rect 3394 1452 3417 1486
rect 3456 1452 3463 1486
rect 3463 1452 3490 1486
rect 3529 1452 3532 1486
rect 3532 1452 3563 1486
rect 3602 1452 3636 1486
rect 3675 1452 3705 1486
rect 3705 1452 3709 1486
rect 3748 1452 3774 1486
rect 3774 1452 3782 1486
rect 3821 1452 3843 1486
rect 3843 1452 3855 1486
rect 3894 1452 3912 1486
rect 3912 1452 3928 1486
rect 3967 1452 3981 1486
rect 3981 1452 4001 1486
rect 4040 1452 4050 1486
rect 4050 1452 4074 1486
rect 4113 1452 4120 1486
rect 4120 1452 4147 1486
rect 4186 1452 4190 1486
rect 4190 1452 4220 1486
rect 4259 1452 4260 1486
rect 4260 1452 4293 1486
rect 4332 1452 4364 1486
rect 4364 1452 4366 1486
rect 4657 1452 4685 1486
rect 4685 1452 4691 1486
rect 4729 1452 4754 1486
rect 4754 1452 4763 1486
rect 5094 1452 5096 1486
rect 5096 1452 5128 1486
rect 5167 1452 5198 1486
rect 5198 1452 5201 1486
rect 5240 1452 5266 1486
rect 5266 1452 5274 1486
rect 5313 1452 5334 1486
rect 5334 1452 5347 1486
rect 5386 1452 5402 1486
rect 5402 1452 5420 1486
rect 5459 1452 5470 1486
rect 5470 1452 5493 1486
rect 5531 1452 5538 1486
rect 5538 1452 5565 1486
rect 5603 1452 5606 1486
rect 5606 1452 5637 1486
rect 5675 1452 5708 1486
rect 5708 1452 5709 1486
rect 5747 1452 5776 1486
rect 5776 1452 5781 1486
rect 3145 1358 3179 1392
rect 3217 1358 3251 1392
rect 3005 1289 3039 1312
rect 3005 1278 3039 1289
rect 3005 1206 3039 1240
rect 3497 1358 3531 1392
rect 3569 1358 3603 1392
rect 3357 1289 3391 1312
rect 3357 1278 3391 1289
rect 3357 1206 3391 1240
rect 3849 1358 3883 1392
rect 3921 1358 3955 1392
rect 3709 1289 3743 1312
rect 3709 1278 3743 1289
rect 3709 1206 3743 1240
rect 4201 1358 4235 1392
rect 4273 1358 4307 1392
rect 4061 1289 4095 1312
rect 4061 1278 4095 1289
rect 4061 1206 4095 1240
rect 4553 1358 4587 1392
rect 4625 1358 4659 1392
rect 4413 1289 4447 1312
rect 4413 1278 4447 1289
rect 4413 1206 4447 1240
rect 4905 1358 4939 1392
rect 4977 1358 5011 1392
rect 4765 1289 4799 1312
rect 4765 1278 4799 1289
rect 4765 1206 4799 1240
rect 5257 1358 5291 1392
rect 5329 1358 5363 1392
rect 5117 1289 5151 1312
rect 5117 1278 5151 1289
rect 5117 1206 5151 1240
rect 5609 1358 5643 1392
rect 5681 1358 5715 1392
rect 5469 1289 5503 1312
rect 5469 1278 5503 1289
rect 5469 1206 5503 1240
rect 5821 1289 5855 1312
rect 5821 1278 5855 1289
rect 5821 1206 5855 1240
<< metal1 >>
rect 3143 2143 5850 2149
rect 3143 2109 3155 2143
rect 3189 2109 3228 2143
rect 3262 2109 3301 2143
rect 3335 2109 3374 2143
rect 3408 2109 3447 2143
rect 3481 2109 3520 2143
rect 3554 2109 3593 2143
rect 3627 2109 3666 2143
rect 3700 2109 3739 2143
rect 3773 2109 3812 2143
rect 3846 2109 3885 2143
rect 3919 2109 3958 2143
rect 3992 2109 4031 2143
rect 4065 2109 4104 2143
rect 4138 2109 4177 2143
rect 4211 2109 4250 2143
rect 4284 2109 4324 2143
rect 4358 2109 4398 2143
rect 4432 2109 4472 2143
rect 4506 2109 4546 2143
rect 4580 2109 4620 2143
rect 4654 2109 4694 2143
rect 4728 2109 4768 2143
rect 4802 2109 4842 2143
rect 4876 2109 4916 2143
rect 4950 2109 4990 2143
rect 5024 2109 5064 2143
rect 5098 2109 5138 2143
rect 5172 2109 5212 2143
rect 5246 2109 5286 2143
rect 5320 2109 5360 2143
rect 5394 2109 5434 2143
rect 5468 2109 5508 2143
rect 5542 2109 5582 2143
rect 5616 2109 5656 2143
rect 5690 2109 5730 2143
rect 5764 2109 5804 2143
rect 5838 2109 5850 2143
rect 3143 2063 5850 2109
rect 3143 2029 3181 2063
rect 3215 2029 3533 2063
rect 3567 2029 3885 2063
rect 3919 2029 4237 2063
rect 4271 2029 5850 2063
rect 3143 1991 5850 2029
rect 3143 1957 3181 1991
rect 3215 1957 3533 1991
rect 3567 1957 3885 1991
rect 3919 1957 4237 1991
rect 4271 1957 5850 1991
rect 3143 1944 5850 1957
rect 2994 1895 5867 1901
rect 2994 1861 3006 1895
rect 3040 1861 3078 1895
rect 3112 1861 3321 1895
rect 3355 1861 3393 1895
rect 3427 1861 3673 1895
rect 3707 1861 3745 1895
rect 3779 1861 4025 1895
rect 4059 1861 4097 1895
rect 4131 1861 4377 1895
rect 4411 1861 4449 1895
rect 4483 1861 4729 1895
rect 4763 1861 4801 1895
rect 4835 1861 5081 1895
rect 5115 1861 5153 1895
rect 5187 1861 5433 1895
rect 5467 1861 5505 1895
rect 5539 1861 5749 1895
rect 5783 1861 5821 1895
rect 5855 1861 5867 1895
rect 2994 1855 5867 1861
rect 4541 1744 5691 1750
rect 4541 1710 4553 1744
rect 4587 1710 4625 1744
rect 4659 1710 4905 1744
rect 4939 1710 4977 1744
rect 5011 1710 5257 1744
rect 5291 1710 5329 1744
rect 5363 1710 5573 1744
rect 5607 1710 5645 1744
rect 5679 1710 5691 1744
rect 4541 1704 5691 1710
rect 3077 1486 4378 1492
rect 3077 1452 3089 1486
rect 3123 1452 3163 1486
rect 3197 1452 3237 1486
rect 3271 1452 3310 1486
rect 3344 1452 3383 1486
rect 3417 1452 3456 1486
rect 3490 1452 3529 1486
rect 3563 1452 3602 1486
rect 3636 1452 3675 1486
rect 3709 1452 3748 1486
rect 3782 1452 3821 1486
rect 3855 1452 3894 1486
rect 3928 1452 3967 1486
rect 4001 1452 4040 1486
rect 4074 1452 4113 1486
rect 4147 1452 4186 1486
rect 4220 1452 4259 1486
rect 4293 1452 4332 1486
rect 4366 1452 4378 1486
rect 3077 1446 4378 1452
rect 4645 1486 4775 1492
rect 4645 1452 4657 1486
rect 4691 1452 4729 1486
rect 4763 1452 4775 1486
rect 4645 1446 4775 1452
rect 4893 1398 5023 1704
rect 5082 1486 5793 1492
rect 5082 1452 5094 1486
rect 5128 1452 5167 1486
rect 5201 1452 5240 1486
rect 5274 1452 5313 1486
rect 5347 1452 5386 1486
rect 5420 1452 5459 1486
rect 5493 1452 5531 1486
rect 5565 1452 5603 1486
rect 5637 1452 5675 1486
rect 5709 1452 5747 1486
rect 5781 1452 5793 1486
rect 5082 1446 5793 1452
rect 3133 1392 5727 1398
rect 3133 1358 3145 1392
rect 3179 1358 3217 1392
rect 3251 1358 3497 1392
rect 3531 1358 3569 1392
rect 3603 1358 3849 1392
rect 3883 1358 3921 1392
rect 3955 1358 4201 1392
rect 4235 1358 4273 1392
rect 4307 1358 4553 1392
rect 4587 1358 4625 1392
rect 4659 1358 4905 1392
rect 4939 1358 4977 1392
rect 5011 1358 5257 1392
rect 5291 1358 5329 1392
rect 5363 1358 5609 1392
rect 5643 1358 5681 1392
rect 5715 1358 5727 1392
rect 3133 1352 5727 1358
rect 2999 1312 5861 1324
rect 2999 1278 3005 1312
rect 3039 1278 3357 1312
rect 3391 1278 3709 1312
rect 3743 1278 4061 1312
rect 4095 1278 4413 1312
rect 4447 1278 4765 1312
rect 4799 1278 5117 1312
rect 5151 1278 5469 1312
rect 5503 1278 5821 1312
rect 5855 1278 5861 1312
rect 2999 1240 5861 1278
rect 2999 1206 3005 1240
rect 3039 1206 3357 1240
rect 3391 1206 3709 1240
rect 3743 1206 4061 1240
rect 4095 1206 4413 1240
rect 4447 1206 4765 1240
rect 4799 1206 5117 1240
rect 5151 1206 5469 1240
rect 5503 1206 5821 1240
rect 5855 1206 5861 1240
rect 2999 1109 5861 1206
use sky130_fd_pr__model__nfet_highvoltage__example_55959141808442  sky130_fd_pr__model__nfet_highvoltage__example_55959141808442_0
timestamp 1666464484
transform 1 0 3050 0 -1 1369
box -1 0 2761 1
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808443  sky130_fd_pr__model__pfet_highvoltage__example_55959141808443_0
timestamp 1666464484
transform 1 0 3050 0 1 1835
box -1 0 2761 1
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808443  sky130_fd_pr__model__pfet_highvoltage__example_55959141808443_1
timestamp 1666464484
transform 1 0 3050 0 1 1567
box -1 0 2761 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1666464484
transform -1 0 4763 0 -1 1486
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_1
timestamp 1666464484
transform -1 0 5011 0 -1 1744
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_2
timestamp 1666464484
transform -1 0 4659 0 -1 1744
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_3
timestamp 1666464484
transform -1 0 5363 0 -1 1744
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_4
timestamp 1666464484
transform -1 0 4307 0 -1 1392
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_5
timestamp 1666464484
transform -1 0 3955 0 -1 1392
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_6
timestamp 1666464484
transform -1 0 3251 0 -1 1392
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_7
timestamp 1666464484
transform -1 0 3603 0 -1 1392
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_8
timestamp 1666464484
transform -1 0 5679 0 -1 1744
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_9
timestamp 1666464484
transform -1 0 5011 0 -1 1392
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_10
timestamp 1666464484
transform 0 -1 3039 -1 0 1312
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_11
timestamp 1666464484
transform -1 0 4659 0 -1 1392
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_12
timestamp 1666464484
transform -1 0 5363 0 -1 1392
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_13
timestamp 1666464484
transform -1 0 5715 0 -1 1392
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_14
timestamp 1666464484
transform -1 0 5855 0 -1 1895
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_15
timestamp 1666464484
transform -1 0 5539 0 -1 1895
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_16
timestamp 1666464484
transform -1 0 4835 0 -1 1895
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_17
timestamp 1666464484
transform -1 0 5187 0 -1 1895
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_18
timestamp 1666464484
transform -1 0 3112 0 -1 1895
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_19
timestamp 1666464484
transform -1 0 3779 0 -1 1895
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_20
timestamp 1666464484
transform -1 0 3427 0 -1 1895
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_21
timestamp 1666464484
transform -1 0 4131 0 -1 1895
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_22
timestamp 1666464484
transform -1 0 4483 0 -1 1895
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_23
timestamp 1666464484
transform 0 -1 5503 -1 0 1312
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_24
timestamp 1666464484
transform 0 -1 5855 -1 0 1312
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_25
timestamp 1666464484
transform 0 -1 3391 -1 0 1312
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_26
timestamp 1666464484
transform 0 -1 5151 -1 0 1312
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_27
timestamp 1666464484
transform 0 -1 4095 -1 0 1312
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_28
timestamp 1666464484
transform 0 -1 3743 -1 0 1312
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_29
timestamp 1666464484
transform 0 -1 4447 -1 0 1312
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_30
timestamp 1666464484
transform 0 -1 4271 1 0 1957
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_31
timestamp 1666464484
transform 0 -1 4799 -1 0 1312
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_32
timestamp 1666464484
transform 0 -1 3919 1 0 1957
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_33
timestamp 1666464484
transform 0 -1 3567 1 0 1957
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_34
timestamp 1666464484
transform 0 -1 3215 1 0 1957
box 0 0 1 1
<< labels >>
flabel metal1 s 4132 1456 4173 1477 3 FreeSans 520 0 0 0 IN0
port 1 nsew
flabel metal1 s 4685 1456 4734 1480 3 FreeSans 520 0 0 0 IN1
port 2 nsew
flabel metal1 s 4083 1157 4209 1270 3 FreeSans 520 0 0 0 VGND
port 3 nsew
flabel metal1 s 3973 2003 4147 2113 3 FreeSans 520 0 0 0 VPWR
port 4 nsew
flabel metal1 s 4928 1717 4971 1742 3 FreeSans 520 0 0 0 OUT
port 5 nsew
<< properties >>
string GDS_END 31873064
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 31855706
<< end >>
