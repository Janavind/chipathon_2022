magic
tech sky130A
magscale 1 2
timestamp 1666199351
<< dnwell >>
rect 1043 23645 8429 24789
rect 1043 21838 17881 23645
rect 14472 21038 17881 21838
rect 17434 20964 17881 21038
<< nwell >>
rect 963 24583 8509 24869
rect 963 22044 1249 24583
rect 8223 23725 8509 24583
rect 8223 23439 17961 23725
rect 963 21758 2317 22044
rect 17675 21170 17961 23439
rect 17434 20884 17961 21170
rect 12737 457 12971 691
<< pwell >>
rect 17194 23353 17280 23362
rect 15384 21253 17280 23353
rect 15384 21247 17142 21253
<< mvnmos >>
rect 15463 23243 17063 23327
rect 15463 23041 17063 23125
rect 15463 22881 17063 22965
rect 15463 22679 17063 22763
rect 15463 22519 17063 22603
rect 15463 22359 17063 22443
rect 15463 22157 17063 22241
rect 15463 21997 17063 22081
rect 15463 21837 17063 21921
rect 15463 21635 17063 21719
rect 15463 21475 17063 21559
rect 15463 21273 17063 21357
<< mvndiff >>
rect 15410 23315 15463 23327
rect 15410 23281 15418 23315
rect 15452 23281 15463 23315
rect 15410 23243 15463 23281
rect 17063 23315 17116 23327
rect 17063 23281 17074 23315
rect 17108 23281 17116 23315
rect 17063 23243 17116 23281
rect 15410 23113 15463 23125
rect 15410 23079 15418 23113
rect 15452 23079 15463 23113
rect 15410 23041 15463 23079
rect 17063 23113 17116 23125
rect 17063 23079 17074 23113
rect 17108 23079 17116 23113
rect 17063 23041 17116 23079
rect 15410 22953 15463 22965
rect 15410 22919 15418 22953
rect 15452 22919 15463 22953
rect 15410 22881 15463 22919
rect 17063 22953 17116 22965
rect 17063 22919 17074 22953
rect 17108 22919 17116 22953
rect 17063 22881 17116 22919
rect 15410 22751 15463 22763
rect 15410 22717 15418 22751
rect 15452 22717 15463 22751
rect 15410 22679 15463 22717
rect 17063 22751 17116 22763
rect 17063 22717 17074 22751
rect 17108 22717 17116 22751
rect 17063 22679 17116 22717
rect 15410 22591 15463 22603
rect 15410 22557 15418 22591
rect 15452 22557 15463 22591
rect 15410 22519 15463 22557
rect 17063 22591 17116 22603
rect 17063 22557 17074 22591
rect 17108 22557 17116 22591
rect 17063 22519 17116 22557
rect 15410 22431 15463 22443
rect 15410 22397 15418 22431
rect 15452 22397 15463 22431
rect 15410 22359 15463 22397
rect 17063 22431 17116 22443
rect 17063 22397 17074 22431
rect 17108 22397 17116 22431
rect 17063 22359 17116 22397
rect 15410 22229 15463 22241
rect 15410 22195 15418 22229
rect 15452 22195 15463 22229
rect 15410 22157 15463 22195
rect 17063 22229 17116 22241
rect 17063 22195 17074 22229
rect 17108 22195 17116 22229
rect 17063 22157 17116 22195
rect 15410 22069 15463 22081
rect 15410 22035 15418 22069
rect 15452 22035 15463 22069
rect 15410 21997 15463 22035
rect 17063 22069 17116 22081
rect 17063 22035 17074 22069
rect 17108 22035 17116 22069
rect 17063 21997 17116 22035
rect 15410 21909 15463 21921
rect 15410 21875 15418 21909
rect 15452 21875 15463 21909
rect 15410 21837 15463 21875
rect 17063 21909 17116 21921
rect 17063 21875 17074 21909
rect 17108 21875 17116 21909
rect 17063 21837 17116 21875
rect 15410 21707 15463 21719
rect 15410 21673 15418 21707
rect 15452 21673 15463 21707
rect 15410 21635 15463 21673
rect 17063 21707 17116 21719
rect 17063 21673 17074 21707
rect 17108 21673 17116 21707
rect 17063 21635 17116 21673
rect 15410 21547 15463 21559
rect 15410 21513 15418 21547
rect 15452 21513 15463 21547
rect 15410 21475 15463 21513
rect 17063 21547 17116 21559
rect 17063 21513 17074 21547
rect 17108 21513 17116 21547
rect 17063 21475 17116 21513
rect 15410 21345 15463 21357
rect 15410 21311 15418 21345
rect 15452 21311 15463 21345
rect 15410 21273 15463 21311
rect 17063 21345 17116 21357
rect 17063 21311 17074 21345
rect 17108 21311 17116 21345
rect 17063 21273 17116 21311
<< mvndiffc >>
rect 15418 23281 15452 23315
rect 17074 23281 17108 23315
rect 15418 23079 15452 23113
rect 17074 23079 17108 23113
rect 15418 22919 15452 22953
rect 17074 22919 17108 22953
rect 15418 22717 15452 22751
rect 17074 22717 17108 22751
rect 15418 22557 15452 22591
rect 17074 22557 17108 22591
rect 15418 22397 15452 22431
rect 17074 22397 17108 22431
rect 15418 22195 15452 22229
rect 17074 22195 17108 22229
rect 15418 22035 15452 22069
rect 17074 22035 17108 22069
rect 15418 21875 15452 21909
rect 17074 21875 17108 21909
rect 15418 21673 15452 21707
rect 17074 21673 17108 21707
rect 15418 21513 15452 21547
rect 17074 21513 17108 21547
rect 15418 21311 15452 21345
rect 17074 21311 17108 21345
<< mvpsubdiff >>
rect 17220 23302 17254 23336
rect 17220 23217 17254 23268
rect 17220 23132 17254 23183
rect 17220 23047 17254 23098
rect 17220 22962 17254 23013
rect 17220 22877 17254 22928
rect 17220 22792 17254 22843
rect 17220 22707 17254 22758
rect 17220 22622 17254 22673
rect 17220 22537 17254 22588
rect 17220 22452 17254 22503
rect 17220 22367 17254 22418
rect 17220 22282 17254 22333
rect 17220 22197 17254 22248
rect 17220 22112 17254 22163
rect 17220 22027 17254 22078
rect 17220 21942 17254 21993
rect 17220 21857 17254 21908
rect 17220 21772 17254 21823
rect 17220 21687 17254 21738
rect 17220 21602 17254 21653
rect 17220 21517 17254 21568
rect 17220 21432 17254 21483
rect 17220 21347 17254 21398
rect 17220 21279 17254 21313
<< mvnsubdiff >>
rect 1089 24709 1209 24743
rect 1243 24709 1277 24743
rect 1311 24709 1345 24743
rect 1379 24709 1413 24743
rect 1447 24709 1481 24743
rect 1515 24709 1549 24743
rect 1583 24709 1617 24743
rect 1651 24709 1685 24743
rect 1719 24709 1753 24743
rect 1787 24709 1821 24743
rect 1855 24709 1889 24743
rect 1923 24709 1957 24743
rect 1991 24709 2025 24743
rect 2059 24709 2093 24743
rect 2127 24709 2161 24743
rect 2195 24709 2229 24743
rect 2263 24709 2297 24743
rect 2331 24709 2365 24743
rect 2399 24709 2433 24743
rect 2467 24709 2501 24743
rect 2535 24709 2569 24743
rect 2603 24709 2637 24743
rect 2671 24709 2705 24743
rect 2739 24709 2773 24743
rect 2807 24709 2841 24743
rect 2875 24709 2909 24743
rect 2943 24709 2977 24743
rect 3011 24709 3045 24743
rect 3079 24709 3113 24743
rect 3147 24709 3181 24743
rect 3215 24709 3249 24743
rect 3283 24709 3317 24743
rect 3351 24709 3385 24743
rect 3419 24709 3453 24743
rect 3487 24709 3521 24743
rect 3555 24709 3589 24743
rect 3623 24709 3657 24743
rect 3691 24709 3725 24743
rect 3759 24709 3793 24743
rect 3827 24709 3861 24743
rect 3895 24709 3929 24743
rect 3963 24709 3997 24743
rect 4031 24709 4065 24743
rect 4099 24709 4133 24743
rect 4167 24709 4201 24743
rect 4235 24709 4269 24743
rect 4303 24709 4337 24743
rect 4371 24709 4405 24743
rect 4439 24709 4473 24743
rect 4507 24709 4541 24743
rect 4575 24709 4609 24743
rect 4643 24709 4677 24743
rect 4711 24709 4745 24743
rect 4779 24709 4813 24743
rect 4847 24709 4881 24743
rect 4915 24709 4949 24743
rect 4983 24709 5017 24743
rect 5051 24709 5085 24743
rect 5119 24709 5153 24743
rect 5187 24709 5221 24743
rect 5255 24709 5289 24743
rect 5323 24709 5357 24743
rect 5391 24709 5425 24743
rect 5459 24709 5493 24743
rect 5527 24709 5561 24743
rect 5595 24709 5629 24743
rect 5663 24709 5697 24743
rect 5731 24709 5765 24743
rect 5799 24709 5833 24743
rect 5867 24709 5901 24743
rect 5935 24709 5969 24743
rect 6003 24709 6037 24743
rect 6071 24709 6105 24743
rect 6139 24709 6173 24743
rect 6207 24709 6241 24743
rect 6275 24709 6309 24743
rect 6343 24709 6377 24743
rect 6411 24709 6445 24743
rect 6479 24709 6513 24743
rect 6547 24709 6581 24743
rect 6615 24709 6649 24743
rect 6683 24709 6717 24743
rect 6751 24709 6785 24743
rect 6819 24709 6853 24743
rect 6887 24709 6921 24743
rect 6955 24709 6989 24743
rect 7023 24709 7057 24743
rect 7091 24709 7125 24743
rect 7159 24709 7193 24743
rect 7227 24709 7261 24743
rect 7295 24709 7329 24743
rect 7363 24709 7397 24743
rect 7431 24709 7465 24743
rect 7499 24709 7533 24743
rect 7567 24709 7601 24743
rect 7635 24709 7669 24743
rect 7703 24709 7737 24743
rect 7771 24709 7805 24743
rect 7839 24709 7873 24743
rect 7907 24709 7941 24743
rect 7975 24709 8009 24743
rect 8043 24709 8077 24743
rect 8111 24709 8145 24743
rect 8179 24709 8213 24743
rect 8247 24709 8281 24743
rect 8315 24709 8383 24743
rect 1089 24675 1123 24709
rect 1089 24607 1123 24641
rect 1089 24539 1123 24573
rect 1089 24471 1123 24505
rect 1089 24403 1123 24437
rect 1089 24335 1123 24369
rect 1089 24267 1123 24301
rect 1089 24199 1123 24233
rect 1089 24131 1123 24165
rect 1089 24063 1123 24097
rect 1089 23995 1123 24029
rect 1089 23927 1123 23961
rect 1089 23859 1123 23893
rect 1089 23791 1123 23825
rect 1089 23723 1123 23757
rect 1089 23655 1123 23689
rect 1089 23587 1123 23621
rect 8349 24619 8383 24709
rect 8349 24551 8383 24585
rect 8349 24483 8383 24517
rect 8349 24415 8383 24449
rect 8349 24347 8383 24381
rect 8349 24279 8383 24313
rect 8349 24211 8383 24245
rect 8349 24143 8383 24177
rect 8349 24075 8383 24109
rect 8349 24007 8383 24041
rect 8349 23939 8383 23973
rect 8349 23871 8383 23905
rect 8349 23803 8383 23837
rect 8349 23735 8383 23769
rect 8349 23667 8383 23701
rect 8349 23599 8383 23633
rect 8349 23565 8417 23599
rect 8451 23565 8485 23599
rect 8519 23565 8553 23599
rect 8587 23565 8621 23599
rect 8655 23565 8689 23599
rect 8723 23565 8757 23599
rect 8791 23565 8825 23599
rect 8859 23565 8893 23599
rect 8927 23565 8961 23599
rect 8995 23565 9029 23599
rect 9063 23565 9097 23599
rect 9131 23565 9165 23599
rect 9199 23565 9233 23599
rect 9267 23565 9301 23599
rect 9335 23565 9369 23599
rect 9403 23565 9437 23599
rect 9471 23565 9505 23599
rect 9539 23565 9573 23599
rect 9607 23565 9641 23599
rect 9675 23565 9709 23599
rect 9743 23565 9777 23599
rect 9811 23565 9845 23599
rect 9879 23565 9913 23599
rect 9947 23565 9981 23599
rect 10015 23565 10049 23599
rect 10083 23565 10117 23599
rect 10151 23565 10185 23599
rect 10219 23565 10253 23599
rect 10287 23565 10321 23599
rect 10355 23565 10389 23599
rect 10423 23565 10457 23599
rect 10491 23565 10525 23599
rect 10559 23565 10593 23599
rect 10627 23565 10661 23599
rect 10695 23565 10729 23599
rect 10763 23565 10797 23599
rect 10831 23565 10865 23599
rect 10899 23565 10933 23599
rect 10967 23565 11001 23599
rect 11035 23565 11069 23599
rect 11103 23565 11137 23599
rect 11171 23565 11205 23599
rect 11239 23565 11273 23599
rect 11307 23565 11341 23599
rect 11375 23565 11409 23599
rect 11443 23565 11477 23599
rect 11511 23565 11545 23599
rect 11579 23565 11613 23599
rect 11647 23565 11681 23599
rect 11715 23565 11749 23599
rect 11783 23565 11817 23599
rect 11851 23565 11885 23599
rect 11919 23565 11953 23599
rect 11987 23565 12021 23599
rect 12055 23565 12089 23599
rect 12123 23565 12157 23599
rect 12191 23565 12225 23599
rect 12259 23565 12293 23599
rect 12327 23565 12361 23599
rect 12395 23565 12429 23599
rect 12463 23565 12497 23599
rect 12531 23565 12565 23599
rect 12599 23565 12633 23599
rect 12667 23565 12701 23599
rect 12735 23565 12769 23599
rect 12803 23565 12837 23599
rect 12871 23565 12905 23599
rect 12939 23565 12973 23599
rect 13007 23565 13041 23599
rect 13075 23565 13109 23599
rect 13143 23565 13177 23599
rect 13211 23565 13245 23599
rect 13279 23565 13313 23599
rect 13347 23565 13381 23599
rect 13415 23565 13449 23599
rect 13483 23565 13517 23599
rect 13551 23565 13585 23599
rect 13619 23565 13653 23599
rect 13687 23565 13721 23599
rect 13755 23565 13789 23599
rect 13823 23565 13857 23599
rect 13891 23565 13925 23599
rect 13959 23565 13993 23599
rect 14027 23565 14061 23599
rect 14095 23565 14129 23599
rect 14163 23565 14197 23599
rect 14231 23565 14265 23599
rect 14299 23565 14333 23599
rect 14367 23565 14401 23599
rect 14435 23565 14469 23599
rect 14503 23565 14537 23599
rect 14571 23565 14605 23599
rect 14639 23565 14673 23599
rect 14707 23565 14741 23599
rect 14775 23565 14809 23599
rect 14843 23565 14877 23599
rect 14911 23565 14945 23599
rect 14979 23565 15013 23599
rect 15047 23565 15081 23599
rect 15115 23565 15149 23599
rect 15183 23565 15217 23599
rect 15251 23565 15285 23599
rect 15319 23565 15353 23599
rect 15387 23565 15421 23599
rect 15455 23565 15489 23599
rect 15523 23565 15557 23599
rect 15591 23565 15625 23599
rect 15659 23565 15693 23599
rect 15727 23565 15761 23599
rect 15795 23565 15829 23599
rect 15863 23565 15897 23599
rect 15931 23565 15965 23599
rect 15999 23565 16033 23599
rect 16067 23565 16101 23599
rect 16135 23565 16169 23599
rect 16203 23565 16237 23599
rect 16271 23565 16305 23599
rect 16339 23565 16373 23599
rect 16407 23565 16441 23599
rect 16475 23565 16509 23599
rect 16543 23565 16577 23599
rect 16611 23565 16645 23599
rect 16679 23565 16713 23599
rect 16747 23565 16781 23599
rect 16815 23565 16849 23599
rect 16883 23565 16917 23599
rect 16951 23565 16985 23599
rect 17019 23565 17053 23599
rect 17087 23565 17121 23599
rect 17155 23565 17189 23599
rect 17223 23565 17257 23599
rect 17291 23565 17325 23599
rect 17359 23565 17393 23599
rect 17427 23565 17461 23599
rect 17495 23565 17529 23599
rect 17563 23565 17597 23599
rect 17631 23565 17665 23599
rect 17699 23565 17733 23599
rect 17767 23565 17835 23599
rect 1089 23519 1123 23553
rect 1089 23451 1123 23485
rect 1089 23383 1123 23417
rect 17801 23492 17835 23565
rect 17801 23424 17835 23458
rect 17801 23356 17835 23390
rect 1089 23315 1123 23349
rect 1089 23247 1123 23281
rect 1089 23179 1123 23213
rect 1089 23111 1123 23145
rect 1089 23043 1123 23077
rect 1089 22975 1123 23009
rect 1089 22907 1123 22941
rect 1089 22839 1123 22873
rect 1089 22771 1123 22805
rect 1089 22703 1123 22737
rect 1089 22635 1123 22669
rect 1089 22567 1123 22601
rect 1089 22499 1123 22533
rect 1089 22431 1123 22465
rect 1089 22363 1123 22397
rect 1089 22295 1123 22329
rect 1089 22227 1123 22261
rect 1089 22159 1123 22193
rect 1089 22010 1123 22125
rect 1089 21918 1123 21976
rect 1089 21884 1157 21918
rect 1191 21884 1225 21918
rect 1259 21884 1293 21918
rect 1327 21884 1361 21918
rect 1395 21884 1429 21918
rect 1463 21884 1497 21918
rect 1531 21884 1565 21918
rect 1599 21884 1633 21918
rect 1667 21884 1701 21918
rect 1735 21884 1769 21918
rect 1803 21884 1837 21918
rect 1871 21884 1905 21918
rect 1939 21884 1973 21918
rect 2007 21884 2041 21918
rect 2075 21884 2109 21918
rect 2143 21884 2177 21918
rect 2211 21884 2245 21918
rect 2279 21884 2317 21918
rect 17801 23288 17835 23322
rect 17801 23220 17835 23254
rect 17801 23152 17835 23186
rect 17801 23084 17835 23118
rect 17801 23016 17835 23050
rect 17801 22948 17835 22982
rect 17801 22880 17835 22914
rect 17801 22812 17835 22846
rect 17801 22744 17835 22778
rect 17801 22676 17835 22710
rect 17801 22608 17835 22642
rect 17801 22540 17835 22574
rect 17801 22472 17835 22506
rect 17801 22404 17835 22438
rect 17801 22336 17835 22370
rect 17801 22268 17835 22302
rect 17801 22200 17835 22234
rect 17801 22132 17835 22166
rect 17801 22064 17835 22098
rect 17801 21996 17835 22030
rect 17801 21928 17835 21962
rect 17801 21860 17835 21894
rect 17801 21792 17835 21826
rect 17801 21724 17835 21758
rect 17801 21656 17835 21690
rect 17801 21588 17835 21622
rect 17801 21520 17835 21554
rect 17801 21452 17835 21486
rect 17801 21384 17835 21418
rect 17801 21316 17835 21350
rect 17801 21248 17835 21282
rect 17801 21180 17835 21214
rect 17801 21112 17835 21146
rect 17801 21044 17835 21078
rect 17434 21010 17468 21044
rect 17502 21010 17536 21044
rect 17570 21010 17604 21044
rect 17638 21010 17672 21044
rect 17706 21010 17835 21044
rect 12803 581 12905 625
rect 12837 547 12871 581
rect 12803 523 12905 547
<< mvpsubdiffcont >>
rect 17220 23268 17254 23302
rect 17220 23183 17254 23217
rect 17220 23098 17254 23132
rect 17220 23013 17254 23047
rect 17220 22928 17254 22962
rect 17220 22843 17254 22877
rect 17220 22758 17254 22792
rect 17220 22673 17254 22707
rect 17220 22588 17254 22622
rect 17220 22503 17254 22537
rect 17220 22418 17254 22452
rect 17220 22333 17254 22367
rect 17220 22248 17254 22282
rect 17220 22163 17254 22197
rect 17220 22078 17254 22112
rect 17220 21993 17254 22027
rect 17220 21908 17254 21942
rect 17220 21823 17254 21857
rect 17220 21738 17254 21772
rect 17220 21653 17254 21687
rect 17220 21568 17254 21602
rect 17220 21483 17254 21517
rect 17220 21398 17254 21432
rect 17220 21313 17254 21347
<< mvnsubdiffcont >>
rect 1209 24709 1243 24743
rect 1277 24709 1311 24743
rect 1345 24709 1379 24743
rect 1413 24709 1447 24743
rect 1481 24709 1515 24743
rect 1549 24709 1583 24743
rect 1617 24709 1651 24743
rect 1685 24709 1719 24743
rect 1753 24709 1787 24743
rect 1821 24709 1855 24743
rect 1889 24709 1923 24743
rect 1957 24709 1991 24743
rect 2025 24709 2059 24743
rect 2093 24709 2127 24743
rect 2161 24709 2195 24743
rect 2229 24709 2263 24743
rect 2297 24709 2331 24743
rect 2365 24709 2399 24743
rect 2433 24709 2467 24743
rect 2501 24709 2535 24743
rect 2569 24709 2603 24743
rect 2637 24709 2671 24743
rect 2705 24709 2739 24743
rect 2773 24709 2807 24743
rect 2841 24709 2875 24743
rect 2909 24709 2943 24743
rect 2977 24709 3011 24743
rect 3045 24709 3079 24743
rect 3113 24709 3147 24743
rect 3181 24709 3215 24743
rect 3249 24709 3283 24743
rect 3317 24709 3351 24743
rect 3385 24709 3419 24743
rect 3453 24709 3487 24743
rect 3521 24709 3555 24743
rect 3589 24709 3623 24743
rect 3657 24709 3691 24743
rect 3725 24709 3759 24743
rect 3793 24709 3827 24743
rect 3861 24709 3895 24743
rect 3929 24709 3963 24743
rect 3997 24709 4031 24743
rect 4065 24709 4099 24743
rect 4133 24709 4167 24743
rect 4201 24709 4235 24743
rect 4269 24709 4303 24743
rect 4337 24709 4371 24743
rect 4405 24709 4439 24743
rect 4473 24709 4507 24743
rect 4541 24709 4575 24743
rect 4609 24709 4643 24743
rect 4677 24709 4711 24743
rect 4745 24709 4779 24743
rect 4813 24709 4847 24743
rect 4881 24709 4915 24743
rect 4949 24709 4983 24743
rect 5017 24709 5051 24743
rect 5085 24709 5119 24743
rect 5153 24709 5187 24743
rect 5221 24709 5255 24743
rect 5289 24709 5323 24743
rect 5357 24709 5391 24743
rect 5425 24709 5459 24743
rect 5493 24709 5527 24743
rect 5561 24709 5595 24743
rect 5629 24709 5663 24743
rect 5697 24709 5731 24743
rect 5765 24709 5799 24743
rect 5833 24709 5867 24743
rect 5901 24709 5935 24743
rect 5969 24709 6003 24743
rect 6037 24709 6071 24743
rect 6105 24709 6139 24743
rect 6173 24709 6207 24743
rect 6241 24709 6275 24743
rect 6309 24709 6343 24743
rect 6377 24709 6411 24743
rect 6445 24709 6479 24743
rect 6513 24709 6547 24743
rect 6581 24709 6615 24743
rect 6649 24709 6683 24743
rect 6717 24709 6751 24743
rect 6785 24709 6819 24743
rect 6853 24709 6887 24743
rect 6921 24709 6955 24743
rect 6989 24709 7023 24743
rect 7057 24709 7091 24743
rect 7125 24709 7159 24743
rect 7193 24709 7227 24743
rect 7261 24709 7295 24743
rect 7329 24709 7363 24743
rect 7397 24709 7431 24743
rect 7465 24709 7499 24743
rect 7533 24709 7567 24743
rect 7601 24709 7635 24743
rect 7669 24709 7703 24743
rect 7737 24709 7771 24743
rect 7805 24709 7839 24743
rect 7873 24709 7907 24743
rect 7941 24709 7975 24743
rect 8009 24709 8043 24743
rect 8077 24709 8111 24743
rect 8145 24709 8179 24743
rect 8213 24709 8247 24743
rect 8281 24709 8315 24743
rect 1089 24641 1123 24675
rect 1089 24573 1123 24607
rect 1089 24505 1123 24539
rect 1089 24437 1123 24471
rect 1089 24369 1123 24403
rect 1089 24301 1123 24335
rect 1089 24233 1123 24267
rect 1089 24165 1123 24199
rect 1089 24097 1123 24131
rect 1089 24029 1123 24063
rect 1089 23961 1123 23995
rect 1089 23893 1123 23927
rect 1089 23825 1123 23859
rect 1089 23757 1123 23791
rect 1089 23689 1123 23723
rect 1089 23621 1123 23655
rect 1089 23553 1123 23587
rect 8349 24585 8383 24619
rect 8349 24517 8383 24551
rect 8349 24449 8383 24483
rect 8349 24381 8383 24415
rect 8349 24313 8383 24347
rect 8349 24245 8383 24279
rect 8349 24177 8383 24211
rect 8349 24109 8383 24143
rect 8349 24041 8383 24075
rect 8349 23973 8383 24007
rect 8349 23905 8383 23939
rect 8349 23837 8383 23871
rect 8349 23769 8383 23803
rect 8349 23701 8383 23735
rect 8349 23633 8383 23667
rect 8417 23565 8451 23599
rect 8485 23565 8519 23599
rect 8553 23565 8587 23599
rect 8621 23565 8655 23599
rect 8689 23565 8723 23599
rect 8757 23565 8791 23599
rect 8825 23565 8859 23599
rect 8893 23565 8927 23599
rect 8961 23565 8995 23599
rect 9029 23565 9063 23599
rect 9097 23565 9131 23599
rect 9165 23565 9199 23599
rect 9233 23565 9267 23599
rect 9301 23565 9335 23599
rect 9369 23565 9403 23599
rect 9437 23565 9471 23599
rect 9505 23565 9539 23599
rect 9573 23565 9607 23599
rect 9641 23565 9675 23599
rect 9709 23565 9743 23599
rect 9777 23565 9811 23599
rect 9845 23565 9879 23599
rect 9913 23565 9947 23599
rect 9981 23565 10015 23599
rect 10049 23565 10083 23599
rect 10117 23565 10151 23599
rect 10185 23565 10219 23599
rect 10253 23565 10287 23599
rect 10321 23565 10355 23599
rect 10389 23565 10423 23599
rect 10457 23565 10491 23599
rect 10525 23565 10559 23599
rect 10593 23565 10627 23599
rect 10661 23565 10695 23599
rect 10729 23565 10763 23599
rect 10797 23565 10831 23599
rect 10865 23565 10899 23599
rect 10933 23565 10967 23599
rect 11001 23565 11035 23599
rect 11069 23565 11103 23599
rect 11137 23565 11171 23599
rect 11205 23565 11239 23599
rect 11273 23565 11307 23599
rect 11341 23565 11375 23599
rect 11409 23565 11443 23599
rect 11477 23565 11511 23599
rect 11545 23565 11579 23599
rect 11613 23565 11647 23599
rect 11681 23565 11715 23599
rect 11749 23565 11783 23599
rect 11817 23565 11851 23599
rect 11885 23565 11919 23599
rect 11953 23565 11987 23599
rect 12021 23565 12055 23599
rect 12089 23565 12123 23599
rect 12157 23565 12191 23599
rect 12225 23565 12259 23599
rect 12293 23565 12327 23599
rect 12361 23565 12395 23599
rect 12429 23565 12463 23599
rect 12497 23565 12531 23599
rect 12565 23565 12599 23599
rect 12633 23565 12667 23599
rect 12701 23565 12735 23599
rect 12769 23565 12803 23599
rect 12837 23565 12871 23599
rect 12905 23565 12939 23599
rect 12973 23565 13007 23599
rect 13041 23565 13075 23599
rect 13109 23565 13143 23599
rect 13177 23565 13211 23599
rect 13245 23565 13279 23599
rect 13313 23565 13347 23599
rect 13381 23565 13415 23599
rect 13449 23565 13483 23599
rect 13517 23565 13551 23599
rect 13585 23565 13619 23599
rect 13653 23565 13687 23599
rect 13721 23565 13755 23599
rect 13789 23565 13823 23599
rect 13857 23565 13891 23599
rect 13925 23565 13959 23599
rect 13993 23565 14027 23599
rect 14061 23565 14095 23599
rect 14129 23565 14163 23599
rect 14197 23565 14231 23599
rect 14265 23565 14299 23599
rect 14333 23565 14367 23599
rect 14401 23565 14435 23599
rect 14469 23565 14503 23599
rect 14537 23565 14571 23599
rect 14605 23565 14639 23599
rect 14673 23565 14707 23599
rect 14741 23565 14775 23599
rect 14809 23565 14843 23599
rect 14877 23565 14911 23599
rect 14945 23565 14979 23599
rect 15013 23565 15047 23599
rect 15081 23565 15115 23599
rect 15149 23565 15183 23599
rect 15217 23565 15251 23599
rect 15285 23565 15319 23599
rect 15353 23565 15387 23599
rect 15421 23565 15455 23599
rect 15489 23565 15523 23599
rect 15557 23565 15591 23599
rect 15625 23565 15659 23599
rect 15693 23565 15727 23599
rect 15761 23565 15795 23599
rect 15829 23565 15863 23599
rect 15897 23565 15931 23599
rect 15965 23565 15999 23599
rect 16033 23565 16067 23599
rect 16101 23565 16135 23599
rect 16169 23565 16203 23599
rect 16237 23565 16271 23599
rect 16305 23565 16339 23599
rect 16373 23565 16407 23599
rect 16441 23565 16475 23599
rect 16509 23565 16543 23599
rect 16577 23565 16611 23599
rect 16645 23565 16679 23599
rect 16713 23565 16747 23599
rect 16781 23565 16815 23599
rect 16849 23565 16883 23599
rect 16917 23565 16951 23599
rect 16985 23565 17019 23599
rect 17053 23565 17087 23599
rect 17121 23565 17155 23599
rect 17189 23565 17223 23599
rect 17257 23565 17291 23599
rect 17325 23565 17359 23599
rect 17393 23565 17427 23599
rect 17461 23565 17495 23599
rect 17529 23565 17563 23599
rect 17597 23565 17631 23599
rect 17665 23565 17699 23599
rect 17733 23565 17767 23599
rect 1089 23485 1123 23519
rect 1089 23417 1123 23451
rect 1089 23349 1123 23383
rect 17801 23458 17835 23492
rect 17801 23390 17835 23424
rect 1089 23281 1123 23315
rect 1089 23213 1123 23247
rect 1089 23145 1123 23179
rect 1089 23077 1123 23111
rect 1089 23009 1123 23043
rect 1089 22941 1123 22975
rect 1089 22873 1123 22907
rect 1089 22805 1123 22839
rect 1089 22737 1123 22771
rect 1089 22669 1123 22703
rect 1089 22601 1123 22635
rect 1089 22533 1123 22567
rect 1089 22465 1123 22499
rect 1089 22397 1123 22431
rect 1089 22329 1123 22363
rect 1089 22261 1123 22295
rect 1089 22193 1123 22227
rect 1089 22125 1123 22159
rect 1089 21976 1123 22010
rect 1157 21884 1191 21918
rect 1225 21884 1259 21918
rect 1293 21884 1327 21918
rect 1361 21884 1395 21918
rect 1429 21884 1463 21918
rect 1497 21884 1531 21918
rect 1565 21884 1599 21918
rect 1633 21884 1667 21918
rect 1701 21884 1735 21918
rect 1769 21884 1803 21918
rect 1837 21884 1871 21918
rect 1905 21884 1939 21918
rect 1973 21884 2007 21918
rect 2041 21884 2075 21918
rect 2109 21884 2143 21918
rect 2177 21884 2211 21918
rect 2245 21884 2279 21918
rect 17801 23322 17835 23356
rect 17801 23254 17835 23288
rect 17801 23186 17835 23220
rect 17801 23118 17835 23152
rect 17801 23050 17835 23084
rect 17801 22982 17835 23016
rect 17801 22914 17835 22948
rect 17801 22846 17835 22880
rect 17801 22778 17835 22812
rect 17801 22710 17835 22744
rect 17801 22642 17835 22676
rect 17801 22574 17835 22608
rect 17801 22506 17835 22540
rect 17801 22438 17835 22472
rect 17801 22370 17835 22404
rect 17801 22302 17835 22336
rect 17801 22234 17835 22268
rect 17801 22166 17835 22200
rect 17801 22098 17835 22132
rect 17801 22030 17835 22064
rect 17801 21962 17835 21996
rect 17801 21894 17835 21928
rect 17801 21826 17835 21860
rect 17801 21758 17835 21792
rect 17801 21690 17835 21724
rect 17801 21622 17835 21656
rect 17801 21554 17835 21588
rect 17801 21486 17835 21520
rect 17801 21418 17835 21452
rect 17801 21350 17835 21384
rect 17801 21282 17835 21316
rect 17801 21214 17835 21248
rect 17801 21146 17835 21180
rect 17801 21078 17835 21112
rect 17468 21010 17502 21044
rect 17536 21010 17570 21044
rect 17604 21010 17638 21044
rect 17672 21010 17706 21044
rect 12803 547 12837 581
rect 12871 547 12905 581
<< poly >>
rect 15463 23327 17063 23353
rect 15463 23201 17063 23243
rect 15463 23167 15506 23201
rect 15540 23167 15576 23201
rect 15610 23167 15646 23201
rect 15680 23167 15716 23201
rect 15750 23167 15786 23201
rect 15820 23167 15856 23201
rect 15890 23167 15926 23201
rect 15960 23167 15996 23201
rect 16030 23167 16066 23201
rect 16100 23167 16136 23201
rect 16170 23167 16206 23201
rect 16240 23167 16276 23201
rect 16310 23167 16346 23201
rect 16380 23167 16416 23201
rect 16450 23167 16486 23201
rect 16520 23167 16556 23201
rect 16590 23167 16626 23201
rect 16660 23167 16696 23201
rect 16730 23167 16766 23201
rect 16800 23167 16836 23201
rect 16870 23167 16906 23201
rect 16940 23167 16976 23201
rect 17010 23167 17063 23201
rect 15463 23125 17063 23167
rect 15463 22965 17063 23041
rect 15463 22836 17063 22881
rect 15463 22802 15506 22836
rect 15540 22802 15576 22836
rect 15610 22802 15646 22836
rect 15680 22802 15716 22836
rect 15750 22802 15786 22836
rect 15820 22802 15856 22836
rect 15890 22802 15926 22836
rect 15960 22802 15996 22836
rect 16030 22802 16066 22836
rect 16100 22802 16136 22836
rect 16170 22802 16206 22836
rect 16240 22802 16276 22836
rect 16310 22802 16346 22836
rect 16380 22802 16416 22836
rect 16450 22802 16486 22836
rect 16520 22802 16556 22836
rect 16590 22802 16626 22836
rect 16660 22802 16696 22836
rect 16730 22802 16766 22836
rect 16800 22802 16836 22836
rect 16870 22802 16906 22836
rect 16940 22802 16976 22836
rect 17010 22802 17063 22836
rect 15463 22763 17063 22802
rect 15463 22603 17063 22679
rect 15463 22443 17063 22519
rect 15463 22317 17063 22359
rect 15463 22283 15506 22317
rect 15540 22283 15576 22317
rect 15610 22283 15646 22317
rect 15680 22283 15716 22317
rect 15750 22283 15786 22317
rect 15820 22283 15856 22317
rect 15890 22283 15926 22317
rect 15960 22283 15996 22317
rect 16030 22283 16066 22317
rect 16100 22283 16136 22317
rect 16170 22283 16206 22317
rect 16240 22283 16276 22317
rect 16310 22283 16346 22317
rect 16380 22283 16416 22317
rect 16450 22283 16486 22317
rect 16520 22283 16556 22317
rect 16590 22283 16626 22317
rect 16660 22283 16696 22317
rect 16730 22283 16766 22317
rect 16800 22283 16836 22317
rect 16870 22283 16906 22317
rect 16940 22283 16976 22317
rect 17010 22283 17063 22317
rect 15463 22241 17063 22283
rect 15463 22081 17063 22157
rect 15463 21921 17063 21997
rect 15463 21795 17063 21837
rect 15463 21761 15506 21795
rect 15540 21761 15576 21795
rect 15610 21761 15646 21795
rect 15680 21761 15716 21795
rect 15750 21761 15786 21795
rect 15820 21761 15856 21795
rect 15890 21761 15926 21795
rect 15960 21761 15996 21795
rect 16030 21761 16066 21795
rect 16100 21761 16136 21795
rect 16170 21761 16206 21795
rect 16240 21761 16276 21795
rect 16310 21761 16346 21795
rect 16380 21761 16416 21795
rect 16450 21761 16486 21795
rect 16520 21761 16556 21795
rect 16590 21761 16626 21795
rect 16660 21761 16696 21795
rect 16730 21761 16766 21795
rect 16800 21761 16836 21795
rect 16870 21761 16906 21795
rect 16940 21761 16976 21795
rect 17010 21761 17063 21795
rect 15463 21719 17063 21761
rect 15463 21559 17063 21635
rect 15463 21433 17063 21475
rect 15463 21399 15506 21433
rect 15540 21399 15576 21433
rect 15610 21399 15646 21433
rect 15680 21399 15716 21433
rect 15750 21399 15786 21433
rect 15820 21399 15856 21433
rect 15890 21399 15926 21433
rect 15960 21399 15996 21433
rect 16030 21399 16066 21433
rect 16100 21399 16136 21433
rect 16170 21399 16206 21433
rect 16240 21399 16276 21433
rect 16310 21399 16346 21433
rect 16380 21399 16416 21433
rect 16450 21399 16486 21433
rect 16520 21399 16556 21433
rect 16590 21399 16626 21433
rect 16660 21399 16696 21433
rect 16730 21399 16766 21433
rect 16800 21399 16836 21433
rect 16870 21399 16906 21433
rect 16940 21399 16976 21433
rect 17010 21399 17063 21433
rect 15463 21357 17063 21399
rect 15463 21247 17063 21273
<< polycont >>
rect 15506 23167 15540 23201
rect 15576 23167 15610 23201
rect 15646 23167 15680 23201
rect 15716 23167 15750 23201
rect 15786 23167 15820 23201
rect 15856 23167 15890 23201
rect 15926 23167 15960 23201
rect 15996 23167 16030 23201
rect 16066 23167 16100 23201
rect 16136 23167 16170 23201
rect 16206 23167 16240 23201
rect 16276 23167 16310 23201
rect 16346 23167 16380 23201
rect 16416 23167 16450 23201
rect 16486 23167 16520 23201
rect 16556 23167 16590 23201
rect 16626 23167 16660 23201
rect 16696 23167 16730 23201
rect 16766 23167 16800 23201
rect 16836 23167 16870 23201
rect 16906 23167 16940 23201
rect 16976 23167 17010 23201
rect 15506 22802 15540 22836
rect 15576 22802 15610 22836
rect 15646 22802 15680 22836
rect 15716 22802 15750 22836
rect 15786 22802 15820 22836
rect 15856 22802 15890 22836
rect 15926 22802 15960 22836
rect 15996 22802 16030 22836
rect 16066 22802 16100 22836
rect 16136 22802 16170 22836
rect 16206 22802 16240 22836
rect 16276 22802 16310 22836
rect 16346 22802 16380 22836
rect 16416 22802 16450 22836
rect 16486 22802 16520 22836
rect 16556 22802 16590 22836
rect 16626 22802 16660 22836
rect 16696 22802 16730 22836
rect 16766 22802 16800 22836
rect 16836 22802 16870 22836
rect 16906 22802 16940 22836
rect 16976 22802 17010 22836
rect 15506 22283 15540 22317
rect 15576 22283 15610 22317
rect 15646 22283 15680 22317
rect 15716 22283 15750 22317
rect 15786 22283 15820 22317
rect 15856 22283 15890 22317
rect 15926 22283 15960 22317
rect 15996 22283 16030 22317
rect 16066 22283 16100 22317
rect 16136 22283 16170 22317
rect 16206 22283 16240 22317
rect 16276 22283 16310 22317
rect 16346 22283 16380 22317
rect 16416 22283 16450 22317
rect 16486 22283 16520 22317
rect 16556 22283 16590 22317
rect 16626 22283 16660 22317
rect 16696 22283 16730 22317
rect 16766 22283 16800 22317
rect 16836 22283 16870 22317
rect 16906 22283 16940 22317
rect 16976 22283 17010 22317
rect 15506 21761 15540 21795
rect 15576 21761 15610 21795
rect 15646 21761 15680 21795
rect 15716 21761 15750 21795
rect 15786 21761 15820 21795
rect 15856 21761 15890 21795
rect 15926 21761 15960 21795
rect 15996 21761 16030 21795
rect 16066 21761 16100 21795
rect 16136 21761 16170 21795
rect 16206 21761 16240 21795
rect 16276 21761 16310 21795
rect 16346 21761 16380 21795
rect 16416 21761 16450 21795
rect 16486 21761 16520 21795
rect 16556 21761 16590 21795
rect 16626 21761 16660 21795
rect 16696 21761 16730 21795
rect 16766 21761 16800 21795
rect 16836 21761 16870 21795
rect 16906 21761 16940 21795
rect 16976 21761 17010 21795
rect 15506 21399 15540 21433
rect 15576 21399 15610 21433
rect 15646 21399 15680 21433
rect 15716 21399 15750 21433
rect 15786 21399 15820 21433
rect 15856 21399 15890 21433
rect 15926 21399 15960 21433
rect 15996 21399 16030 21433
rect 16066 21399 16100 21433
rect 16136 21399 16170 21433
rect 16206 21399 16240 21433
rect 16276 21399 16310 21433
rect 16346 21399 16380 21433
rect 16416 21399 16450 21433
rect 16486 21399 16520 21433
rect 16556 21399 16590 21433
rect 16626 21399 16660 21433
rect 16696 21399 16730 21433
rect 16766 21399 16800 21433
rect 16836 21399 16870 21433
rect 16906 21399 16940 21433
rect 16976 21399 17010 21433
<< locali >>
rect 1089 24709 1209 24743
rect 1243 24709 1277 24743
rect 1311 24709 1345 24743
rect 1379 24709 1413 24743
rect 1447 24709 1481 24743
rect 1515 24709 1549 24743
rect 1583 24709 1617 24743
rect 1651 24709 1685 24743
rect 1719 24709 1753 24743
rect 1787 24709 1821 24743
rect 1855 24709 1889 24743
rect 1923 24709 1957 24743
rect 1991 24709 2025 24743
rect 2059 24709 2093 24743
rect 2127 24709 2161 24743
rect 2195 24709 2229 24743
rect 2263 24709 2297 24743
rect 2331 24709 2365 24743
rect 2399 24709 2433 24743
rect 2467 24709 2501 24743
rect 2535 24709 2569 24743
rect 2603 24709 2637 24743
rect 2671 24709 2705 24743
rect 2739 24709 2773 24743
rect 2807 24709 2841 24743
rect 2875 24709 2909 24743
rect 2943 24709 2977 24743
rect 3011 24709 3045 24743
rect 3079 24709 3113 24743
rect 3147 24709 3181 24743
rect 3215 24709 3249 24743
rect 3283 24709 3317 24743
rect 3351 24709 3385 24743
rect 3419 24709 3453 24743
rect 3487 24709 3521 24743
rect 3555 24709 3589 24743
rect 3623 24709 3657 24743
rect 3691 24709 3725 24743
rect 3759 24709 3793 24743
rect 3827 24709 3861 24743
rect 3895 24709 3929 24743
rect 3963 24709 3997 24743
rect 4031 24709 4065 24743
rect 4099 24709 4133 24743
rect 4167 24709 4201 24743
rect 4235 24709 4269 24743
rect 4303 24709 4337 24743
rect 4371 24709 4405 24743
rect 4439 24709 4473 24743
rect 4507 24709 4541 24743
rect 4575 24709 4609 24743
rect 4643 24709 4677 24743
rect 4711 24709 4745 24743
rect 4779 24709 4813 24743
rect 4847 24709 4881 24743
rect 4915 24709 4949 24743
rect 4983 24709 5017 24743
rect 5051 24709 5085 24743
rect 5119 24709 5153 24743
rect 5187 24709 5221 24743
rect 5255 24709 5289 24743
rect 5323 24709 5357 24743
rect 5391 24709 5425 24743
rect 5459 24709 5493 24743
rect 5527 24709 5561 24743
rect 5595 24709 5629 24743
rect 5663 24709 5697 24743
rect 5731 24709 5765 24743
rect 5799 24709 5833 24743
rect 5867 24709 5901 24743
rect 5935 24709 5969 24743
rect 6003 24709 6037 24743
rect 6071 24709 6105 24743
rect 6139 24709 6173 24743
rect 6207 24709 6241 24743
rect 6275 24709 6309 24743
rect 6343 24709 6377 24743
rect 6411 24709 6445 24743
rect 6479 24709 6513 24743
rect 6547 24709 6581 24743
rect 6615 24709 6649 24743
rect 6683 24709 6717 24743
rect 6751 24709 6785 24743
rect 6819 24709 6853 24743
rect 6887 24709 6921 24743
rect 6955 24709 6989 24743
rect 7023 24709 7057 24743
rect 7091 24709 7125 24743
rect 7159 24709 7193 24743
rect 7227 24709 7261 24743
rect 7295 24709 7329 24743
rect 7363 24709 7397 24743
rect 7431 24709 7465 24743
rect 7499 24709 7533 24743
rect 7567 24709 7601 24743
rect 7635 24709 7669 24743
rect 7703 24709 7737 24743
rect 7771 24709 7805 24743
rect 7839 24709 7873 24743
rect 7907 24709 7941 24743
rect 7975 24709 8009 24743
rect 8043 24709 8077 24743
rect 8111 24709 8145 24743
rect 8179 24709 8213 24743
rect 8247 24709 8281 24743
rect 8315 24709 8383 24743
rect 1089 24675 1123 24709
rect 1089 24607 1123 24641
rect 1089 24539 1123 24573
rect 1089 24471 1123 24505
rect 1089 24403 1123 24437
rect 1089 24335 1123 24369
rect 1089 24267 1123 24301
rect 1089 24199 1123 24233
rect 1089 24131 1123 24165
rect 1089 24063 1123 24097
rect 1089 23995 1123 24029
rect 1089 23927 1123 23961
rect 1089 23859 1123 23893
rect 1089 23791 1123 23825
rect 1089 23723 1123 23757
rect 1089 23655 1123 23689
rect 1089 23587 1123 23621
rect 8349 24619 8383 24709
rect 8349 24551 8383 24585
rect 8349 24483 8383 24517
rect 8349 24415 8383 24449
rect 8349 24347 8383 24381
rect 8349 24279 8383 24313
rect 8349 24211 8383 24245
rect 8349 24143 8383 24177
rect 8349 24075 8383 24109
rect 8349 24007 8383 24041
rect 8349 23939 8383 23973
rect 8349 23871 8383 23905
rect 8349 23803 8383 23837
rect 8349 23735 8383 23769
rect 8349 23667 8383 23701
rect 8349 23599 8383 23633
rect 8349 23565 8417 23599
rect 8451 23565 8485 23599
rect 8519 23565 8553 23599
rect 8587 23565 8621 23599
rect 8655 23565 8689 23599
rect 8723 23565 8757 23599
rect 8791 23565 8825 23599
rect 8859 23565 8893 23599
rect 8927 23565 8961 23599
rect 8995 23565 9029 23599
rect 9063 23565 9097 23599
rect 9131 23565 9165 23599
rect 9199 23565 9233 23599
rect 9267 23565 9301 23599
rect 9335 23565 9369 23599
rect 9403 23565 9437 23599
rect 9471 23565 9505 23599
rect 9539 23565 9573 23599
rect 9607 23565 9641 23599
rect 9675 23565 9709 23599
rect 9743 23565 9777 23599
rect 9811 23565 9845 23599
rect 9879 23565 9913 23599
rect 9947 23565 9981 23599
rect 10015 23565 10049 23599
rect 10083 23565 10117 23599
rect 10151 23565 10185 23599
rect 10219 23565 10253 23599
rect 10287 23565 10321 23599
rect 10355 23565 10389 23599
rect 10423 23565 10457 23599
rect 10491 23565 10525 23599
rect 10559 23565 10593 23599
rect 10627 23565 10661 23599
rect 10695 23565 10729 23599
rect 10763 23565 10797 23599
rect 10831 23565 10865 23599
rect 10899 23565 10933 23599
rect 10967 23565 11001 23599
rect 11035 23565 11069 23599
rect 11103 23565 11137 23599
rect 11171 23565 11205 23599
rect 11239 23565 11273 23599
rect 11307 23565 11341 23599
rect 11375 23565 11409 23599
rect 11443 23565 11477 23599
rect 11511 23565 11545 23599
rect 11579 23565 11613 23599
rect 11647 23565 11681 23599
rect 11715 23565 11749 23599
rect 11783 23565 11817 23599
rect 11851 23565 11885 23599
rect 11919 23565 11953 23599
rect 11987 23565 12021 23599
rect 12055 23565 12089 23599
rect 12123 23565 12157 23599
rect 12191 23565 12225 23599
rect 12259 23565 12293 23599
rect 12327 23565 12361 23599
rect 12395 23565 12429 23599
rect 12463 23565 12497 23599
rect 12531 23565 12565 23599
rect 12599 23565 12633 23599
rect 12667 23565 12701 23599
rect 12735 23565 12769 23599
rect 12803 23565 12837 23599
rect 12871 23565 12905 23599
rect 12939 23565 12973 23599
rect 13007 23565 13041 23599
rect 13075 23565 13109 23599
rect 13143 23565 13177 23599
rect 13211 23565 13245 23599
rect 13279 23565 13313 23599
rect 13347 23565 13381 23599
rect 13415 23565 13449 23599
rect 13483 23565 13517 23599
rect 13551 23565 13585 23599
rect 13619 23565 13653 23599
rect 13687 23565 13721 23599
rect 13755 23565 13789 23599
rect 13823 23565 13857 23599
rect 13891 23565 13925 23599
rect 13959 23565 13993 23599
rect 14027 23565 14061 23599
rect 14095 23565 14129 23599
rect 14163 23565 14197 23599
rect 14231 23565 14265 23599
rect 14299 23565 14333 23599
rect 14367 23565 14401 23599
rect 14435 23565 14469 23599
rect 14503 23565 14537 23599
rect 14571 23565 14605 23599
rect 14639 23565 14673 23599
rect 14707 23565 14741 23599
rect 14775 23565 14809 23599
rect 14843 23565 14877 23599
rect 14911 23565 14945 23599
rect 14979 23565 15013 23599
rect 15047 23565 15081 23599
rect 15115 23565 15149 23599
rect 15183 23565 15217 23599
rect 15251 23565 15285 23599
rect 15319 23565 15353 23599
rect 15387 23565 15421 23599
rect 15455 23565 15489 23599
rect 15523 23565 15557 23599
rect 15591 23565 15625 23599
rect 15659 23565 15693 23599
rect 15727 23565 15761 23599
rect 15795 23565 15829 23599
rect 15863 23565 15897 23599
rect 15931 23565 15965 23599
rect 15999 23565 16033 23599
rect 16067 23565 16101 23599
rect 16135 23565 16169 23599
rect 16203 23565 16237 23599
rect 16271 23565 16305 23599
rect 16339 23565 16373 23599
rect 16407 23565 16441 23599
rect 16475 23565 16509 23599
rect 16543 23565 16577 23599
rect 16611 23565 16645 23599
rect 16679 23565 16713 23599
rect 16747 23565 16781 23599
rect 16815 23565 16849 23599
rect 16883 23565 16917 23599
rect 16951 23565 16985 23599
rect 17019 23565 17053 23599
rect 17087 23565 17121 23599
rect 17155 23565 17189 23599
rect 17223 23565 17257 23599
rect 17291 23565 17325 23599
rect 17359 23565 17393 23599
rect 17427 23565 17461 23599
rect 17495 23565 17529 23599
rect 17563 23565 17597 23599
rect 17631 23565 17665 23599
rect 17699 23565 17733 23599
rect 17767 23565 17835 23599
rect 1089 23519 1123 23553
rect 1089 23451 1123 23485
rect 1089 23383 1123 23417
rect 17801 23492 17835 23565
rect 17801 23424 17835 23458
rect 1089 23315 1123 23349
rect 1089 23247 1123 23281
rect 15418 23315 15452 23349
rect 17801 23356 17835 23390
rect 15418 23265 15452 23277
rect 17074 23315 17180 23331
rect 17108 23281 17180 23315
rect 1089 23179 1123 23213
rect 17074 23209 17180 23281
rect 15490 23167 15506 23201
rect 15540 23167 15576 23201
rect 15610 23167 15646 23201
rect 15680 23167 15716 23201
rect 15750 23167 15786 23201
rect 15820 23167 15856 23201
rect 15890 23167 15926 23201
rect 15960 23167 15996 23201
rect 16030 23167 16066 23201
rect 16100 23167 16136 23201
rect 16170 23167 16206 23201
rect 16240 23167 16276 23201
rect 16310 23167 16346 23201
rect 16380 23167 16416 23201
rect 16450 23167 16486 23201
rect 16520 23167 16556 23201
rect 16590 23167 16626 23201
rect 16660 23167 16696 23201
rect 16730 23167 16766 23201
rect 16800 23167 16836 23201
rect 16870 23167 16906 23201
rect 16940 23167 16976 23201
rect 17010 23167 17026 23201
rect 17108 23175 17146 23209
rect 17220 23325 17254 23336
rect 17220 23302 17226 23325
rect 17254 23268 17260 23291
rect 17220 23252 17260 23268
rect 17220 23218 17226 23252
rect 17220 23217 17260 23218
rect 17254 23183 17260 23217
rect 17220 23179 17260 23183
rect 1089 23111 1123 23145
rect 1089 23043 1123 23077
rect 15418 23113 15452 23125
rect 1089 22975 1123 23009
rect 1089 22907 1123 22941
rect 15418 22953 15452 22965
rect 1089 22839 1123 22873
rect 1089 22771 1123 22805
rect 15490 22836 17026 23167
rect 17220 23145 17226 23179
rect 17220 23132 17260 23145
rect 17074 23113 17108 23129
rect 17108 23077 17146 23111
rect 17254 23106 17260 23132
rect 17074 23063 17108 23077
rect 17220 23072 17226 23098
rect 17220 23047 17260 23072
rect 17254 23033 17260 23047
rect 17220 22999 17226 23013
rect 17074 22953 17108 22969
rect 17220 22962 17260 22999
rect 17254 22960 17260 22962
rect 17108 22913 17146 22947
rect 17220 22926 17226 22928
rect 17074 22903 17108 22913
rect 15490 22802 15506 22836
rect 15540 22802 15576 22836
rect 15610 22802 15646 22836
rect 15680 22802 15716 22836
rect 15750 22802 15786 22836
rect 15820 22802 15856 22836
rect 15890 22802 15926 22836
rect 15960 22802 15996 22836
rect 16030 22802 16066 22836
rect 16100 22802 16136 22836
rect 16170 22802 16206 22836
rect 16240 22802 16276 22836
rect 16310 22802 16346 22836
rect 16380 22802 16416 22836
rect 16450 22802 16486 22836
rect 16520 22802 16556 22836
rect 16590 22802 16626 22836
rect 16660 22802 16696 22836
rect 16730 22802 16766 22836
rect 16800 22802 16836 22836
rect 16870 22802 16906 22836
rect 16940 22802 16976 22836
rect 17010 22802 17026 22836
rect 1089 22703 1123 22737
rect 15418 22751 15452 22763
rect 1089 22635 1123 22669
rect 1089 22567 1123 22601
rect 1089 22499 1123 22533
rect 15418 22591 15452 22603
rect 1089 22431 1123 22465
rect 1089 22363 1123 22397
rect 15418 22435 15452 22447
rect 15418 22363 15452 22397
rect 1089 22295 1123 22329
rect 15490 22317 17026 22802
rect 17220 22887 17260 22926
rect 17220 22877 17226 22887
rect 17254 22843 17260 22853
rect 17220 22814 17260 22843
rect 17220 22792 17226 22814
rect 17073 22758 17220 22767
rect 17254 22758 17260 22780
rect 17073 22751 17260 22758
rect 17073 22717 17074 22751
rect 17108 22741 17260 22751
rect 17108 22717 17226 22741
rect 17073 22712 17226 22717
rect 17073 22678 17120 22712
rect 17154 22707 17226 22712
rect 17154 22678 17220 22707
rect 17073 22673 17220 22678
rect 17254 22673 17260 22707
rect 17073 22668 17260 22673
rect 17073 22634 17226 22668
rect 17073 22622 17260 22634
rect 17073 22591 17120 22622
rect 17073 22557 17074 22591
rect 17108 22588 17120 22591
rect 17154 22588 17220 22622
rect 17254 22595 17260 22622
rect 17108 22561 17226 22588
rect 17108 22557 17260 22561
rect 17073 22537 17260 22557
rect 17073 22532 17220 22537
rect 17073 22498 17120 22532
rect 17154 22503 17220 22532
rect 17254 22522 17260 22537
rect 17154 22498 17226 22503
rect 17073 22488 17226 22498
rect 17073 22452 17260 22488
rect 17073 22442 17220 22452
rect 17254 22449 17260 22452
rect 17073 22431 17120 22442
rect 17073 22397 17074 22431
rect 17108 22408 17120 22431
rect 17154 22418 17220 22442
rect 17154 22415 17226 22418
rect 17154 22408 17260 22415
rect 17108 22397 17260 22408
rect 17073 22376 17260 22397
rect 17073 22367 17226 22376
rect 17073 22347 17220 22367
rect 15490 22283 15506 22317
rect 15540 22283 15576 22317
rect 15610 22283 15646 22317
rect 15680 22283 15716 22317
rect 15750 22283 15786 22317
rect 15820 22283 15856 22317
rect 15890 22283 15926 22317
rect 15960 22283 15996 22317
rect 16030 22283 16066 22317
rect 16100 22283 16136 22317
rect 16170 22283 16206 22317
rect 16240 22283 16276 22317
rect 16310 22283 16346 22317
rect 16380 22283 16416 22317
rect 16450 22283 16486 22317
rect 16520 22283 16556 22317
rect 16590 22283 16626 22317
rect 16660 22283 16696 22317
rect 16730 22283 16766 22317
rect 16800 22283 16836 22317
rect 16870 22283 16906 22317
rect 16940 22283 16976 22317
rect 17010 22283 17026 22317
rect 1089 22227 1123 22261
rect 1089 22159 1123 22193
rect 15418 22229 15452 22237
rect 1089 22010 1123 22125
rect 15418 22027 15452 22035
rect 1089 21918 1123 21976
rect 1089 21884 1157 21918
rect 1191 21884 1225 21918
rect 1259 21884 1293 21918
rect 1327 21884 1361 21918
rect 1395 21884 1429 21918
rect 1463 21884 1497 21918
rect 1531 21884 1565 21918
rect 1599 21884 1633 21918
rect 1667 21884 1701 21918
rect 1735 21884 1769 21918
rect 1803 21884 1837 21918
rect 1871 21884 1905 21918
rect 1939 21884 1973 21918
rect 2007 21884 2041 21918
rect 2075 21884 2109 21918
rect 2143 21884 2177 21918
rect 2211 21884 2245 21918
rect 2279 21884 2317 21918
rect 15418 21867 15452 21875
rect 15490 21795 17026 22283
rect 17254 22333 17260 22342
rect 17220 22303 17260 22333
rect 17220 22282 17226 22303
rect 17254 22248 17260 22269
rect 17074 22229 17108 22245
rect 17220 22230 17260 22248
rect 17108 22195 17146 22229
rect 17220 22197 17226 22230
rect 17074 22179 17108 22195
rect 17254 22163 17260 22196
rect 17220 22157 17260 22163
rect 17074 22069 17108 22091
rect 17220 22123 17226 22157
rect 17220 22112 17260 22123
rect 17254 22084 17260 22112
rect 17220 22050 17226 22078
rect 17220 22027 17260 22050
rect 17254 22011 17260 22027
rect 17220 21977 17226 21993
rect 17074 21909 17108 21931
rect 17220 21942 17260 21977
rect 17254 21937 17260 21942
rect 17220 21903 17226 21908
rect 17220 21863 17260 21903
rect 15490 21761 15506 21795
rect 15540 21761 15576 21795
rect 15610 21761 15646 21795
rect 15680 21761 15716 21795
rect 15750 21761 15786 21795
rect 15820 21761 15856 21795
rect 15890 21761 15926 21795
rect 15960 21761 15996 21795
rect 16030 21761 16066 21795
rect 16100 21761 16136 21795
rect 16170 21761 16181 21795
rect 16240 21761 16254 21795
rect 16310 21761 16327 21795
rect 16380 21761 16400 21795
rect 16450 21761 16473 21795
rect 16520 21761 16546 21795
rect 16590 21761 16619 21795
rect 16660 21761 16692 21795
rect 16730 21761 16764 21795
rect 16800 21761 16836 21795
rect 16870 21761 16906 21795
rect 16942 21761 16976 21795
rect 17014 21761 17026 21795
rect 15418 21707 15452 21720
rect 15418 21547 15452 21550
rect 15418 21512 15452 21513
rect 15490 21440 17026 21761
rect 17220 21857 17226 21863
rect 17254 21823 17260 21829
rect 17220 21789 17260 21823
rect 17220 21772 17226 21789
rect 17254 21738 17260 21755
rect 15490 21433 16179 21440
rect 16213 21433 16252 21440
rect 16286 21433 16325 21440
rect 16359 21433 16398 21440
rect 16432 21433 16471 21440
rect 16505 21433 16544 21440
rect 16578 21433 16617 21440
rect 16651 21433 16690 21440
rect 16724 21433 16763 21440
rect 16797 21433 16836 21440
rect 16870 21433 16908 21440
rect 16942 21433 16980 21440
rect 15490 21399 15506 21433
rect 15540 21399 15576 21433
rect 15610 21399 15646 21433
rect 15680 21399 15716 21433
rect 15750 21399 15786 21433
rect 15820 21399 15856 21433
rect 15890 21399 15926 21433
rect 15960 21399 15996 21433
rect 16030 21399 16066 21433
rect 16100 21399 16136 21433
rect 16170 21406 16179 21433
rect 16240 21406 16252 21433
rect 16310 21406 16325 21433
rect 16380 21406 16398 21433
rect 16450 21406 16471 21433
rect 16520 21406 16544 21433
rect 16590 21406 16617 21433
rect 16660 21406 16690 21433
rect 16730 21406 16763 21433
rect 16170 21399 16206 21406
rect 16240 21399 16276 21406
rect 16310 21399 16346 21406
rect 16380 21399 16416 21406
rect 16450 21399 16486 21406
rect 16520 21399 16556 21406
rect 16590 21399 16626 21406
rect 16660 21399 16696 21406
rect 16730 21399 16766 21406
rect 16800 21399 16836 21433
rect 16870 21399 16906 21433
rect 16942 21406 16976 21433
rect 17014 21406 17026 21440
rect 16940 21399 16976 21406
rect 17010 21399 17026 21406
rect 17066 21716 17186 21725
rect 17066 21682 17073 21716
rect 17107 21707 17145 21716
rect 17108 21682 17145 21707
rect 17179 21682 17186 21716
rect 17066 21673 17074 21682
rect 17108 21673 17186 21682
rect 17066 21638 17186 21673
rect 17066 21604 17073 21638
rect 17107 21604 17145 21638
rect 17179 21604 17186 21638
rect 17066 21560 17186 21604
rect 17066 21526 17073 21560
rect 17107 21547 17145 21560
rect 17108 21526 17145 21547
rect 17179 21526 17186 21560
rect 17066 21513 17074 21526
rect 17108 21513 17186 21526
rect 17066 21481 17186 21513
rect 17066 21447 17073 21481
rect 17107 21447 17145 21481
rect 17179 21447 17186 21481
rect 17066 21402 17186 21447
rect 15418 21305 15452 21311
rect 17066 21368 17073 21402
rect 17107 21368 17145 21402
rect 17179 21368 17186 21402
rect 17066 21345 17186 21368
rect 17066 21323 17074 21345
rect 17108 21323 17186 21345
rect 17066 21289 17073 21323
rect 17108 21311 17145 21323
rect 17107 21289 17145 21311
rect 17179 21289 17186 21323
rect 17066 21280 17186 21289
rect 17220 21715 17260 21738
rect 17220 21687 17226 21715
rect 17254 21653 17260 21681
rect 17220 21641 17260 21653
rect 17220 21607 17226 21641
rect 17220 21602 17260 21607
rect 17254 21568 17260 21602
rect 17220 21567 17260 21568
rect 17220 21533 17226 21567
rect 17220 21517 17260 21533
rect 17254 21493 17260 21517
rect 17220 21459 17226 21483
rect 17220 21432 17260 21459
rect 17254 21419 17260 21432
rect 17220 21385 17226 21398
rect 17220 21347 17260 21385
rect 17254 21345 17260 21347
rect 17220 21311 17226 21313
rect 17220 21279 17260 21311
rect 17226 21271 17260 21279
rect 17801 23288 17835 23322
rect 17801 23220 17835 23254
rect 17801 23152 17835 23186
rect 17801 23084 17835 23118
rect 17801 23016 17835 23050
rect 17801 22948 17835 22982
rect 17801 22880 17835 22914
rect 17801 22812 17835 22846
rect 17801 22744 17835 22778
rect 17801 22676 17835 22710
rect 17801 22608 17835 22642
rect 17801 22540 17835 22574
rect 17801 22472 17835 22506
rect 17801 22404 17835 22438
rect 17801 22336 17835 22370
rect 17801 22268 17835 22302
rect 17801 22200 17835 22234
rect 17801 22132 17835 22166
rect 17801 22064 17835 22098
rect 17801 21996 17835 22030
rect 17801 21928 17835 21962
rect 17801 21860 17835 21894
rect 17801 21792 17835 21826
rect 17801 21724 17835 21758
rect 17801 21656 17835 21690
rect 17801 21588 17835 21622
rect 17801 21520 17835 21554
rect 17801 21452 17835 21486
rect 17801 21384 17835 21418
rect 17801 21316 17835 21350
rect 17801 21248 17835 21282
rect 17801 21180 17835 21214
rect 17801 21112 17835 21146
rect 17801 21044 17835 21078
rect 17434 21010 17468 21044
rect 17502 21010 17536 21044
rect 17570 21010 17604 21044
rect 17638 21010 17672 21044
rect 17706 21010 17835 21044
rect 22920 9800 22958 9834
rect 22868 9559 22902 9597
rect 12803 581 12905 625
rect 12837 547 12871 581
rect 12803 523 12905 547
<< viali >>
rect 15418 23349 15452 23383
rect 15418 23281 15452 23311
rect 15418 23277 15452 23281
rect 17074 23175 17108 23209
rect 17146 23175 17180 23209
rect 17226 23302 17260 23325
rect 17226 23291 17254 23302
rect 17254 23291 17260 23302
rect 17226 23218 17260 23252
rect 15418 23125 15452 23159
rect 15418 23079 15452 23087
rect 15418 23053 15452 23079
rect 15418 22965 15452 22999
rect 15418 22919 15452 22927
rect 15418 22893 15452 22919
rect 17226 23145 17260 23179
rect 17074 23079 17108 23111
rect 17074 23077 17108 23079
rect 17146 23077 17180 23111
rect 17226 23098 17254 23106
rect 17254 23098 17260 23106
rect 17226 23072 17260 23098
rect 17226 23013 17254 23033
rect 17254 23013 17260 23033
rect 17226 22999 17260 23013
rect 17074 22919 17108 22947
rect 17074 22913 17108 22919
rect 17146 22913 17180 22947
rect 17226 22928 17254 22960
rect 17254 22928 17260 22960
rect 17226 22926 17260 22928
rect 15418 22763 15452 22797
rect 15418 22717 15452 22725
rect 15418 22691 15452 22717
rect 15418 22603 15452 22637
rect 15418 22557 15452 22565
rect 15418 22531 15452 22557
rect 15418 22431 15452 22435
rect 15418 22401 15452 22431
rect 15418 22329 15452 22363
rect 17226 22877 17260 22887
rect 17226 22853 17254 22877
rect 17254 22853 17260 22877
rect 17226 22792 17260 22814
rect 17226 22780 17254 22792
rect 17254 22780 17260 22792
rect 17120 22678 17154 22712
rect 17226 22707 17260 22741
rect 17226 22634 17260 22668
rect 17120 22588 17154 22622
rect 17226 22588 17254 22595
rect 17254 22588 17260 22595
rect 17226 22561 17260 22588
rect 17120 22498 17154 22532
rect 17226 22503 17254 22522
rect 17254 22503 17260 22522
rect 17226 22488 17260 22503
rect 17120 22408 17154 22442
rect 17226 22418 17254 22449
rect 17254 22418 17260 22449
rect 17226 22415 17260 22418
rect 17226 22367 17260 22376
rect 15418 22237 15452 22271
rect 15418 22195 15452 22199
rect 15418 22165 15452 22195
rect 15418 22069 15452 22099
rect 15418 22065 15452 22069
rect 15418 21993 15452 22027
rect 15418 21909 15452 21939
rect 15418 21905 15452 21909
rect 15418 21833 15452 21867
rect 17226 22342 17254 22367
rect 17254 22342 17260 22367
rect 17226 22282 17260 22303
rect 17226 22269 17254 22282
rect 17254 22269 17260 22282
rect 17074 22195 17108 22229
rect 17146 22195 17180 22229
rect 17226 22197 17260 22230
rect 17226 22196 17254 22197
rect 17254 22196 17260 22197
rect 17074 22091 17108 22125
rect 17074 22035 17108 22053
rect 17074 22019 17108 22035
rect 17226 22123 17260 22157
rect 17226 22078 17254 22084
rect 17254 22078 17260 22084
rect 17226 22050 17260 22078
rect 17226 21993 17254 22011
rect 17254 21993 17260 22011
rect 17226 21977 17260 21993
rect 17074 21931 17108 21965
rect 17074 21875 17108 21893
rect 17074 21859 17108 21875
rect 17226 21908 17254 21937
rect 17254 21908 17260 21937
rect 17226 21903 17260 21908
rect 16181 21761 16206 21795
rect 16206 21761 16215 21795
rect 16254 21761 16276 21795
rect 16276 21761 16288 21795
rect 16327 21761 16346 21795
rect 16346 21761 16361 21795
rect 16400 21761 16416 21795
rect 16416 21761 16434 21795
rect 16473 21761 16486 21795
rect 16486 21761 16507 21795
rect 16546 21761 16556 21795
rect 16556 21761 16580 21795
rect 16619 21761 16626 21795
rect 16626 21761 16653 21795
rect 16692 21761 16696 21795
rect 16696 21761 16726 21795
rect 16764 21761 16766 21795
rect 16766 21761 16798 21795
rect 16836 21761 16870 21795
rect 16908 21761 16940 21795
rect 16940 21761 16942 21795
rect 16980 21761 17010 21795
rect 17010 21761 17014 21795
rect 15418 21720 15452 21754
rect 15418 21673 15452 21682
rect 15418 21648 15452 21673
rect 15418 21550 15452 21584
rect 15418 21478 15452 21512
rect 17226 21857 17260 21863
rect 17226 21829 17254 21857
rect 17254 21829 17260 21857
rect 17226 21772 17260 21789
rect 17226 21755 17254 21772
rect 17254 21755 17260 21772
rect 16179 21433 16213 21440
rect 16252 21433 16286 21440
rect 16325 21433 16359 21440
rect 16398 21433 16432 21440
rect 16471 21433 16505 21440
rect 16544 21433 16578 21440
rect 16617 21433 16651 21440
rect 16690 21433 16724 21440
rect 16763 21433 16797 21440
rect 16836 21433 16870 21440
rect 16908 21433 16942 21440
rect 16980 21433 17014 21440
rect 16179 21406 16206 21433
rect 16206 21406 16213 21433
rect 16252 21406 16276 21433
rect 16276 21406 16286 21433
rect 16325 21406 16346 21433
rect 16346 21406 16359 21433
rect 16398 21406 16416 21433
rect 16416 21406 16432 21433
rect 16471 21406 16486 21433
rect 16486 21406 16505 21433
rect 16544 21406 16556 21433
rect 16556 21406 16578 21433
rect 16617 21406 16626 21433
rect 16626 21406 16651 21433
rect 16690 21406 16696 21433
rect 16696 21406 16724 21433
rect 16763 21406 16766 21433
rect 16766 21406 16797 21433
rect 16836 21406 16870 21433
rect 16908 21406 16940 21433
rect 16940 21406 16942 21433
rect 16980 21406 17010 21433
rect 17010 21406 17014 21433
rect 17073 21707 17107 21716
rect 17073 21682 17074 21707
rect 17074 21682 17107 21707
rect 17145 21682 17179 21716
rect 17073 21604 17107 21638
rect 17145 21604 17179 21638
rect 17073 21547 17107 21560
rect 17073 21526 17074 21547
rect 17074 21526 17107 21547
rect 17145 21526 17179 21560
rect 17073 21447 17107 21481
rect 17145 21447 17179 21481
rect 15418 21345 15452 21377
rect 15418 21343 15452 21345
rect 15418 21271 15452 21305
rect 17073 21368 17107 21402
rect 17145 21368 17179 21402
rect 17073 21311 17074 21323
rect 17074 21311 17107 21323
rect 17073 21289 17107 21311
rect 17145 21289 17179 21323
rect 17226 21687 17260 21715
rect 17226 21681 17254 21687
rect 17254 21681 17260 21687
rect 17226 21607 17260 21641
rect 17226 21533 17260 21567
rect 17226 21483 17254 21493
rect 17254 21483 17260 21493
rect 17226 21459 17260 21483
rect 17226 21398 17254 21419
rect 17254 21398 17260 21419
rect 17226 21385 17260 21398
rect 17226 21313 17254 21345
rect 17254 21313 17260 21345
rect 17226 21311 17260 21313
rect 17226 21237 17260 21271
rect 22886 9800 22920 9834
rect 22958 9800 22992 9834
rect 24964 9756 25070 9862
rect 22868 9597 22902 9631
rect 22868 9525 22902 9559
rect 24955 9524 25061 9630
<< metal1 >>
rect 15412 23383 15653 23395
rect 15412 23349 15418 23383
rect 15452 23366 15653 23383
tri 15653 23366 15682 23395 sw
rect 15452 23349 15682 23366
rect 15412 23311 15682 23349
rect 15412 23277 15418 23311
rect 15452 23277 15682 23311
rect 15412 23265 15682 23277
tri 15594 23252 15607 23265 ne
rect 15607 23252 15682 23265
tri 15607 23223 15636 23252 ne
rect 15412 23166 15571 23171
tri 15571 23166 15576 23171 sw
rect 15412 23159 15576 23166
rect 15412 23125 15418 23159
rect 15452 23145 15576 23159
tri 15576 23145 15597 23166 sw
rect 15452 23134 15597 23145
tri 15597 23134 15608 23145 sw
rect 15452 23125 15608 23134
rect 15412 23087 15608 23125
rect 15412 23053 15418 23087
rect 15452 23053 15608 23087
rect 15412 23041 15608 23053
tri 15524 23033 15532 23041 ne
rect 15532 23033 15608 23041
tri 15532 23011 15554 23033 ne
rect 15554 23011 15608 23033
rect 15412 22999 15458 23011
tri 15554 23003 15562 23011 ne
rect 15412 22965 15418 22999
rect 15452 22965 15458 22999
rect 15412 22927 15458 22965
rect 15412 22893 15418 22927
rect 15452 22893 15458 22927
rect 15412 22797 15458 22893
rect 15412 22763 15418 22797
rect 15452 22763 15458 22797
rect 15412 22725 15458 22763
rect 15412 22691 15418 22725
rect 15452 22691 15458 22725
rect 15412 22679 15458 22691
tri 15559 22668 15562 22671 se
rect 15562 22668 15608 23011
tri 15540 22649 15559 22668 se
rect 15559 22649 15608 22668
rect 15412 22637 15608 22649
rect 15412 22603 15418 22637
rect 15452 22603 15608 22637
rect 15412 22565 15608 22603
rect 15412 22531 15418 22565
rect 15452 22535 15608 22565
rect 15452 22532 15605 22535
tri 15605 22532 15608 22535 nw
rect 15452 22531 15592 22532
rect 15412 22519 15592 22531
tri 15592 22519 15605 22532 nw
tri 15616 22449 15636 22469 se
rect 15636 22449 15682 23252
rect 17220 23325 17266 23337
rect 17220 23291 17226 23325
rect 17260 23291 17266 23325
rect 17220 23252 17266 23291
rect 17220 23218 17226 23252
rect 17260 23218 17266 23252
rect 17062 23166 17068 23218
rect 17120 23166 17132 23218
rect 17184 23166 17192 23218
rect 17220 23179 17266 23218
rect 17220 23145 17226 23179
rect 17260 23145 17266 23179
rect 17062 23068 17068 23120
rect 17120 23068 17132 23120
rect 17184 23068 17192 23120
rect 17220 23106 17266 23145
rect 17220 23072 17226 23106
rect 17260 23072 17266 23106
rect 17220 23033 17266 23072
rect 17220 22999 17226 23033
rect 17260 22999 17266 23033
rect 17220 22960 17266 22999
rect 16252 22880 16258 22932
rect 16310 22880 16348 22932
rect 16400 22880 16438 22932
rect 16490 22880 16527 22932
rect 16579 22913 16659 22932
tri 16659 22913 16678 22932 sw
rect 16579 22904 16678 22913
tri 16678 22904 16687 22913 sw
rect 17062 22904 17068 22956
rect 17120 22904 17132 22956
rect 17184 22904 17192 22956
rect 17220 22926 17226 22960
rect 17260 22926 17266 22960
rect 16579 22887 16687 22904
tri 16687 22887 16704 22904 sw
rect 17220 22887 17266 22926
rect 16579 22880 16704 22887
rect 16252 22853 16704 22880
tri 16704 22853 16738 22887 sw
tri 17215 22853 17220 22858 se
rect 17220 22853 17226 22887
rect 17260 22853 17266 22887
rect 16252 22840 16738 22853
rect 16252 22788 16258 22840
rect 16310 22788 16348 22840
rect 16400 22788 16438 22840
rect 16490 22788 16527 22840
rect 16579 22814 16738 22840
tri 16738 22814 16777 22853 sw
tri 17176 22814 17215 22853 se
rect 17215 22814 17266 22853
rect 16579 22788 16777 22814
rect 16252 22780 16777 22788
tri 16777 22780 16811 22814 sw
tri 17142 22780 17176 22814 se
rect 17176 22780 17226 22814
rect 17260 22780 17266 22814
rect 16252 22748 16811 22780
rect 16252 22696 16258 22748
rect 16310 22696 16348 22748
rect 16400 22696 16438 22748
rect 16490 22696 16527 22748
rect 16579 22741 16811 22748
tri 16811 22741 16850 22780 sw
tri 17103 22741 17142 22780 se
rect 17142 22741 17266 22780
rect 16579 22724 16850 22741
tri 16850 22724 16867 22741 sw
tri 17086 22724 17103 22741 se
rect 17103 22724 17226 22741
rect 16579 22712 17226 22724
rect 16579 22696 17120 22712
rect 16252 22678 17120 22696
rect 17154 22707 17226 22712
rect 17260 22707 17266 22741
rect 17154 22678 17266 22707
rect 16252 22668 17266 22678
rect 16252 22656 17226 22668
rect 16252 22604 16258 22656
rect 16310 22604 16348 22656
rect 16400 22604 16438 22656
rect 16490 22604 16527 22656
rect 16579 22634 17226 22656
rect 17260 22634 17266 22668
rect 16579 22622 17266 22634
rect 16579 22604 17120 22622
tri 16523 22588 16539 22604 ne
rect 16539 22588 17120 22604
rect 17154 22595 17266 22622
rect 17154 22588 17226 22595
tri 16539 22561 16566 22588 ne
rect 16566 22561 17226 22588
rect 17260 22561 17266 22595
tri 16566 22532 16595 22561 ne
rect 16595 22532 17266 22561
tri 16595 22498 16629 22532 ne
rect 16629 22498 17120 22532
rect 17154 22522 17266 22532
rect 17154 22498 17226 22522
tri 16629 22488 16639 22498 ne
rect 16639 22488 17226 22498
rect 17260 22488 17266 22522
tri 16639 22449 16678 22488 ne
rect 16678 22449 17266 22488
tri 15614 22447 15616 22449 se
rect 15616 22447 15682 22449
rect 15412 22435 15682 22447
tri 16678 22442 16685 22449 ne
rect 16685 22442 17226 22449
rect 15412 22401 15418 22435
rect 15452 22401 15682 22435
tri 16685 22408 16719 22442 ne
rect 16719 22408 17120 22442
rect 17154 22415 17226 22442
rect 17260 22415 17266 22449
rect 17154 22408 17266 22415
rect 15412 22363 15682 22401
tri 16719 22396 16731 22408 ne
rect 16731 22396 17266 22408
tri 17086 22376 17106 22396 ne
rect 17106 22376 17266 22396
rect 15412 22329 15418 22363
rect 15452 22335 15682 22363
tri 17106 22342 17140 22376 ne
rect 17140 22342 17226 22376
rect 17260 22342 17266 22376
rect 15452 22329 15664 22335
rect 15412 22317 15664 22329
tri 15664 22317 15682 22335 nw
tri 17140 22327 17155 22342 ne
rect 17155 22327 17266 22342
tri 16521 22317 16531 22327 se
rect 16531 22317 16947 22327
tri 16947 22317 16957 22327 sw
tri 17155 22317 17165 22327 ne
rect 17165 22317 17266 22327
tri 16507 22303 16521 22317 se
rect 16521 22303 16957 22317
tri 16957 22303 16971 22317 sw
tri 17165 22303 17179 22317 ne
rect 17179 22303 17266 22317
tri 16505 22301 16507 22303 se
rect 16507 22301 16971 22303
tri 16971 22301 16973 22303 sw
tri 17179 22301 17181 22303 ne
rect 17181 22301 17226 22303
tri 16487 22283 16505 22301 se
rect 16505 22283 16973 22301
tri 16973 22283 16991 22301 sw
tri 17181 22283 17199 22301 ne
rect 17199 22283 17226 22301
rect 15412 22271 15653 22283
rect 15412 22237 15418 22271
rect 15452 22269 15653 22271
tri 15653 22269 15667 22283 sw
tri 16473 22269 16487 22283 se
rect 16487 22281 16991 22283
rect 16487 22269 16539 22281
tri 16539 22269 16551 22281 nw
tri 16927 22269 16939 22281 ne
rect 16939 22269 16991 22281
tri 16991 22269 17005 22283 sw
tri 17199 22269 17213 22283 ne
rect 17213 22269 17226 22283
rect 17260 22269 17266 22303
rect 15452 22254 15667 22269
tri 15667 22254 15682 22269 sw
tri 16465 22261 16473 22269 se
rect 16473 22261 16531 22269
tri 16531 22261 16539 22269 nw
tri 16939 22261 16947 22269 ne
rect 16947 22261 17005 22269
rect 15452 22237 15682 22254
rect 15412 22199 15682 22237
rect 15412 22165 15418 22199
rect 15452 22165 15682 22199
rect 15412 22153 15682 22165
tri 15594 22125 15622 22153 ne
rect 15622 22125 15682 22153
tri 15622 22111 15636 22125 ne
rect 15412 22099 15571 22111
rect 15412 22065 15418 22099
rect 15452 22091 15571 22099
tri 15571 22091 15591 22111 sw
rect 15452 22084 15591 22091
tri 15591 22084 15598 22091 sw
rect 15452 22074 15598 22084
tri 15598 22074 15608 22084 sw
rect 15452 22065 15608 22074
rect 15412 22027 15608 22065
rect 15412 21993 15418 22027
rect 15452 21993 15608 22027
rect 15412 21981 15608 21993
tri 15524 21977 15528 21981 ne
rect 15528 21977 15608 21981
tri 15528 21965 15540 21977 ne
rect 15540 21965 15608 21977
tri 15540 21951 15554 21965 ne
rect 15554 21951 15608 21965
rect 15412 21939 15458 21951
tri 15554 21943 15562 21951 ne
rect 15412 21905 15418 21939
rect 15452 21905 15458 21939
rect 15412 21867 15458 21905
rect 15412 21833 15418 21867
rect 15452 21833 15458 21867
rect 14624 21809 14759 21815
rect 14624 21757 14641 21809
rect 14693 21757 14707 21809
rect 14624 21726 14759 21757
rect 14624 21674 14641 21726
rect 14693 21674 14707 21726
rect 14624 21643 14759 21674
rect 14624 21591 14641 21643
rect 14693 21591 14707 21643
rect 15412 21754 15458 21833
rect 15412 21720 15418 21754
rect 15452 21720 15458 21754
rect 15412 21682 15458 21720
rect 15412 21648 15418 21682
rect 15452 21648 15458 21682
rect 15412 21636 15458 21648
tri 15555 21604 15562 21611 se
rect 15562 21604 15608 21951
tri 15547 21596 15555 21604 se
rect 15555 21596 15608 21604
rect 14624 21560 14759 21591
rect 14624 21508 14641 21560
rect 14693 21508 14707 21560
rect 14624 21377 14759 21508
rect 15412 21584 15608 21596
rect 15412 21550 15418 21584
rect 15452 21550 15608 21584
rect 15412 21512 15608 21550
rect 15412 21478 15418 21512
rect 15452 21478 15608 21512
rect 15412 21475 15608 21478
rect 15412 21466 15599 21475
tri 15599 21466 15608 21475 nw
tri 15631 21406 15636 21411 se
rect 15636 21406 15682 22125
tri 16439 22235 16465 22261 se
rect 16465 22235 16505 22261
tri 16505 22235 16531 22261 nw
tri 16947 22235 16973 22261 ne
rect 16973 22235 17005 22261
tri 17005 22235 17039 22269 sw
tri 17213 22262 17220 22269 ne
rect 16439 22230 16500 22235
tri 16500 22230 16505 22235 nw
tri 16973 22230 16978 22235 ne
rect 16978 22230 17192 22235
rect 16439 22229 16499 22230
tri 16499 22229 16500 22230 nw
tri 16978 22229 16979 22230 ne
rect 16979 22229 17192 22230
tri 16421 21911 16439 21929 se
rect 16439 21911 16485 22229
tri 16485 22215 16499 22229 nw
tri 16979 22215 16993 22229 ne
rect 16993 22215 17074 22229
tri 16993 22195 17013 22215 ne
rect 17013 22195 17074 22215
rect 17108 22195 17146 22229
rect 17180 22195 17192 22229
tri 17013 22189 17019 22195 ne
rect 17019 22189 17192 22195
rect 17220 22230 17266 22269
rect 17220 22196 17226 22230
rect 17260 22196 17266 22230
rect 17220 22157 17266 22196
tri 17057 22125 17068 22136 se
rect 17068 22125 17114 22137
tri 17054 22122 17057 22125 se
rect 17057 22122 17074 22125
tri 16789 22091 16820 22122 se
rect 16820 22091 17074 22122
rect 17108 22091 17114 22125
tri 16782 22084 16789 22091 se
rect 16789 22084 17114 22091
tri 16751 22053 16782 22084 se
rect 16782 22070 17114 22084
rect 16782 22053 16825 22070
tri 16825 22053 16842 22070 nw
tri 17032 22053 17049 22070 ne
rect 17049 22053 17114 22070
tri 16746 22048 16751 22053 se
rect 16751 22048 16820 22053
tri 16820 22048 16825 22053 nw
tri 17049 22048 17054 22053 ne
rect 17054 22048 17074 22053
tri 16717 22019 16746 22048 se
rect 16746 22019 16791 22048
tri 16791 22019 16820 22048 nw
tri 17054 22034 17068 22048 ne
rect 17068 22019 17074 22048
rect 17108 22019 17114 22053
tri 16709 22011 16717 22019 se
rect 16717 22011 16787 22019
tri 16787 22015 16791 22019 nw
tri 16705 22007 16709 22011 se
rect 16709 22007 16787 22011
rect 17068 22007 17114 22019
rect 17220 22123 17226 22157
rect 17260 22123 17266 22157
rect 17220 22084 17266 22123
rect 17220 22050 17226 22084
rect 17260 22050 17266 22084
rect 17220 22011 17266 22050
tri 16675 21977 16705 22007 se
rect 16705 21977 16787 22007
rect 17220 21977 17226 22011
rect 17260 21977 17266 22011
tri 16663 21965 16675 21977 se
rect 16675 21965 16787 21977
tri 17056 21965 17068 21977 se
rect 17068 21965 17114 21977
tri 16661 21963 16663 21965 se
rect 16663 21963 16787 21965
tri 17054 21963 17056 21965 se
rect 17056 21963 17074 21965
tri 16485 21911 16503 21929 sw
rect 16659 21911 16665 21963
rect 16717 21911 16729 21963
rect 16781 21911 16787 21963
rect 16849 21911 16855 21963
rect 16907 21911 16919 21963
rect 16971 21931 17074 21963
rect 17108 21931 17114 21965
rect 16971 21911 17114 21931
tri 16413 21903 16421 21911 se
rect 16421 21903 16503 21911
tri 16503 21903 16511 21911 sw
tri 17023 21903 17031 21911 ne
rect 17031 21903 17114 21911
tri 16405 21895 16413 21903 se
rect 16413 21895 16511 21903
tri 16511 21895 16519 21903 sw
tri 17031 21895 17039 21903 ne
rect 17039 21895 17114 21903
rect 16404 21843 16410 21895
rect 16462 21843 16476 21895
rect 16528 21843 16534 21895
tri 17039 21893 17041 21895 ne
rect 17041 21893 17114 21895
tri 17041 21866 17068 21893 ne
rect 17068 21859 17074 21893
rect 17108 21859 17114 21893
rect 17068 21847 17114 21859
rect 17220 21937 17266 21977
rect 17220 21903 17226 21937
rect 17260 21903 17266 21937
rect 17220 21863 17266 21903
rect 17220 21829 17226 21863
rect 17260 21829 17266 21863
rect 16169 21795 17026 21801
rect 16169 21761 16181 21795
rect 16215 21761 16254 21795
rect 16288 21761 16327 21795
rect 16361 21761 16400 21795
rect 16434 21761 16473 21795
rect 16507 21761 16546 21795
rect 16580 21761 16619 21795
rect 16653 21761 16692 21795
rect 16726 21761 16764 21795
rect 16798 21761 16836 21795
rect 16870 21761 16908 21795
rect 16942 21761 16980 21795
rect 17014 21761 17026 21795
rect 16169 21755 17026 21761
rect 17220 21789 17266 21829
rect 17220 21755 17226 21789
rect 17260 21755 17266 21789
rect 17067 21716 17185 21728
rect 17067 21682 17073 21716
rect 17107 21682 17145 21716
rect 17179 21682 17185 21716
rect 17067 21638 17185 21682
rect 17067 21604 17073 21638
rect 17107 21604 17145 21638
rect 17179 21604 17185 21638
rect 17067 21560 17185 21604
rect 17067 21526 17073 21560
rect 17107 21526 17145 21560
rect 17179 21526 17185 21560
rect 17067 21481 17185 21526
tri 16844 21447 16846 21449 se
rect 16846 21447 17024 21449
tri 16843 21446 16844 21447 se
rect 16844 21446 17024 21447
rect 17067 21447 17073 21481
rect 17107 21447 17145 21481
rect 17179 21447 17185 21481
tri 15627 21402 15631 21406 se
rect 15631 21402 15682 21406
tri 15625 21400 15627 21402 se
rect 15627 21400 15682 21402
rect 16167 21440 17026 21446
rect 16167 21406 16179 21440
rect 16213 21406 16252 21440
rect 16286 21406 16325 21440
rect 16359 21406 16398 21440
rect 16432 21406 16471 21440
rect 16505 21406 16544 21440
rect 16578 21406 16617 21440
rect 16651 21406 16690 21440
rect 16724 21406 16763 21440
rect 16797 21406 16836 21440
rect 16870 21406 16908 21440
rect 16942 21406 16980 21440
rect 17014 21406 17026 21440
rect 16167 21400 17026 21406
rect 17067 21402 17185 21447
tri 15621 21396 15625 21400 se
rect 15625 21396 15682 21400
tri 16843 21397 16846 21400 ne
rect 16846 21397 17024 21400
tri 14759 21377 14778 21396 sw
tri 15614 21389 15621 21396 se
rect 15621 21389 15682 21396
rect 15412 21377 15682 21389
rect 14624 21343 14778 21377
tri 14778 21343 14812 21377 sw
rect 15412 21343 15418 21377
rect 15452 21343 15682 21377
rect 14624 21225 15330 21343
rect 15412 21305 15682 21343
rect 15412 21271 15418 21305
rect 15452 21277 15682 21305
rect 17067 21368 17073 21402
rect 17107 21368 17145 21402
rect 17179 21368 17185 21402
rect 17067 21323 17185 21368
rect 17067 21289 17073 21323
rect 17107 21289 17145 21323
rect 17179 21289 17185 21323
rect 17067 21277 17185 21289
rect 17220 21715 17266 21755
rect 17486 21746 17492 21798
rect 17544 21746 17558 21798
rect 17610 21746 17625 21798
tri 17542 21715 17573 21746 ne
rect 17220 21681 17226 21715
rect 17260 21681 17266 21715
rect 17220 21641 17266 21681
rect 17220 21607 17226 21641
rect 17260 21607 17266 21641
rect 17220 21567 17266 21607
rect 17220 21533 17226 21567
rect 17260 21533 17266 21567
rect 17220 21493 17266 21533
rect 17220 21459 17226 21493
rect 17260 21459 17266 21493
rect 17220 21419 17266 21459
rect 17220 21385 17226 21419
rect 17260 21385 17266 21419
rect 17220 21345 17266 21385
rect 17220 21311 17226 21345
rect 17260 21311 17266 21345
rect 15452 21271 15676 21277
tri 15676 21271 15682 21277 nw
rect 17220 21271 17266 21311
rect 15412 21259 15664 21271
tri 15664 21259 15676 21271 nw
rect 17220 21237 17226 21271
rect 17260 21237 17266 21271
rect 17220 21225 17266 21237
rect 17573 21050 17625 21746
rect 17573 20984 17625 20998
rect 17573 20926 17625 20932
rect 17570 20507 17614 20598
rect 3273 20179 3398 20254
rect 5424 11472 5526 11561
rect 24958 9867 25076 9874
rect 22874 9791 22880 9843
rect 22932 9791 22946 9843
rect 22998 9791 23004 9843
rect 25074 9751 25076 9867
rect 24958 9744 25076 9751
rect 22862 9642 22908 9643
rect 22862 9636 22914 9642
rect 22862 9572 22914 9584
rect 22862 9514 22914 9520
rect 24949 9636 25070 9642
rect 24949 9520 24954 9636
rect 24949 9514 25070 9520
rect 22862 9513 22908 9514
rect 24949 9512 25067 9514
rect 24579 9329 24698 9447
rect 24954 9441 25070 9447
tri 24944 9319 24954 9329 ne
rect 24954 9319 25070 9325
rect 22483 9085 22600 9201
rect 9030 7637 9094 7669
rect 7384 6988 7424 7020
rect 9728 5453 9923 5547
rect 1370 2094 1679 2262
rect 970 1127 1110 1265
tri 6487 -4438 6498 -4427 se
rect 6498 -4438 6549 -4427
rect 6270 -4628 6549 -4438
tri 6445 -4629 6446 -4628 ne
rect 6446 -4629 6549 -4628
rect 6605 -4561 6611 -4509
rect 6663 -4561 6678 -4509
rect 6730 -4561 6745 -4509
rect 6797 -4561 6812 -4509
rect 6864 -4561 6879 -4509
rect 6931 -4561 6945 -4509
rect 6997 -4561 7003 -4509
rect 6605 -4577 7003 -4561
rect 6605 -4629 6611 -4577
rect 6663 -4629 6678 -4577
rect 6730 -4629 6745 -4577
rect 6797 -4629 6812 -4577
rect 6864 -4629 6879 -4577
rect 6931 -4629 6945 -4577
rect 6997 -4629 7003 -4577
rect 3007 -4934 3013 -4882
rect 3065 -4934 3077 -4882
rect 3129 -4934 3135 -4882
rect 12490 -4939 12496 -4887
rect 12548 -4939 12588 -4887
rect 12640 -4939 12680 -4887
rect 12732 -4939 12771 -4887
rect 12823 -4939 12862 -4887
rect 12914 -4939 12920 -4887
rect 12490 -4991 12920 -4939
rect 12490 -5043 12496 -4991
rect 12548 -5043 12588 -4991
rect 12640 -5043 12680 -4991
rect 12732 -5043 12771 -4991
rect 12823 -5043 12862 -4991
rect 12914 -5043 12920 -4991
rect 12490 -5095 12920 -5043
rect 8128 -5153 8134 -5101
rect 8186 -5153 8226 -5101
rect 8278 -5153 8318 -5101
rect 8370 -5153 8376 -5101
rect 12490 -5147 12496 -5095
rect 12548 -5147 12588 -5095
rect 12640 -5147 12680 -5095
rect 12732 -5147 12771 -5095
rect 12823 -5147 12862 -5095
rect 12914 -5147 12920 -5095
rect 10260 -5648 10303 -5610
rect 10548 -5620 10591 -5581
rect 11678 -5712 11739 -5680
rect 4994 -5823 5000 -5771
rect 5052 -5823 5099 -5771
rect 5151 -5823 5197 -5771
rect 5249 -5823 5255 -5771
rect 4994 -5845 5255 -5823
rect 4994 -5897 5000 -5845
rect 5052 -5897 5099 -5845
rect 5151 -5897 5197 -5845
rect 5249 -5897 5255 -5845
rect 4994 -5919 5255 -5897
rect 4994 -5971 5000 -5919
rect 5052 -5971 5099 -5919
rect 5151 -5971 5197 -5919
rect 5249 -5971 5255 -5919
rect 5440 -5825 5446 -5773
rect 5498 -5825 5511 -5773
rect 5440 -5837 5511 -5825
rect 5440 -5889 5446 -5837
rect 5498 -5889 5511 -5837
rect 5440 -5901 5511 -5889
rect 5440 -5953 5446 -5901
rect 5498 -5953 5511 -5901
rect 5755 -5953 5761 -5773
rect 6605 -6403 6611 -6351
rect 6663 -6403 6678 -6351
rect 6730 -6403 6745 -6351
rect 6797 -6403 6812 -6351
rect 6864 -6403 6879 -6351
rect 6931 -6403 6945 -6351
rect 6997 -6403 7003 -6351
rect 6605 -6419 7003 -6403
rect 6605 -6471 6611 -6419
rect 6663 -6471 6678 -6419
rect 6730 -6471 6745 -6419
rect 6797 -6471 6812 -6419
rect 6864 -6471 6879 -6419
rect 6931 -6471 6945 -6419
rect 6997 -6471 7003 -6419
<< via1 >>
rect 17068 23209 17120 23218
rect 17068 23175 17074 23209
rect 17074 23175 17108 23209
rect 17108 23175 17120 23209
rect 17068 23166 17120 23175
rect 17132 23209 17184 23218
rect 17132 23175 17146 23209
rect 17146 23175 17180 23209
rect 17180 23175 17184 23209
rect 17132 23166 17184 23175
rect 17068 23111 17120 23120
rect 17068 23077 17074 23111
rect 17074 23077 17108 23111
rect 17108 23077 17120 23111
rect 17068 23068 17120 23077
rect 17132 23111 17184 23120
rect 17132 23077 17146 23111
rect 17146 23077 17180 23111
rect 17180 23077 17184 23111
rect 17132 23068 17184 23077
rect 16258 22880 16310 22932
rect 16348 22880 16400 22932
rect 16438 22880 16490 22932
rect 16527 22880 16579 22932
rect 17068 22947 17120 22956
rect 17068 22913 17074 22947
rect 17074 22913 17108 22947
rect 17108 22913 17120 22947
rect 17068 22904 17120 22913
rect 17132 22947 17184 22956
rect 17132 22913 17146 22947
rect 17146 22913 17180 22947
rect 17180 22913 17184 22947
rect 17132 22904 17184 22913
rect 16258 22788 16310 22840
rect 16348 22788 16400 22840
rect 16438 22788 16490 22840
rect 16527 22788 16579 22840
rect 16258 22696 16310 22748
rect 16348 22696 16400 22748
rect 16438 22696 16490 22748
rect 16527 22696 16579 22748
rect 16258 22604 16310 22656
rect 16348 22604 16400 22656
rect 16438 22604 16490 22656
rect 16527 22604 16579 22656
rect 14641 21757 14693 21809
rect 14707 21757 14759 21809
rect 14641 21674 14693 21726
rect 14707 21674 14759 21726
rect 14641 21591 14693 21643
rect 14707 21591 14759 21643
rect 14641 21508 14693 21560
rect 14707 21508 14759 21560
rect 16665 21911 16717 21963
rect 16729 21911 16781 21963
rect 16855 21911 16907 21963
rect 16919 21911 16971 21963
rect 16410 21843 16462 21895
rect 16476 21843 16528 21895
rect 17492 21746 17544 21798
rect 17558 21746 17610 21798
rect 17573 20998 17625 21050
rect 17573 20932 17625 20984
rect 24958 9862 25074 9867
rect 22880 9834 22932 9843
rect 22880 9800 22886 9834
rect 22886 9800 22920 9834
rect 22920 9800 22932 9834
rect 22880 9791 22932 9800
rect 22946 9834 22998 9843
rect 22946 9800 22958 9834
rect 22958 9800 22992 9834
rect 22992 9800 22998 9834
rect 22946 9791 22998 9800
rect 24958 9756 24964 9862
rect 24964 9756 25070 9862
rect 25070 9756 25074 9862
rect 24958 9751 25074 9756
rect 22862 9631 22914 9636
rect 22862 9597 22868 9631
rect 22868 9597 22902 9631
rect 22902 9597 22914 9631
rect 22862 9584 22914 9597
rect 22862 9559 22914 9572
rect 22862 9525 22868 9559
rect 22868 9525 22902 9559
rect 22902 9525 22914 9559
rect 22862 9520 22914 9525
rect 24954 9630 25070 9636
rect 24954 9524 24955 9630
rect 24955 9524 25061 9630
rect 25061 9524 25070 9630
rect 24954 9520 25070 9524
rect 24954 9325 25070 9441
rect 6611 -4561 6663 -4509
rect 6678 -4561 6730 -4509
rect 6745 -4561 6797 -4509
rect 6812 -4561 6864 -4509
rect 6879 -4561 6931 -4509
rect 6945 -4561 6997 -4509
rect 6611 -4629 6663 -4577
rect 6678 -4629 6730 -4577
rect 6745 -4629 6797 -4577
rect 6812 -4629 6864 -4577
rect 6879 -4629 6931 -4577
rect 6945 -4629 6997 -4577
rect 3013 -4934 3065 -4882
rect 3077 -4934 3129 -4882
rect 12496 -4939 12548 -4887
rect 12588 -4939 12640 -4887
rect 12680 -4939 12732 -4887
rect 12771 -4939 12823 -4887
rect 12862 -4939 12914 -4887
rect 12496 -5043 12548 -4991
rect 12588 -5043 12640 -4991
rect 12680 -5043 12732 -4991
rect 12771 -5043 12823 -4991
rect 12862 -5043 12914 -4991
rect 8134 -5153 8186 -5101
rect 8226 -5153 8278 -5101
rect 8318 -5153 8370 -5101
rect 12496 -5147 12548 -5095
rect 12588 -5147 12640 -5095
rect 12680 -5147 12732 -5095
rect 12771 -5147 12823 -5095
rect 12862 -5147 12914 -5095
rect 5000 -5823 5052 -5771
rect 5099 -5823 5151 -5771
rect 5197 -5823 5249 -5771
rect 5000 -5897 5052 -5845
rect 5099 -5897 5151 -5845
rect 5197 -5897 5249 -5845
rect 5000 -5971 5052 -5919
rect 5099 -5971 5151 -5919
rect 5197 -5971 5249 -5919
rect 5446 -5825 5498 -5773
rect 5446 -5889 5498 -5837
rect 5446 -5953 5498 -5901
rect 5511 -5953 5755 -5773
rect 6611 -6403 6663 -6351
rect 6678 -6403 6730 -6351
rect 6745 -6403 6797 -6351
rect 6812 -6403 6864 -6351
rect 6879 -6403 6931 -6351
rect 6945 -6403 6997 -6351
rect 6611 -6471 6663 -6419
rect 6678 -6471 6730 -6419
rect 6745 -6471 6797 -6419
rect 6812 -6471 6864 -6419
rect 6879 -6471 6931 -6419
rect 6945 -6471 6997 -6419
<< metal2 >>
rect 18254 23676 18263 23732
rect 18319 23676 18343 23732
rect 18399 23676 18408 23732
tri 16959 23203 16974 23218 se
rect 16974 23203 17068 23218
rect 16959 23166 17068 23203
rect 17120 23166 17132 23218
rect 17184 23166 17190 23218
rect 15752 22922 16258 22932
rect 15752 22866 15768 22922
rect 15824 22866 15899 22922
rect 15955 22866 16030 22922
rect 16086 22866 16161 22922
rect 16217 22880 16258 22922
rect 16310 22880 16348 22932
rect 16400 22880 16438 22932
rect 16490 22880 16527 22932
rect 16579 22880 16585 22932
rect 16217 22866 16585 22880
rect 15752 22840 16585 22866
rect 15752 22796 16258 22840
rect 15752 22740 15768 22796
rect 15824 22740 15899 22796
rect 15955 22740 16030 22796
rect 16086 22740 16161 22796
rect 16217 22788 16258 22796
rect 16310 22788 16348 22840
rect 16400 22788 16438 22840
rect 16490 22788 16527 22840
rect 16579 22788 16585 22840
rect 16217 22748 16585 22788
rect 16217 22740 16258 22748
rect 15752 22696 16258 22740
rect 16310 22696 16348 22748
rect 16400 22696 16438 22748
rect 16490 22696 16527 22748
rect 16579 22696 16585 22748
rect 15752 22670 16585 22696
rect 15752 22614 15768 22670
rect 15824 22614 15899 22670
rect 15955 22614 16030 22670
rect 16086 22614 16161 22670
rect 16217 22656 16585 22670
rect 16217 22614 16258 22656
rect 15752 22604 16258 22614
rect 16310 22604 16348 22656
rect 16400 22604 16438 22656
rect 16490 22604 16527 22656
rect 16579 22604 16585 22656
rect 16959 22637 17011 23166
tri 17011 23136 17041 23166 nw
rect 17062 23068 17068 23120
rect 17120 23068 17132 23120
rect 17184 23068 17208 23120
tri 17186 23054 17200 23068 ne
rect 17200 23054 17208 23068
tri 17208 23054 17274 23120 sw
tri 17200 23046 17208 23054 ne
rect 17208 23046 17274 23054
tri 17208 23032 17222 23046 ne
rect 17062 22904 17068 22956
rect 17120 22904 17132 22956
rect 17184 22904 17190 22956
tri 17102 22868 17138 22904 ne
tri 16959 22632 16964 22637 ne
rect 16964 22632 17011 22637
tri 17011 22632 17042 22663 sw
rect 17138 22649 17190 22904
rect 17222 22740 17274 23046
rect 17780 22816 17836 22825
tri 17274 22740 17290 22756 sw
rect 17222 22734 17290 22740
tri 17222 22727 17229 22734 ne
rect 17229 22727 17290 22734
tri 17290 22727 17303 22740 sw
rect 17780 22736 17836 22760
tri 17229 22682 17274 22727 ne
rect 17274 22682 17780 22727
tri 17274 22671 17285 22682 ne
rect 17285 22680 17780 22682
rect 17285 22671 17836 22680
rect 17906 22731 17962 22740
tri 17190 22649 17212 22671 sw
rect 17906 22651 17962 22675
tri 17138 22632 17155 22649 ne
rect 17155 22642 17212 22649
tri 17212 22642 17219 22649 sw
rect 17155 22632 17906 22642
tri 16964 22604 16992 22632 ne
rect 16992 22604 17042 22632
tri 16992 22585 17011 22604 ne
rect 17011 22586 17042 22604
tri 17042 22586 17088 22632 sw
tri 17155 22586 17201 22632 ne
rect 17201 22595 17906 22632
rect 17201 22586 17962 22595
rect 17011 22585 17088 22586
tri 17011 22554 17042 22585 ne
rect 17042 22554 17088 22585
tri 17088 22554 17120 22586 sw
tri 17042 22498 17098 22554 ne
rect 17098 22545 17708 22554
rect 17098 22498 17652 22545
rect 17652 22465 17708 22489
rect 17652 22400 17708 22409
rect 16643 21909 16652 21965
rect 16708 21963 16732 21965
rect 16717 21911 16729 21963
rect 16708 21909 16732 21911
rect 16788 21909 16797 21965
rect 16849 21963 16858 21965
rect 16914 21963 16938 21965
rect 16849 21911 16855 21963
rect 16914 21911 16919 21963
rect 16849 21909 16858 21911
rect 16914 21909 16938 21911
rect 16994 21909 17003 21965
rect 16400 21843 16410 21895
rect 16462 21843 16476 21895
rect 16528 21843 16584 21895
tri 16584 21843 16636 21895 sw
rect 16400 21839 16636 21843
tri 16636 21839 16640 21843 sw
rect 16400 21835 17616 21839
tri 16558 21815 16578 21835 ne
rect 16578 21815 17616 21835
rect 13852 21809 14774 21815
rect 13852 21805 14641 21809
rect 13852 21749 13861 21805
rect 13917 21749 13949 21805
rect 14005 21749 14037 21805
rect 14093 21749 14125 21805
rect 14181 21749 14213 21805
rect 14269 21749 14300 21805
rect 14356 21749 14387 21805
rect 14443 21757 14641 21805
rect 14693 21757 14707 21809
rect 14759 21757 14774 21809
tri 16578 21798 16595 21815 ne
rect 16595 21798 17616 21815
tri 16595 21787 16606 21798 ne
rect 16606 21787 17492 21798
rect 14443 21749 14774 21757
rect 13852 21726 14774 21749
tri 17445 21746 17486 21787 ne
rect 17486 21746 17492 21787
rect 17544 21746 17558 21798
rect 17610 21746 17616 21798
rect 13852 21689 14641 21726
rect 13852 21633 13861 21689
rect 13917 21633 13949 21689
rect 14005 21633 14037 21689
rect 14093 21633 14125 21689
rect 14181 21633 14213 21689
rect 14269 21633 14300 21689
rect 14356 21633 14387 21689
rect 14443 21674 14641 21689
rect 14693 21674 14707 21726
rect 14759 21674 14774 21726
rect 14443 21643 14774 21674
rect 14443 21633 14641 21643
rect 13852 21591 14641 21633
rect 14693 21591 14707 21643
rect 14759 21591 14774 21643
rect 13852 21573 14774 21591
rect 17302 21575 17311 21711
rect 17447 21575 17456 21711
rect 13852 21517 13861 21573
rect 13917 21517 13949 21573
rect 14005 21517 14037 21573
rect 14093 21517 14125 21573
rect 14181 21517 14213 21573
rect 14269 21517 14300 21573
rect 14356 21517 14387 21573
rect 14443 21560 14774 21573
rect 14443 21517 14641 21560
rect 13852 21508 14641 21517
rect 14693 21508 14707 21560
rect 14759 21508 14774 21560
rect 13852 21502 14774 21508
rect 17310 21315 17377 21367
rect 17310 21235 17378 21275
rect 17573 21050 17625 21056
tri 17568 20998 17573 21003 se
tri 17554 20984 17568 20998 se
rect 17568 20984 17625 20998
tri 17533 20963 17554 20984 se
rect 17554 20963 17573 20984
tri 6281 20932 6312 20963 se
rect 6312 20932 17573 20963
tri 6275 20926 6281 20932 se
rect 6281 20926 17625 20932
tri 6217 20868 6275 20926 se
rect 6275 20868 6312 20926
tri 6312 20868 6370 20926 nw
tri 6185 20836 6217 20868 se
rect 6217 20836 6280 20868
tri 6280 20836 6312 20868 nw
rect 17308 20844 17377 20896
rect 3017 20790 6234 20836
tri 6234 20790 6280 20836 nw
rect 3017 20752 3174 20790
rect 3103 20244 3174 20752
tri 3174 20751 3213 20790 nw
rect 17306 20177 17391 20255
rect 24958 9867 25074 9873
rect 22874 9791 22880 9843
rect 22932 9791 22946 9843
rect 22998 9791 23004 9843
rect 24958 9745 25074 9751
rect 22844 9663 22900 9672
rect 22900 9636 22914 9642
rect 22844 9584 22862 9607
rect 22844 9583 22914 9584
rect 22900 9572 22914 9583
rect 22844 9520 22862 9527
rect 22844 9518 22914 9520
rect 22862 9514 22914 9518
rect 24954 9636 25070 9642
rect 24954 9514 25070 9520
rect 24954 9464 25074 9473
rect 24954 9441 24986 9464
rect 25042 9441 25074 9464
rect 25070 9325 25074 9441
rect 24954 9319 25074 9325
rect 1891 7803 1943 7841
rect 1799 7756 1851 7790
rect 2520 7745 2572 7785
rect 2075 6895 2127 6945
rect 1799 6793 1851 6848
rect 1523 5869 1575 5947
rect 1853 3279 1880 3306
tri 12608 553 12702 647 se
rect 12702 637 16399 647
rect 12702 608 16254 637
tri 12702 553 12757 608 nw
tri 16203 581 16230 608 ne
rect 16230 581 16254 608
rect 16310 581 16334 637
rect 16390 581 16399 637
rect 16451 581 16460 637
rect 16516 581 16540 637
rect 16596 605 17220 637
tri 17220 605 17252 637 sw
rect 16596 581 17252 605
tri 17166 553 17194 581 ne
rect 17194 553 17252 581
tri 12514 459 12608 553 se
tri 12608 459 12702 553 nw
tri 17194 549 17198 553 ne
tri 12455 400 12514 459 se
rect 12514 400 12549 459
tri 12549 400 12608 459 nw
rect 12455 301 12511 400
tri 12511 362 12549 400 nw
tri 17169 -575 17198 -546 se
rect 17198 -575 17252 553
tri 17252 -575 17281 -546 sw
rect 6605 -4561 6611 -4509
rect 6663 -4542 6678 -4509
rect 6730 -4542 6745 -4509
rect 6797 -4542 6812 -4509
rect 6864 -4542 6879 -4509
rect 6931 -4542 6945 -4509
rect 6671 -4561 6678 -4542
rect 6931 -4561 6937 -4542
rect 6997 -4561 7003 -4509
rect 6605 -4577 6615 -4561
rect 6671 -4577 6696 -4561
rect 6752 -4577 6777 -4561
rect 6833 -4577 6857 -4561
rect 6913 -4577 6937 -4561
rect 6993 -4577 7003 -4561
rect 6605 -4629 6611 -4577
rect 6671 -4598 6678 -4577
rect 6931 -4598 6937 -4577
rect 6663 -4629 6678 -4598
rect 6730 -4629 6745 -4598
rect 6797 -4629 6812 -4598
rect 6864 -4629 6879 -4598
rect 6931 -4629 6945 -4598
rect 6997 -4629 7003 -4577
rect 3016 -4856 3072 -4847
rect 3007 -4934 3013 -4882
rect 3072 -4912 3077 -4882
rect 3065 -4934 3077 -4912
rect 3129 -4934 3135 -4882
rect 12485 -4885 12927 -4884
rect 3016 -4936 3072 -4934
rect 3016 -5001 3072 -4992
rect 12485 -4941 12494 -4885
rect 12550 -4887 12617 -4885
rect 12673 -4887 12740 -4885
rect 12796 -4887 12862 -4885
rect 12550 -4939 12588 -4887
rect 12673 -4939 12680 -4887
rect 12732 -4939 12740 -4887
rect 12823 -4939 12862 -4887
rect 12550 -4941 12617 -4939
rect 12673 -4941 12740 -4939
rect 12796 -4941 12862 -4939
rect 12918 -4941 12927 -4885
rect 12485 -4989 12927 -4941
rect 12485 -5045 12494 -4989
rect 12550 -4991 12617 -4989
rect 12673 -4991 12740 -4989
rect 12796 -4991 12862 -4989
rect 12550 -5043 12588 -4991
rect 12673 -5043 12680 -4991
rect 12732 -5043 12740 -4991
rect 12823 -5043 12862 -4991
rect 12550 -5045 12617 -5043
rect 12673 -5045 12740 -5043
rect 12796 -5045 12862 -5043
rect 12918 -5045 12927 -4989
rect 12485 -5093 12927 -5045
rect 8114 -5155 8123 -5099
rect 8179 -5101 8220 -5099
rect 8276 -5101 8316 -5099
rect 8186 -5153 8220 -5101
rect 8278 -5153 8316 -5101
rect 8179 -5155 8220 -5153
rect 8276 -5155 8316 -5153
rect 8372 -5155 8381 -5099
rect 12485 -5149 12494 -5093
rect 12550 -5095 12617 -5093
rect 12673 -5095 12740 -5093
rect 12796 -5095 12862 -5093
rect 12550 -5147 12588 -5095
rect 12673 -5147 12680 -5095
rect 12732 -5147 12740 -5095
rect 12823 -5147 12862 -5095
rect 12550 -5149 12617 -5147
rect 12673 -5149 12740 -5147
rect 12796 -5149 12862 -5147
rect 12918 -5149 12927 -5093
rect 12485 -5150 12927 -5149
rect 4981 -5812 4990 -5756
rect 5046 -5771 5101 -5756
rect 5157 -5771 5212 -5756
rect 4981 -5823 5000 -5812
rect 5052 -5823 5099 -5771
rect 5157 -5812 5197 -5771
rect 5268 -5812 5277 -5756
rect 5151 -5823 5197 -5812
rect 5249 -5823 5277 -5812
rect 4981 -5840 5277 -5823
rect 4981 -5896 4990 -5840
rect 5046 -5845 5101 -5840
rect 5157 -5845 5212 -5840
rect 4981 -5897 5000 -5896
rect 5052 -5897 5099 -5845
rect 5157 -5896 5197 -5845
rect 5268 -5896 5277 -5840
rect 5151 -5897 5197 -5896
rect 5249 -5897 5277 -5896
rect 4981 -5919 5277 -5897
rect 4981 -5924 5000 -5919
rect 4981 -5980 4990 -5924
rect 5052 -5971 5099 -5919
rect 5151 -5924 5197 -5919
rect 5249 -5924 5277 -5919
rect 5157 -5971 5197 -5924
rect 5046 -5980 5101 -5971
rect 5157 -5980 5212 -5971
rect 5268 -5980 5277 -5924
rect 5433 -5829 5442 -5773
rect 5498 -5829 5511 -5773
rect 5761 -5829 5770 -5773
rect 8198 -5785 8304 -5776
rect 8198 -5794 8223 -5785
rect 5433 -5837 5511 -5829
rect 5433 -5889 5446 -5837
rect 5498 -5889 5511 -5837
rect 5433 -5897 5511 -5889
rect 5755 -5897 5770 -5829
rect 8166 -5841 8223 -5794
rect 8279 -5841 8304 -5785
rect 8166 -5846 8304 -5841
tri 8166 -5873 8193 -5846 ne
rect 8193 -5865 8304 -5846
rect 5433 -5953 5442 -5897
rect 5498 -5953 5511 -5897
rect 5761 -5953 5770 -5897
rect 8193 -5921 8223 -5865
rect 8279 -5921 8304 -5865
rect 8193 -5922 8304 -5921
rect 8198 -5930 8304 -5922
rect 6605 -6403 6611 -6351
rect 6663 -6383 6678 -6351
rect 6730 -6383 6745 -6351
rect 6797 -6383 6812 -6351
rect 6864 -6383 6879 -6351
rect 6931 -6383 6945 -6351
rect 6671 -6403 6678 -6383
rect 6931 -6403 6937 -6383
rect 6997 -6403 7003 -6351
rect 6605 -6419 6615 -6403
rect 6671 -6419 6696 -6403
rect 6752 -6419 6777 -6403
rect 6833 -6419 6857 -6403
rect 6913 -6419 6937 -6403
rect 6993 -6419 7003 -6403
rect 6605 -6471 6611 -6419
rect 6671 -6439 6678 -6419
rect 6931 -6439 6937 -6419
rect 6663 -6471 6678 -6439
rect 6730 -6471 6745 -6439
rect 6797 -6471 6812 -6439
rect 6864 -6471 6879 -6439
rect 6931 -6471 6945 -6439
rect 6997 -6471 7003 -6419
<< via2 >>
rect 18263 23676 18319 23732
rect 18343 23676 18399 23732
rect 15768 22866 15824 22922
rect 15899 22866 15955 22922
rect 16030 22866 16086 22922
rect 16161 22866 16217 22922
rect 15768 22740 15824 22796
rect 15899 22740 15955 22796
rect 16030 22740 16086 22796
rect 16161 22740 16217 22796
rect 15768 22614 15824 22670
rect 15899 22614 15955 22670
rect 16030 22614 16086 22670
rect 16161 22614 16217 22670
rect 17780 22760 17836 22816
rect 17780 22680 17836 22736
rect 17906 22675 17962 22731
rect 17906 22595 17962 22651
rect 17652 22489 17708 22545
rect 17652 22409 17708 22465
rect 16652 21963 16708 21965
rect 16732 21963 16788 21965
rect 16652 21911 16665 21963
rect 16665 21911 16708 21963
rect 16732 21911 16781 21963
rect 16781 21911 16788 21963
rect 16652 21909 16708 21911
rect 16732 21909 16788 21911
rect 16858 21963 16914 21965
rect 16938 21963 16994 21965
rect 16858 21911 16907 21963
rect 16907 21911 16914 21963
rect 16938 21911 16971 21963
rect 16971 21911 16994 21963
rect 16858 21909 16914 21911
rect 16938 21909 16994 21911
rect 13861 21749 13917 21805
rect 13949 21749 14005 21805
rect 14037 21749 14093 21805
rect 14125 21749 14181 21805
rect 14213 21749 14269 21805
rect 14300 21749 14356 21805
rect 14387 21749 14443 21805
rect 13861 21633 13917 21689
rect 13949 21633 14005 21689
rect 14037 21633 14093 21689
rect 14125 21633 14181 21689
rect 14213 21633 14269 21689
rect 14300 21633 14356 21689
rect 14387 21633 14443 21689
rect 17311 21575 17447 21711
rect 13861 21517 13917 21573
rect 13949 21517 14005 21573
rect 14037 21517 14093 21573
rect 14125 21517 14181 21573
rect 14213 21517 14269 21573
rect 14300 21517 14356 21573
rect 14387 21517 14443 21573
rect 22844 9636 22900 9663
rect 22844 9607 22862 9636
rect 22862 9607 22900 9636
rect 22844 9572 22900 9583
rect 22844 9527 22862 9572
rect 22862 9527 22900 9572
rect 24986 9441 25042 9464
rect 24986 9408 25042 9441
rect 24986 9328 25042 9384
rect 16254 581 16310 637
rect 16334 581 16390 637
rect 16460 581 16516 637
rect 16540 581 16596 637
rect 6615 -4561 6663 -4542
rect 6663 -4561 6671 -4542
rect 6696 -4561 6730 -4542
rect 6730 -4561 6745 -4542
rect 6745 -4561 6752 -4542
rect 6777 -4561 6797 -4542
rect 6797 -4561 6812 -4542
rect 6812 -4561 6833 -4542
rect 6857 -4561 6864 -4542
rect 6864 -4561 6879 -4542
rect 6879 -4561 6913 -4542
rect 6937 -4561 6945 -4542
rect 6945 -4561 6993 -4542
rect 6615 -4577 6671 -4561
rect 6696 -4577 6752 -4561
rect 6777 -4577 6833 -4561
rect 6857 -4577 6913 -4561
rect 6937 -4577 6993 -4561
rect 6615 -4598 6663 -4577
rect 6663 -4598 6671 -4577
rect 6696 -4598 6730 -4577
rect 6730 -4598 6745 -4577
rect 6745 -4598 6752 -4577
rect 6777 -4598 6797 -4577
rect 6797 -4598 6812 -4577
rect 6812 -4598 6833 -4577
rect 6857 -4598 6864 -4577
rect 6864 -4598 6879 -4577
rect 6879 -4598 6913 -4577
rect 6937 -4598 6945 -4577
rect 6945 -4598 6993 -4577
rect 3016 -4882 3072 -4856
rect 3016 -4912 3065 -4882
rect 3065 -4912 3072 -4882
rect 3016 -4992 3072 -4936
rect 12494 -4887 12550 -4885
rect 12617 -4887 12673 -4885
rect 12740 -4887 12796 -4885
rect 12862 -4887 12918 -4885
rect 12494 -4939 12496 -4887
rect 12496 -4939 12548 -4887
rect 12548 -4939 12550 -4887
rect 12617 -4939 12640 -4887
rect 12640 -4939 12673 -4887
rect 12740 -4939 12771 -4887
rect 12771 -4939 12796 -4887
rect 12862 -4939 12914 -4887
rect 12914 -4939 12918 -4887
rect 12494 -4941 12550 -4939
rect 12617 -4941 12673 -4939
rect 12740 -4941 12796 -4939
rect 12862 -4941 12918 -4939
rect 12494 -4991 12550 -4989
rect 12617 -4991 12673 -4989
rect 12740 -4991 12796 -4989
rect 12862 -4991 12918 -4989
rect 12494 -5043 12496 -4991
rect 12496 -5043 12548 -4991
rect 12548 -5043 12550 -4991
rect 12617 -5043 12640 -4991
rect 12640 -5043 12673 -4991
rect 12740 -5043 12771 -4991
rect 12771 -5043 12796 -4991
rect 12862 -5043 12914 -4991
rect 12914 -5043 12918 -4991
rect 12494 -5045 12550 -5043
rect 12617 -5045 12673 -5043
rect 12740 -5045 12796 -5043
rect 12862 -5045 12918 -5043
rect 8123 -5101 8179 -5099
rect 8220 -5101 8276 -5099
rect 8316 -5101 8372 -5099
rect 8123 -5153 8134 -5101
rect 8134 -5153 8179 -5101
rect 8220 -5153 8226 -5101
rect 8226 -5153 8276 -5101
rect 8316 -5153 8318 -5101
rect 8318 -5153 8370 -5101
rect 8370 -5153 8372 -5101
rect 8123 -5155 8179 -5153
rect 8220 -5155 8276 -5153
rect 8316 -5155 8372 -5153
rect 12494 -5095 12550 -5093
rect 12617 -5095 12673 -5093
rect 12740 -5095 12796 -5093
rect 12862 -5095 12918 -5093
rect 12494 -5147 12496 -5095
rect 12496 -5147 12548 -5095
rect 12548 -5147 12550 -5095
rect 12617 -5147 12640 -5095
rect 12640 -5147 12673 -5095
rect 12740 -5147 12771 -5095
rect 12771 -5147 12796 -5095
rect 12862 -5147 12914 -5095
rect 12914 -5147 12918 -5095
rect 12494 -5149 12550 -5147
rect 12617 -5149 12673 -5147
rect 12740 -5149 12796 -5147
rect 12862 -5149 12918 -5147
rect 4990 -5771 5046 -5756
rect 5101 -5771 5157 -5756
rect 5212 -5771 5268 -5756
rect 4990 -5812 5000 -5771
rect 5000 -5812 5046 -5771
rect 5101 -5812 5151 -5771
rect 5151 -5812 5157 -5771
rect 5212 -5812 5249 -5771
rect 5249 -5812 5268 -5771
rect 4990 -5845 5046 -5840
rect 5101 -5845 5157 -5840
rect 5212 -5845 5268 -5840
rect 4990 -5896 5000 -5845
rect 5000 -5896 5046 -5845
rect 5101 -5896 5151 -5845
rect 5151 -5896 5157 -5845
rect 5212 -5896 5249 -5845
rect 5249 -5896 5268 -5845
rect 4990 -5971 5000 -5924
rect 5000 -5971 5046 -5924
rect 5101 -5971 5151 -5924
rect 5151 -5971 5157 -5924
rect 5212 -5971 5249 -5924
rect 5249 -5971 5268 -5924
rect 4990 -5980 5046 -5971
rect 5101 -5980 5157 -5971
rect 5212 -5980 5268 -5971
rect 5442 -5825 5446 -5773
rect 5446 -5825 5498 -5773
rect 5442 -5829 5498 -5825
rect 5530 -5829 5586 -5773
rect 5618 -5829 5674 -5773
rect 5705 -5829 5755 -5773
rect 5755 -5829 5761 -5773
rect 8223 -5841 8279 -5785
rect 5442 -5901 5498 -5897
rect 5442 -5953 5446 -5901
rect 5446 -5953 5498 -5901
rect 5530 -5953 5586 -5897
rect 5618 -5953 5674 -5897
rect 5705 -5953 5755 -5897
rect 5755 -5953 5761 -5897
rect 8223 -5921 8279 -5865
rect 6615 -6403 6663 -6383
rect 6663 -6403 6671 -6383
rect 6696 -6403 6730 -6383
rect 6730 -6403 6745 -6383
rect 6745 -6403 6752 -6383
rect 6777 -6403 6797 -6383
rect 6797 -6403 6812 -6383
rect 6812 -6403 6833 -6383
rect 6857 -6403 6864 -6383
rect 6864 -6403 6879 -6383
rect 6879 -6403 6913 -6383
rect 6937 -6403 6945 -6383
rect 6945 -6403 6993 -6383
rect 6615 -6419 6671 -6403
rect 6696 -6419 6752 -6403
rect 6777 -6419 6833 -6403
rect 6857 -6419 6913 -6403
rect 6937 -6419 6993 -6403
rect 6615 -6439 6663 -6419
rect 6663 -6439 6671 -6419
rect 6696 -6439 6730 -6419
rect 6730 -6439 6745 -6419
rect 6745 -6439 6752 -6419
rect 6777 -6439 6797 -6419
rect 6797 -6439 6812 -6419
rect 6812 -6439 6833 -6419
rect 6857 -6439 6864 -6419
rect 6864 -6439 6879 -6419
rect 6879 -6439 6913 -6419
rect 6937 -6439 6945 -6419
rect 6945 -6439 6993 -6419
<< metal3 >>
rect 18258 23732 18404 23737
rect 18258 23676 18263 23732
rect 18319 23676 18343 23732
rect 18399 23676 18404 23732
rect 18258 23671 18404 23676
rect 15763 22922 16222 22928
rect 15763 22866 15768 22922
rect 15824 22866 15899 22922
rect 15955 22866 16030 22922
rect 16086 22866 16161 22922
rect 16217 22866 16222 22922
rect 15763 22796 16222 22866
rect 15763 22740 15768 22796
rect 15824 22740 15899 22796
rect 15955 22740 16030 22796
rect 16086 22740 16161 22796
rect 16217 22740 16222 22796
rect 15763 22670 16222 22740
rect 17775 22816 17841 22821
rect 17775 22760 17780 22816
rect 17836 22760 17841 22816
rect 17775 22736 17841 22760
rect 17775 22680 17780 22736
rect 17836 22680 17841 22736
rect 17775 22675 17841 22680
rect 17901 22731 17967 22736
rect 17901 22675 17906 22731
rect 17962 22675 17967 22731
rect 15763 22614 15768 22670
rect 15824 22614 15899 22670
rect 15955 22614 16030 22670
rect 16086 22614 16161 22670
rect 16217 22614 16222 22670
rect 15763 22608 16222 22614
rect 17901 22651 17967 22675
rect 17901 22595 17906 22651
rect 17962 22595 17967 22651
rect 17901 22590 17967 22595
rect 17647 22545 17713 22550
rect 17647 22489 17652 22545
rect 17708 22489 17713 22545
rect 17647 22465 17713 22489
rect 17647 22409 17652 22465
rect 17708 22409 17713 22465
rect 17647 22404 17713 22409
tri 16776 22096 16816 22136 se
rect 16816 22096 17105 22136
tri 17105 22096 17145 22136 sw
tri 16715 22035 16776 22096 se
rect 16776 22069 17145 22096
rect 16776 22035 16816 22069
tri 16816 22035 16850 22069 nw
tri 17045 22035 17079 22069 ne
rect 17079 22035 17145 22069
tri 16650 21970 16715 22035 se
rect 16715 21970 16793 22035
tri 16793 22012 16816 22035 nw
tri 17079 22029 17085 22035 ne
rect 16647 21965 16793 21970
rect 16647 21909 16652 21965
rect 16708 21909 16732 21965
rect 16788 21909 16793 21965
rect 16647 21904 16793 21909
rect 16853 21965 17000 21970
rect 16853 21909 16858 21965
rect 16914 21909 16938 21965
rect 16994 21909 17000 21965
rect 16853 21904 17000 21909
tri 16885 21856 16933 21904 ne
rect 16933 21856 17000 21904
rect 17085 21873 17145 22035
tri 17145 21873 17155 21883 sw
rect 17085 21857 17155 21873
tri 17085 21856 17086 21857 ne
rect 17086 21856 17155 21857
tri 17155 21856 17172 21873 sw
tri 16933 21849 16940 21856 ne
rect 16940 21830 17000 21856
tri 16940 21821 16949 21830 ne
rect 16949 21821 17000 21830
tri 17000 21821 17035 21856 sw
tri 17086 21821 17121 21856 ne
rect 17121 21821 17172 21856
tri 17172 21821 17207 21856 sw
tri 16949 21811 16959 21821 ne
rect 16959 21811 17035 21821
tri 17035 21811 17045 21821 sw
tri 17121 21811 17131 21821 ne
rect 17131 21811 17207 21821
tri 17207 21811 17217 21821 sw
rect 13856 21805 14448 21811
rect 13856 21749 13861 21805
rect 13917 21749 13949 21805
rect 14005 21749 14037 21805
rect 14093 21749 14125 21805
rect 14181 21749 14213 21805
rect 14269 21749 14300 21805
rect 14356 21749 14387 21805
rect 14443 21749 14448 21805
tri 16959 21770 17000 21811 ne
rect 17000 21787 17045 21811
tri 17045 21787 17069 21811 sw
tri 17131 21787 17155 21811 ne
rect 17155 21787 17217 21811
tri 17217 21787 17241 21811 sw
rect 17000 21770 17069 21787
rect 13856 21689 14448 21749
tri 17000 21735 17035 21770 ne
rect 17035 21735 17069 21770
tri 17069 21735 17121 21787 sw
tri 17155 21761 17181 21787 ne
tri 17035 21716 17054 21735 ne
rect 17054 21716 17121 21735
tri 17054 21711 17059 21716 ne
rect 17059 21711 17121 21716
tri 17059 21709 17061 21711 ne
rect 13856 21633 13861 21689
rect 13917 21633 13949 21689
rect 14005 21633 14037 21689
rect 14093 21633 14125 21689
rect 14181 21633 14213 21689
rect 14269 21633 14300 21689
rect 14356 21633 14387 21689
rect 14443 21633 14448 21689
rect 13856 21573 14448 21633
rect 13856 21517 13861 21573
rect 13917 21517 13949 21573
rect 14005 21517 14037 21573
rect 14093 21517 14125 21573
rect 14181 21517 14213 21573
rect 14269 21517 14300 21573
rect 14356 21517 14387 21573
rect 14443 21517 14448 21573
rect 13856 21511 14448 21517
tri 17010 9607 17061 9658 se
rect 17061 9632 17121 21711
rect 17061 9607 17096 9632
tri 17096 9607 17121 9632 nw
tri 16986 9583 17010 9607 se
rect 17010 9606 17095 9607
tri 17095 9606 17096 9607 nw
rect 17010 9583 17072 9606
tri 17072 9583 17095 9606 nw
tri 17158 9583 17181 9606 se
rect 17181 9583 17241 21787
rect 17306 21711 17452 21716
rect 17306 21703 17311 21711
rect 17447 21703 17452 21711
rect 17306 21603 17311 21639
rect 17447 21603 17452 21639
rect 17370 21539 17388 21575
rect 17306 21503 17452 21539
rect 17370 21439 17388 21503
rect 17306 21403 17452 21439
rect 17370 21339 17388 21403
rect 17306 21303 17452 21339
rect 17370 21239 17388 21303
rect 17306 21233 17452 21239
tri 22377 21660 22382 21665 se
rect 22382 21660 22682 21665
tri 22682 21660 22687 21665 sw
rect 22377 21174 22687 21660
tri 22377 21169 22382 21174 ne
rect 22382 21169 22682 21174
tri 22682 21169 22687 21174 nw
tri 22377 20314 22382 20319 se
rect 22382 20314 22682 20319
tri 22682 20314 22687 20319 sw
rect 22377 19828 22687 20314
tri 22377 19827 22378 19828 ne
rect 22378 19827 22686 19828
tri 22686 19827 22687 19828 nw
rect 23036 10304 23183 10322
rect 23100 10240 23118 10304
rect 23182 10240 23183 10304
rect 23036 10222 23183 10240
rect 23100 10158 23118 10222
rect 23182 10158 23183 10222
rect 23036 10139 23183 10158
rect 23100 10075 23118 10139
rect 23182 10075 23183 10139
rect 23036 10056 23183 10075
rect 23100 9992 23118 10056
rect 23182 9992 23183 10056
rect 23036 9973 23183 9992
rect 23100 9909 23118 9973
rect 23182 9909 23183 9973
rect 23036 9890 23183 9909
rect 23100 9826 23118 9890
rect 23182 9826 23183 9890
rect 23036 9807 23183 9826
rect 23100 9743 23118 9807
rect 23182 9743 23183 9807
rect 23036 9724 23183 9743
tri 16975 9572 16986 9583 se
rect 16986 9572 17061 9583
tri 17061 9572 17072 9583 nw
tri 17147 9572 17158 9583 se
rect 17158 9580 17241 9583
rect 17158 9572 17188 9580
tri 16930 9527 16975 9572 se
rect 16975 9527 17016 9572
tri 17016 9527 17061 9572 nw
tri 17102 9527 17147 9572 se
rect 17147 9527 17188 9572
tri 17188 9527 17241 9580 nw
rect 22839 9663 22905 9668
rect 22839 9607 22844 9663
rect 22900 9607 22905 9663
rect 22839 9583 22905 9607
rect 22839 9527 22844 9583
rect 22900 9527 22905 9583
tri 16889 9486 16930 9527 se
rect 16930 9520 17009 9527
tri 17009 9520 17016 9527 nw
tri 17095 9520 17102 9527 se
rect 17102 9520 17181 9527
tri 17181 9520 17188 9527 nw
rect 22839 9522 22905 9527
rect 23100 9660 23118 9724
rect 23182 9660 23183 9724
rect 23036 9641 23183 9660
rect 23100 9577 23118 9641
rect 23182 9577 23183 9641
rect 16930 9486 16975 9520
tri 16975 9486 17009 9520 nw
tri 17061 9486 17095 9520 se
rect 17095 9486 17125 9520
tri 16867 9464 16889 9486 se
rect 16889 9464 16953 9486
tri 16953 9464 16975 9486 nw
tri 17039 9464 17061 9486 se
rect 17061 9464 17125 9486
tri 17125 9464 17181 9520 nw
tri 16811 9408 16867 9464 se
rect 16867 9434 16923 9464
tri 16923 9434 16953 9464 nw
tri 17009 9434 17039 9464 se
rect 17039 9434 17095 9464
tri 17095 9434 17125 9464 nw
rect 16867 9408 16897 9434
tri 16897 9408 16923 9434 nw
tri 16983 9408 17009 9434 se
rect 17009 9408 17069 9434
tri 17069 9408 17095 9434 nw
tri 16803 9400 16811 9408 se
rect 16811 9400 16889 9408
tri 16889 9400 16897 9408 nw
tri 16975 9400 16983 9408 se
rect 16983 9400 17045 9408
tri 16787 9384 16803 9400 se
rect 16803 9384 16873 9400
tri 16873 9384 16889 9400 nw
tri 16959 9384 16975 9400 se
rect 16975 9384 17045 9400
tri 17045 9384 17069 9408 nw
tri 16731 9328 16787 9384 se
rect 16787 9348 16837 9384
tri 16837 9348 16873 9384 nw
tri 16923 9348 16959 9384 se
rect 16959 9348 17009 9384
tri 17009 9348 17045 9384 nw
rect 16787 9328 16817 9348
tri 16817 9328 16837 9348 nw
tri 16903 9328 16923 9348 se
rect 16923 9328 16989 9348
tri 16989 9328 17009 9348 nw
tri 16717 9314 16731 9328 se
rect 16731 9314 16803 9328
tri 16803 9314 16817 9328 nw
tri 16889 9314 16903 9328 se
rect 16903 9314 16923 9328
tri 16631 9228 16717 9314 se
rect 16717 9262 16751 9314
tri 16751 9262 16803 9314 nw
tri 16837 9262 16889 9314 se
rect 16889 9262 16923 9314
tri 16923 9262 16989 9328 nw
tri 16717 9228 16751 9262 nw
tri 16803 9228 16837 9262 se
tri 16545 9142 16631 9228 se
rect 16631 9176 16665 9228
tri 16665 9176 16717 9228 nw
tri 16751 9176 16803 9228 se
rect 16803 9176 16837 9228
tri 16837 9176 16923 9262 nw
tri 16631 9142 16665 9176 nw
tri 16717 9142 16751 9176 se
tri 16459 9056 16545 9142 se
rect 16545 9090 16579 9142
tri 16579 9090 16631 9142 nw
tri 16665 9090 16717 9142 se
rect 16717 9090 16751 9142
tri 16751 9090 16837 9176 nw
tri 16545 9056 16579 9090 nw
tri 16631 9056 16665 9090 se
tri 16373 8970 16459 9056 se
rect 16459 9004 16493 9056
tri 16493 9004 16545 9056 nw
tri 16579 9004 16631 9056 se
rect 16631 9004 16665 9056
tri 16665 9004 16751 9090 nw
tri 16459 8970 16493 9004 nw
tri 16545 8970 16579 9004 se
tri 16287 8884 16373 8970 se
rect 16373 8918 16407 8970
tri 16407 8918 16459 8970 nw
tri 16493 8918 16545 8970 se
rect 16545 8918 16579 8970
tri 16579 8918 16665 9004 nw
tri 16373 8884 16407 8918 nw
tri 16459 8884 16493 8918 se
tri 16230 8827 16287 8884 se
rect 16287 8832 16321 8884
tri 16321 8832 16373 8884 nw
tri 16407 8832 16459 8884 se
rect 16459 8832 16493 8884
tri 16493 8832 16579 8918 nw
rect 16287 8827 16316 8832
tri 16316 8827 16321 8832 nw
tri 16402 8827 16407 8832 se
rect 16407 8827 16436 8832
rect 16230 3811 16290 8827
tri 16290 8801 16316 8827 nw
tri 16376 8801 16402 8827 se
rect 16402 8801 16436 8827
tri 16350 8775 16376 8801 se
rect 16376 8775 16436 8801
tri 16436 8775 16493 8832 nw
rect 16350 3863 16410 8775
tri 16410 8749 16436 8775 nw
tri 16410 3863 16436 3889 sw
tri 16350 3837 16376 3863 ne
rect 16376 3837 16436 3863
tri 16290 3811 16316 3837 sw
tri 16376 3811 16402 3837 ne
rect 16402 3811 16436 3837
tri 16230 3725 16316 3811 ne
tri 16316 3777 16350 3811 sw
tri 16402 3777 16436 3811 ne
tri 16436 3798 16501 3863 sw
rect 16436 3777 16501 3798
rect 16316 3746 16350 3777
tri 16350 3746 16381 3777 sw
tri 16436 3772 16441 3777 ne
rect 16316 3725 16381 3746
tri 16316 3720 16321 3725 ne
rect 16321 1308 16381 3725
rect 16441 1428 16501 3777
tri 16501 1428 16515 1442 sw
rect 16441 1368 16515 1428
tri 16441 1354 16455 1368 ne
tri 16381 1308 16395 1322 sw
rect 11713 1167 12602 1295
rect 16321 1248 16395 1308
tri 16321 1234 16335 1248 ne
tri 11713 1096 11784 1167 ne
rect 3003 -4856 3089 646
rect 3003 -4912 3016 -4856
rect 3072 -4912 3089 -4856
rect 3003 -4936 3089 -4912
rect 3003 -4992 3016 -4936
rect 3072 -4992 3089 -4936
rect 3003 -5049 3089 -4992
tri 3128 -6314 3151 -6291 se
rect 3151 -6380 3237 646
rect 11784 129 12602 1167
tri 16275 642 16335 702 se
rect 16335 642 16395 1248
rect 16249 637 16395 642
rect 16249 581 16254 637
rect 16310 581 16334 637
rect 16390 581 16395 637
rect 16249 576 16395 581
rect 16455 642 16515 1368
tri 16515 642 16572 699 sw
rect 16455 637 16601 642
rect 16455 581 16460 637
rect 16516 581 16540 637
rect 16596 581 16601 637
rect 16455 576 16601 581
tri 22873 149 23036 312 se
rect 23036 151 23183 9577
rect 24949 9464 25079 9469
rect 24949 9408 24986 9464
rect 25042 9408 25079 9464
rect 24949 9384 25079 9408
rect 24949 9328 24986 9384
rect 25042 9328 25079 9384
rect 24949 9323 25079 9328
rect 23036 149 23040 151
rect 23161 149 23181 151
tri 23181 149 23183 151 nw
rect 23161 139 23171 149
tri 23171 139 23181 149 nw
tri 12602 129 12612 139 sw
tri 23161 129 23171 139 nw
rect 11784 85 12612 129
tri 11784 -197 12066 85 ne
rect 12066 -197 12612 85
tri 12612 -197 12938 129 sw
tri 12066 -612 12481 -197 ne
rect 4917 -4941 5246 -4487
rect 6610 -4542 6998 -4507
rect 6610 -4598 6615 -4542
rect 6671 -4598 6696 -4542
rect 6752 -4598 6777 -4542
rect 6833 -4598 6857 -4542
rect 6913 -4598 6937 -4542
rect 6993 -4598 6998 -4542
tri 5246 -4941 5249 -4938 sw
rect 4917 -4989 5249 -4941
tri 5249 -4989 5297 -4941 sw
rect 4917 -4994 5297 -4989
tri 5297 -4994 5302 -4989 sw
rect 4917 -5045 5302 -4994
tri 5302 -5045 5353 -4994 sw
rect 4917 -5073 5353 -5045
tri 4917 -5093 4937 -5073 ne
rect 4937 -5093 5353 -5073
tri 5353 -5093 5401 -5045 sw
tri 4937 -5099 4943 -5093 ne
rect 4943 -5099 5401 -5093
tri 5401 -5099 5407 -5093 sw
tri 4943 -5155 4999 -5099 ne
rect 4999 -5155 5407 -5099
tri 5407 -5155 5463 -5099 sw
tri 4999 -5458 5302 -5155 ne
rect 5302 -5458 5463 -5155
tri 5463 -5458 5766 -5155 sw
tri 5302 -5593 5437 -5458 ne
rect 4985 -5756 5273 -5751
rect 4985 -5812 4990 -5756
rect 5046 -5812 5101 -5756
rect 5157 -5812 5212 -5756
rect 5268 -5812 5273 -5756
rect 4985 -5840 5273 -5812
rect 4985 -5896 4990 -5840
rect 5046 -5896 5101 -5840
rect 5157 -5896 5212 -5840
rect 5268 -5896 5273 -5840
rect 4985 -5924 5273 -5896
rect 4985 -5980 4990 -5924
rect 5046 -5980 5101 -5924
rect 5157 -5980 5212 -5924
rect 5268 -5980 5273 -5924
rect 5437 -5773 5766 -5458
rect 5437 -5829 5442 -5773
rect 5498 -5829 5530 -5773
rect 5586 -5829 5618 -5773
rect 5674 -5829 5705 -5773
rect 5761 -5829 5766 -5773
rect 5437 -5897 5766 -5829
rect 5437 -5953 5442 -5897
rect 5498 -5953 5530 -5897
rect 5586 -5953 5618 -5897
rect 5674 -5953 5705 -5897
rect 5761 -5953 5766 -5897
rect 5437 -5958 5766 -5953
tri 6398 -5958 6430 -5926 se
rect 6430 -5958 6468 -5926
rect 4985 -6134 5273 -5980
tri 6371 -5985 6398 -5958 se
rect 6398 -5985 6468 -5958
tri 6274 -6082 6371 -5985 se
rect 6371 -6082 6468 -5985
tri 5273 -6134 5325 -6082 sw
tri 6222 -6134 6274 -6082 se
rect 6274 -6134 6468 -6082
rect 4985 -6200 6468 -6134
tri 4985 -6277 5062 -6200 ne
rect 5062 -6277 6468 -6200
tri 3237 -6314 3274 -6277 sw
tri 5062 -6314 5099 -6277 ne
rect 5099 -6314 6468 -6277
tri 5099 -6380 5165 -6314 ne
rect 5165 -6380 6468 -6314
tri 5165 -6383 5168 -6380 ne
rect 5168 -6383 6468 -6380
tri 5168 -6422 5207 -6383 ne
rect 5207 -6422 6468 -6383
tri 6228 -6439 6245 -6422 ne
rect 6245 -6439 6468 -6422
tri 6245 -6474 6280 -6439 ne
rect 6280 -6474 6468 -6439
rect 6610 -6383 6998 -4598
rect 12481 -4885 12938 -197
rect 12481 -4941 12494 -4885
rect 12550 -4941 12617 -4885
rect 12673 -4941 12740 -4885
rect 12796 -4941 12862 -4885
rect 12918 -4941 12938 -4885
rect 12481 -4989 12938 -4941
rect 12481 -5045 12494 -4989
rect 12550 -5045 12617 -4989
rect 12673 -5045 12740 -4989
rect 12796 -5045 12862 -4989
rect 12918 -5045 12938 -4989
rect 12481 -5093 12938 -5045
rect 8118 -5099 8377 -5094
rect 8118 -5155 8123 -5099
rect 8179 -5155 8220 -5099
rect 8276 -5155 8316 -5099
rect 8372 -5155 8377 -5099
rect 12481 -5149 12494 -5093
rect 12550 -5149 12617 -5093
rect 12673 -5149 12740 -5093
rect 12796 -5149 12862 -5093
rect 12918 -5149 12938 -5093
rect 12481 -5155 12938 -5149
rect 8118 -5175 8377 -5155
tri 8118 -5250 8193 -5175 ne
rect 8193 -5785 8309 -5175
tri 8309 -5243 8377 -5175 nw
rect 8193 -5841 8223 -5785
rect 8279 -5841 8309 -5785
rect 8193 -5865 8309 -5841
rect 8193 -5921 8223 -5865
rect 8279 -5921 8309 -5865
rect 8193 -5926 8309 -5921
rect 6610 -6439 6615 -6383
rect 6671 -6439 6696 -6383
rect 6752 -6439 6777 -6383
rect 6833 -6439 6857 -6383
rect 6913 -6439 6937 -6383
rect 6993 -6439 6998 -6383
rect 6610 -6474 6998 -6439
tri 6280 -6624 6430 -6474 ne
rect 6430 -6624 6468 -6474
<< via3 >>
rect 17306 21639 17311 21703
rect 17311 21639 17370 21703
rect 17388 21639 17447 21703
rect 17447 21639 17452 21703
rect 17306 21575 17311 21603
rect 17311 21575 17370 21603
rect 17388 21575 17447 21603
rect 17447 21575 17452 21603
rect 17306 21539 17370 21575
rect 17388 21539 17452 21575
rect 17306 21439 17370 21503
rect 17388 21439 17452 21503
rect 17306 21339 17370 21403
rect 17388 21339 17452 21403
rect 17306 21239 17370 21303
rect 17388 21239 17452 21303
rect 23036 10240 23100 10304
rect 23118 10240 23182 10304
rect 23036 10158 23100 10222
rect 23118 10158 23182 10222
rect 23036 10075 23100 10139
rect 23118 10075 23182 10139
rect 23036 9992 23100 10056
rect 23118 9992 23182 10056
rect 23036 9909 23100 9973
rect 23118 9909 23182 9973
rect 23036 9826 23100 9890
rect 23118 9826 23182 9890
rect 23036 9743 23100 9807
rect 23118 9743 23182 9807
rect 23036 9660 23100 9724
rect 23118 9660 23182 9724
rect 23036 9577 23100 9641
rect 23118 9577 23182 9641
<< metal4 >>
rect 5832 23936 6724 24872
rect 17305 21703 22189 21704
rect 17305 21639 17306 21703
rect 17370 21639 17388 21703
rect 17452 21639 22189 21703
rect 17305 21603 22189 21639
rect 17305 21539 17306 21603
rect 17370 21539 17388 21603
rect 17452 21539 22189 21603
rect 17305 21503 22189 21539
rect 17305 21439 17306 21503
rect 17370 21439 17388 21503
rect 17452 21439 22189 21503
rect 17305 21403 22189 21439
rect 17305 21339 17306 21403
rect 17370 21339 17388 21403
rect 17452 21339 22189 21403
rect 17305 21303 22189 21339
rect 17305 21239 17306 21303
rect 17370 21239 17388 21303
rect 17452 21242 22189 21303
tri 22189 21242 22651 21704 sw
rect 17452 21239 22651 21242
rect 17305 21238 22651 21239
tri 21772 20507 22503 21238 ne
rect 22503 10993 22651 21238
tri 22503 10943 22553 10993 ne
rect 22553 10943 22651 10993
tri 22651 10943 22763 11055 sw
tri 22553 10845 22651 10943 ne
rect 22651 10845 22763 10943
tri 22651 10733 22763 10845 ne
tri 22763 10733 22973 10943 sw
tri 22763 10523 22973 10733 ne
tri 22973 10523 23183 10733 sw
tri 22973 10465 23031 10523 ne
rect 23031 10304 23183 10523
rect 23031 10240 23036 10304
rect 23100 10240 23118 10304
rect 23182 10240 23183 10304
rect 23031 10222 23183 10240
rect 23031 10158 23036 10222
rect 23100 10158 23118 10222
rect 23182 10158 23183 10222
rect 23031 10139 23183 10158
rect 23031 10075 23036 10139
rect 23100 10075 23118 10139
rect 23182 10075 23183 10139
rect 23031 10056 23183 10075
rect 23031 9992 23036 10056
rect 23100 9992 23118 10056
rect 23182 9992 23183 10056
rect 23031 9973 23183 9992
rect 23031 9909 23036 9973
rect 23100 9909 23118 9973
rect 23182 9909 23183 9973
rect 23031 9890 23183 9909
rect 23031 9826 23036 9890
rect 23100 9826 23118 9890
rect 23182 9826 23183 9890
rect 23031 9807 23183 9826
rect 23031 9743 23036 9807
rect 23100 9743 23118 9807
rect 23182 9743 23183 9807
rect 23031 9724 23183 9743
rect 23031 9660 23036 9724
rect 23100 9660 23118 9724
rect 23182 9660 23183 9724
rect 23031 9641 23183 9660
rect 23031 9577 23036 9641
rect 23100 9577 23118 9641
rect 23182 9577 23183 9641
rect 23031 9566 23183 9577
rect 11341 8252 11824 8755
rect 15128 3154 16231 4179
use sky130_fd_io__gpio_ovtv2_hotswap_i2c_fix_leak_fix  sky130_fd_io__gpio_ovtv2_hotswap_i2c_fix_leak_fix_0
timestamp 1666199351
transform 1 0 -151 0 1 2514
box 0 -9138 27348 17659
use sky130_fd_io__gpio_ovtv2_odrvr_sub_leak_fix  sky130_fd_io__gpio_ovtv2_odrvr_sub_leak_fix_0
timestamp 1666199351
transform 1 0 -1014 0 1 -176
box 137 -2507 28211 26296
use sky130_fd_pr__nfet_01v8__example_55959141808182  sky130_fd_pr__nfet_01v8__example_55959141808182_0
timestamp 1666199351
transform -1 0 17063 0 -1 21559
box -1 0 1601 1
use sky130_fd_pr__nfet_01v8__example_55959141808182  sky130_fd_pr__nfet_01v8__example_55959141808182_1
timestamp 1666199351
transform -1 0 17063 0 -1 21357
box -1 0 1601 1
use sky130_fd_pr__nfet_01v8__example_55959141808182  sky130_fd_pr__nfet_01v8__example_55959141808182_2
timestamp 1666199351
transform -1 0 17063 0 -1 23327
box -1 0 1601 1
use sky130_fd_pr__nfet_01v8__example_55959141808182  sky130_fd_pr__nfet_01v8__example_55959141808182_3
timestamp 1666199351
transform -1 0 17063 0 -1 22603
box -1 0 1601 1
use sky130_fd_pr__nfet_01v8__example_55959141808182  sky130_fd_pr__nfet_01v8__example_55959141808182_4
timestamp 1666199351
transform -1 0 17063 0 -1 22443
box -1 0 1601 1
use sky130_fd_pr__nfet_01v8__example_55959141808182  sky130_fd_pr__nfet_01v8__example_55959141808182_5
timestamp 1666199351
transform -1 0 17063 0 -1 23125
box -1 0 1601 1
use sky130_fd_pr__nfet_01v8__example_55959141808182  sky130_fd_pr__nfet_01v8__example_55959141808182_6
timestamp 1666199351
transform -1 0 17063 0 -1 22965
box -1 0 1601 1
use sky130_fd_pr__nfet_01v8__example_55959141808182  sky130_fd_pr__nfet_01v8__example_55959141808182_7
timestamp 1666199351
transform -1 0 17063 0 -1 22763
box -1 0 1601 1
use sky130_fd_pr__nfet_01v8__example_55959141808182  sky130_fd_pr__nfet_01v8__example_55959141808182_8
timestamp 1666199351
transform -1 0 17063 0 -1 21719
box -1 0 1601 1
use sky130_fd_pr__nfet_01v8__example_55959141808182  sky130_fd_pr__nfet_01v8__example_55959141808182_9
timestamp 1666199351
transform -1 0 17063 0 -1 21921
box -1 0 1601 1
use sky130_fd_pr__nfet_01v8__example_55959141808182  sky130_fd_pr__nfet_01v8__example_55959141808182_10
timestamp 1666199351
transform -1 0 17063 0 -1 22081
box -1 0 1601 1
use sky130_fd_pr__nfet_01v8__example_55959141808182  sky130_fd_pr__nfet_01v8__example_55959141808182_11
timestamp 1666199351
transform -1 0 17063 0 -1 22241
box -1 0 1601 1
<< labels >>
flabel metal3 s 17095 21879 17134 21939 3 FreeSans 520 90 0 0 NGB_PAD_VPMP_H
port 1 nsew
flabel metal3 s 16949 21884 16994 21944 3 FreeSans 520 90 0 0 NGA_PAD_VPMP_H
port 2 nsew
flabel metal4 s 15128 3154 16231 4179 3 FreeSans 200 0 0 0 VDDIO
port 3 nsew
flabel metal4 s 5832 23936 6724 24872 3 FreeSans 600 0 0 0 VSSIO
port 4 nsew
flabel metal4 s 11341 8252 11824 8755 3 FreeSans 600 0 0 0 PAD
port 5 nsew
flabel metal2 s 1853 3279 1880 3306 0 FreeSans 200 90 0 0 NGHS_H
port 6 nsew
flabel metal2 s 17308 20844 17377 20896 3 FreeSans 200 0 0 0 PD_H[2]
port 7 nsew
flabel metal2 s 17306 20177 17391 20255 3 FreeSans 200 0 0 0 PD_H[3]
port 8 nsew
flabel metal2 s 1523 5869 1575 5947 3 FreeSans 200 0 0 0 PU_CSD_H
port 9 nsew
flabel metal2 s 1799 7756 1851 7790 3 FreeSans 200 0 0 0 PU_H_N[0]
port 10 nsew
flabel metal2 s 1891 7803 1943 7841 3 FreeSans 200 0 0 0 PU_H_N[1]
port 11 nsew
flabel metal2 s 1799 6793 1851 6848 3 FreeSans 200 0 0 0 PU_H_N[2]
port 12 nsew
flabel metal2 s 2075 6895 2127 6945 3 FreeSans 200 0 0 0 PU_H_N[3]
port 13 nsew
flabel metal2 s 2520 7745 2572 7785 3 FreeSans 200 0 0 0 PGHS_H
port 14 nsew
flabel metal2 s 17310 21315 17377 21367 3 FreeSans 200 0 0 0 PD_H[0]
port 15 nsew
flabel metal2 s 17310 21235 17378 21275 3 FreeSans 200 0 0 0 PD_H[1]
port 16 nsew
flabel metal1 s 970 1127 1110 1265 3 FreeSans 200 0 0 0 VSSD
port 17 nsew
flabel metal1 s 5424 11472 5526 11561 3 FreeSans 200 0 0 0 VSSIO_AMX
port 18 nsew
flabel metal1 s 24579 9329 24698 9447 3 FreeSans 200 0 0 0 TIE_HI_ESD
port 19 nsew
flabel metal1 s 17570 20507 17614 20598 3 FreeSans 200 0 0 0 TIE_LO_ESD
port 20 nsew
flabel metal1 s 9030 7637 9094 7669 3 FreeSans 200 0 0 0 PUG_H[5]
port 21 nsew
flabel metal1 s 7384 6988 7424 7020 3 FreeSans 200 0 0 0 PUG_H[6]
port 22 nsew
flabel metal1 s 9728 5453 9923 5547 3 FreeSans 200 0 0 0 VDDIO_AMX
port 23 nsew
flabel metal1 s 1370 2094 1679 2262 3 FreeSans 200 0 0 0 VPB_DRVR
port 24 nsew
flabel metal1 s 10260 -5648 10303 -5610 3 FreeSans 200 0 0 0 FORCE_H[1]
port 25 nsew
flabel metal1 s 11678 -5712 11739 -5680 3 FreeSans 200 0 0 0 OD_H
port 26 nsew
flabel metal1 s 10548 -5620 10591 -5581 3 FreeSans 200 0 0 0 OE_HS_H
port 27 nsew
flabel metal1 s 3273 20179 3398 20254 3 FreeSans 200 0 0 0 PD_CSD_H
port 28 nsew
flabel comment s 3202 -5556 3202 -5556 0 FreeSans 400 0 0 0 PADLO
<< properties >>
string GDS_END 42123658
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 42046144
<< end >>
