magic
tech sky130B
magscale 1 2
timestamp 1666199351
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 3 21 643 203
rect 28 -17 62 21
<< locali >>
rect 199 393 259 425
rect 482 393 529 493
rect 199 357 529 393
rect 24 289 419 323
rect 24 211 90 289
rect 124 215 284 255
rect 320 215 419 289
rect 487 119 529 357
rect 563 153 626 280
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 21 357 87 527
rect 121 459 343 493
rect 121 357 165 459
rect 305 427 343 459
rect 382 435 448 527
rect 21 143 453 177
rect 21 51 87 143
rect 123 17 157 109
rect 193 51 259 143
rect 305 17 339 109
rect 387 85 453 143
rect 563 314 625 527
rect 563 85 625 119
rect 387 51 625 85
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel locali s 320 215 419 289 6 A1
port 1 nsew signal input
rlabel locali s 24 211 90 289 6 A1
port 1 nsew signal input
rlabel locali s 24 289 419 323 6 A1
port 1 nsew signal input
rlabel locali s 124 215 284 255 6 A2
port 2 nsew signal input
rlabel locali s 563 153 626 280 6 B1
port 3 nsew signal input
rlabel metal1 s 0 -48 644 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 28 -17 62 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 3 21 643 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 682 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 644 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 487 119 529 357 6 Y
port 8 nsew signal output
rlabel locali s 199 357 529 393 6 Y
port 8 nsew signal output
rlabel locali s 482 393 529 493 6 Y
port 8 nsew signal output
rlabel locali s 199 393 259 425 6 Y
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 644 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1313876
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1307432
<< end >>
