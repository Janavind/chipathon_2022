magic
tech sky130B
magscale 1 2
timestamp 1666464484
<< nwell >>
rect -38 261 498 582
<< pwell >>
rect 1 67 368 203
rect 30 21 368 67
rect 30 -17 64 21
<< locali >>
rect 200 401 266 493
rect 200 367 434 401
rect 18 215 88 263
rect 122 215 217 263
rect 360 109 434 367
rect 284 51 434 109
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 116 367 166 527
rect 300 435 343 527
rect 18 333 74 365
rect 18 299 285 333
rect 251 265 285 299
rect 251 215 326 265
rect 251 181 285 215
rect 18 147 285 181
rect 18 105 72 147
rect 116 17 182 109
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
rlabel locali s 18 215 88 263 6 A_N
port 1 nsew signal input
rlabel locali s 122 215 217 263 6 B
port 2 nsew signal input
rlabel metal1 s 0 -48 460 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 30 21 368 67 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 1 67 368 203 6 VNB
port 4 nsew ground bidirectional
rlabel nwell s -38 261 498 582 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 496 460 592 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 284 51 434 109 6 Y
port 7 nsew signal output
rlabel locali s 360 109 434 367 6 Y
port 7 nsew signal output
rlabel locali s 200 367 434 401 6 Y
port 7 nsew signal output
rlabel locali s 200 401 266 493 6 Y
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 460 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1804548
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1800018
<< end >>
