magic
tech sky130A
magscale 1 2
timestamp 1666464484
<< nwell >>
rect -54 284 852 454
rect -59 116 857 284
rect -54 -54 852 116
<< scpmos >>
rect 60 0 90 400
rect 168 0 198 400
rect 276 0 306 400
rect 384 0 414 400
rect 492 0 522 400
rect 600 0 630 400
rect 708 0 738 400
<< pdiff >>
rect 0 217 60 400
rect 0 183 8 217
rect 42 183 60 217
rect 0 0 60 183
rect 90 217 168 400
rect 90 183 112 217
rect 146 183 168 217
rect 90 0 168 183
rect 198 217 276 400
rect 198 183 220 217
rect 254 183 276 217
rect 198 0 276 183
rect 306 217 384 400
rect 306 183 328 217
rect 362 183 384 217
rect 306 0 384 183
rect 414 217 492 400
rect 414 183 436 217
rect 470 183 492 217
rect 414 0 492 183
rect 522 217 600 400
rect 522 183 544 217
rect 578 183 600 217
rect 522 0 600 183
rect 630 217 708 400
rect 630 183 652 217
rect 686 183 708 217
rect 630 0 708 183
rect 738 217 798 400
rect 738 183 756 217
rect 790 183 798 217
rect 738 0 798 183
<< pdiffc >>
rect 8 183 42 217
rect 112 183 146 217
rect 220 183 254 217
rect 328 183 362 217
rect 436 183 470 217
rect 544 183 578 217
rect 652 183 686 217
rect 756 183 790 217
<< poly >>
rect 60 400 90 426
rect 168 400 198 426
rect 276 400 306 426
rect 384 400 414 426
rect 492 400 522 426
rect 600 400 630 426
rect 708 400 738 426
rect 60 -26 90 0
rect 168 -26 198 0
rect 276 -26 306 0
rect 384 -26 414 0
rect 492 -26 522 0
rect 600 -26 630 0
rect 708 -26 738 0
rect 60 -56 738 -26
<< locali >>
rect 8 217 42 233
rect 8 167 42 183
rect 112 217 146 233
rect 112 133 146 183
rect 220 217 254 233
rect 220 167 254 183
rect 328 217 362 233
rect 328 133 362 183
rect 436 217 470 233
rect 436 167 470 183
rect 544 217 578 233
rect 544 133 578 183
rect 652 217 686 233
rect 652 167 686 183
rect 756 217 790 233
rect 756 133 790 183
rect 112 99 790 133
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_0
timestamp 1666464484
transform 1 0 748 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_1
timestamp 1666464484
transform 1 0 644 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_2
timestamp 1666464484
transform 1 0 536 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_3
timestamp 1666464484
transform 1 0 428 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_4
timestamp 1666464484
transform 1 0 320 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_5
timestamp 1666464484
transform 1 0 212 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_6
timestamp 1666464484
transform 1 0 104 0 1 167
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_12  sky130_sram_2kbyte_1rw1r_32x512_8_contact_12_7
timestamp 1666464484
transform 1 0 0 0 1 167
box 0 0 1 1
<< labels >>
rlabel locali s 25 200 25 200 4 S
port 1 nsew
rlabel locali s 237 200 237 200 4 S
port 1 nsew
rlabel locali s 669 200 669 200 4 S
port 1 nsew
rlabel locali s 453 200 453 200 4 S
port 1 nsew
rlabel locali s 451 116 451 116 4 D
port 2 nsew
rlabel poly s 399 -41 399 -41 4 G
port 3 nsew
<< properties >>
string FIXED_BBOX -54 -56 852 116
string GDS_END 51848
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_2kbyte_1rw1r_32x512_8.gds
string GDS_START 49580
<< end >>
