magic
tech sky130B
magscale 1 2
timestamp 1666464484
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 107 157 618 203
rect 1 21 827 157
rect 30 -17 64 21
<< scnmos >>
rect 81 47 111 131
rect 183 47 283 177
rect 442 47 542 177
rect 608 47 638 131
rect 693 47 723 131
<< scpmoshvt >>
rect 81 297 111 497
rect 183 333 283 497
rect 442 333 542 497
rect 608 297 638 497
rect 693 297 723 497
<< ndiff >>
rect 133 131 183 177
rect 27 111 81 131
rect 27 77 36 111
rect 70 77 81 111
rect 27 47 81 77
rect 111 102 183 131
rect 111 68 133 102
rect 167 68 183 102
rect 111 47 183 68
rect 283 104 336 177
rect 283 70 294 104
rect 328 70 336 104
rect 283 47 336 70
rect 390 111 442 177
rect 390 77 398 111
rect 432 77 442 111
rect 390 47 442 77
rect 542 131 592 177
rect 542 97 608 131
rect 542 63 553 97
rect 587 63 608 97
rect 542 47 608 63
rect 638 111 693 131
rect 638 77 649 111
rect 683 77 693 111
rect 638 47 693 77
rect 723 111 801 131
rect 723 77 759 111
rect 793 77 801 111
rect 723 47 801 77
<< pdiff >>
rect 27 478 81 497
rect 27 444 36 478
rect 70 444 81 478
rect 27 410 81 444
rect 27 376 36 410
rect 70 376 81 410
rect 27 297 81 376
rect 111 478 183 497
rect 111 444 136 478
rect 170 444 183 478
rect 111 410 183 444
rect 111 376 136 410
rect 170 376 183 410
rect 111 333 183 376
rect 283 478 336 497
rect 283 444 294 478
rect 328 444 336 478
rect 283 410 336 444
rect 283 376 294 410
rect 328 376 336 410
rect 283 333 336 376
rect 390 477 442 497
rect 390 443 398 477
rect 432 443 442 477
rect 390 409 442 443
rect 390 375 398 409
rect 432 375 442 409
rect 390 333 442 375
rect 542 478 608 497
rect 542 444 553 478
rect 587 444 608 478
rect 542 410 608 444
rect 542 376 553 410
rect 587 376 608 410
rect 542 333 608 376
rect 111 297 161 333
rect 558 297 608 333
rect 638 477 693 497
rect 638 443 649 477
rect 683 443 693 477
rect 638 409 693 443
rect 638 375 649 409
rect 683 375 693 409
rect 638 297 693 375
rect 723 478 801 497
rect 723 444 759 478
rect 793 444 801 478
rect 723 410 801 444
rect 723 376 759 410
rect 793 376 801 410
rect 723 297 801 376
<< ndiffc >>
rect 36 77 70 111
rect 133 68 167 102
rect 294 70 328 104
rect 398 77 432 111
rect 553 63 587 97
rect 649 77 683 111
rect 759 77 793 111
<< pdiffc >>
rect 36 444 70 478
rect 36 376 70 410
rect 136 444 170 478
rect 136 376 170 410
rect 294 444 328 478
rect 294 376 328 410
rect 398 443 432 477
rect 398 375 432 409
rect 553 444 587 478
rect 553 376 587 410
rect 649 443 683 477
rect 649 375 683 409
rect 759 444 793 478
rect 759 376 793 410
<< poly >>
rect 81 497 111 523
rect 183 497 283 523
rect 442 497 542 523
rect 608 497 638 523
rect 693 497 723 523
rect 81 261 111 297
rect 30 249 111 261
rect 183 259 283 333
rect 442 261 542 333
rect 608 265 638 297
rect 30 215 46 249
rect 80 215 111 249
rect 30 203 111 215
rect 153 249 287 259
rect 153 215 169 249
rect 203 215 237 249
rect 271 215 287 249
rect 153 205 287 215
rect 395 249 542 261
rect 395 215 411 249
rect 445 215 542 249
rect 81 131 111 203
rect 183 177 283 205
rect 395 203 542 215
rect 442 177 542 203
rect 584 259 638 265
rect 693 259 723 297
rect 584 249 723 259
rect 584 215 594 249
rect 628 215 723 249
rect 584 205 723 215
rect 584 199 638 205
rect 608 131 638 199
rect 693 131 723 205
rect 81 21 111 47
rect 183 21 283 47
rect 442 21 542 47
rect 608 21 638 47
rect 693 21 723 47
<< polycont >>
rect 46 215 80 249
rect 169 215 203 249
rect 237 215 271 249
rect 411 215 445 249
rect 594 215 628 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 17 478 86 493
rect 17 444 36 478
rect 70 444 86 478
rect 17 410 86 444
rect 17 376 36 410
rect 70 376 86 410
rect 17 326 86 376
rect 120 478 186 527
rect 120 444 136 478
rect 170 444 186 478
rect 120 410 186 444
rect 120 376 136 410
rect 170 376 186 410
rect 120 360 186 376
rect 278 478 359 493
rect 278 444 294 478
rect 328 444 359 478
rect 278 410 359 444
rect 278 376 294 410
rect 328 376 359 410
rect 278 357 359 376
rect 17 291 254 326
rect 17 249 96 257
rect 170 249 254 291
rect 325 249 359 357
rect 397 477 447 493
rect 397 443 398 477
rect 432 443 447 477
rect 397 409 447 443
rect 397 375 398 409
rect 432 375 447 409
rect 397 326 447 375
rect 537 478 603 527
rect 537 444 553 478
rect 587 444 603 478
rect 537 410 603 444
rect 537 376 553 410
rect 587 376 603 410
rect 537 360 603 376
rect 637 477 725 493
rect 637 443 649 477
rect 683 443 725 477
rect 637 409 725 443
rect 637 375 649 409
rect 683 375 725 409
rect 397 292 529 326
rect 637 306 725 375
rect 759 478 811 527
rect 793 444 811 478
rect 759 410 811 444
rect 793 376 811 410
rect 759 360 811 376
rect 495 265 529 292
rect 495 249 635 265
rect 17 215 46 249
rect 80 215 96 249
rect 153 215 169 249
rect 203 215 237 249
rect 271 215 287 249
rect 325 215 411 249
rect 445 215 461 249
rect 495 215 594 249
rect 628 215 635 249
rect 170 181 254 215
rect 17 147 254 181
rect 325 180 359 215
rect 495 199 635 215
rect 495 181 529 199
rect 17 111 83 147
rect 17 77 36 111
rect 70 77 83 111
rect 17 54 83 77
rect 117 102 183 113
rect 117 68 133 102
rect 167 68 183 102
rect 117 17 183 68
rect 288 104 359 180
rect 288 70 294 104
rect 328 70 359 104
rect 288 54 359 70
rect 397 147 529 181
rect 397 111 447 147
rect 669 128 725 306
rect 397 77 398 111
rect 432 77 447 111
rect 397 54 447 77
rect 537 97 603 113
rect 537 63 553 97
rect 587 63 603 97
rect 537 17 603 63
rect 637 111 725 128
rect 637 77 649 111
rect 683 77 725 111
rect 637 54 725 77
rect 759 111 811 127
rect 793 77 811 111
rect 759 17 811 77
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
flabel locali s 30 221 64 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 678 425 712 459 0 FreeSans 400 0 0 0 X
port 6 nsew signal output
flabel locali s 678 357 712 391 0 FreeSans 400 0 0 0 X
port 6 nsew signal output
flabel locali s 678 289 712 323 0 FreeSans 400 0 0 0 X
port 6 nsew signal output
flabel locali s 678 221 712 255 0 FreeSans 400 0 0 0 X
port 6 nsew signal output
flabel locali s 678 153 712 187 0 FreeSans 400 0 0 0 X
port 6 nsew signal output
flabel locali s 678 85 712 119 0 FreeSans 400 0 0 0 X
port 6 nsew signal output
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 clkdlybuf4s50_2
rlabel metal1 s 0 -48 828 48 1 VGND
port 2 nsew ground bidirectional abutment
rlabel metal1 s 0 496 828 592 1 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 828 544
string GDS_END 3303806
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3297206
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 20.700 0.000 
<< end >>
