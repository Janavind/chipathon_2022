magic
tech sky130A
magscale 1 2
timestamp 1666199351
use sky130_fd_pr__dfl1sd2__example_55959141808191  sky130_fd_pr__dfl1sd2__example_55959141808191_0
timestamp 1666199351
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808191  sky130_fd_pr__dfl1sd2__example_55959141808191_1
timestamp 1666199351
transform 1 0 256 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808191  sky130_fd_pr__dfl1sd2__example_55959141808191_2
timestamp 1666199351
transform 1 0 412 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808191  sky130_fd_pr__dfl1sd2__example_55959141808191_3
timestamp 1666199351
transform 1 0 568 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_55959141808190  sky130_fd_pr__dfl1sd__example_55959141808190_0
timestamp 1666199351
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_55959141808190  sky130_fd_pr__dfl1sd__example_55959141808190_1
timestamp 1666199351
transform 1 0 724 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 42328024
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 42324910
<< end >>
