// This is the unpowered netlist.
module macro_2to3 (io_active,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input io_active;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [127:0] la_data_in;
 output [127:0] la_data_out;
 input [127:0] la_oenb;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire active;

 sky130_fd_sc_hd__inv_2 _170_ (.A(active),
    .Y(_137_));
 sky130_fd_sc_hd__buf_1 _171_ (.A(active),
    .X(_099_));
 sky130_fd_sc_hd__buf_1 _172_ (.A(_099_),
    .X(_100_));
 sky130_fd_sc_hd__buf_1 _173_ (.A(_100_),
    .X(_101_));
 sky130_fd_sc_hd__inv_2 _174_ (.A(_101_),
    .Y(_136_));
 sky130_fd_sc_hd__inv_2 _175_ (.A(_101_),
    .Y(_135_));
 sky130_fd_sc_hd__inv_2 _176_ (.A(_101_),
    .Y(_134_));
 sky130_fd_sc_hd__inv_2 _177_ (.A(_101_),
    .Y(_133_));
 sky130_fd_sc_hd__inv_2 _178_ (.A(_101_),
    .Y(_132_));
 sky130_fd_sc_hd__buf_1 _179_ (.A(_100_),
    .X(_102_));
 sky130_fd_sc_hd__inv_2 _180_ (.A(_102_),
    .Y(_131_));
 sky130_fd_sc_hd__inv_2 _181_ (.A(_102_),
    .Y(_130_));
 sky130_fd_sc_hd__inv_2 _182_ (.A(_102_),
    .Y(_129_));
 sky130_fd_sc_hd__inv_2 _183_ (.A(_102_),
    .Y(_128_));
 sky130_fd_sc_hd__inv_2 _184_ (.A(_102_),
    .Y(_127_));
 sky130_fd_sc_hd__buf_1 _185_ (.A(_100_),
    .X(_103_));
 sky130_fd_sc_hd__inv_2 _186_ (.A(_103_),
    .Y(_126_));
 sky130_fd_sc_hd__inv_2 _187_ (.A(_103_),
    .Y(_125_));
 sky130_fd_sc_hd__inv_2 _188_ (.A(_103_),
    .Y(_124_));
 sky130_fd_sc_hd__inv_2 _189_ (.A(_103_),
    .Y(_123_));
 sky130_fd_sc_hd__inv_2 _190_ (.A(_103_),
    .Y(_122_));
 sky130_fd_sc_hd__buf_1 _191_ (.A(_100_),
    .X(_104_));
 sky130_fd_sc_hd__inv_2 _192_ (.A(_104_),
    .Y(_121_));
 sky130_fd_sc_hd__inv_2 _193_ (.A(_104_),
    .Y(_120_));
 sky130_fd_sc_hd__inv_2 _194_ (.A(_104_),
    .Y(_119_));
 sky130_fd_sc_hd__inv_2 _195_ (.A(_104_),
    .Y(_118_));
 sky130_fd_sc_hd__inv_2 _196_ (.A(_104_),
    .Y(_117_));
 sky130_fd_sc_hd__buf_1 _197_ (.A(_099_),
    .X(_105_));
 sky130_fd_sc_hd__inv_2 _198_ (.A(_105_),
    .Y(_116_));
 sky130_fd_sc_hd__inv_2 _199_ (.A(_105_),
    .Y(_115_));
 sky130_fd_sc_hd__inv_2 _200_ (.A(_105_),
    .Y(_114_));
 sky130_fd_sc_hd__inv_2 _201_ (.A(_105_),
    .Y(_113_));
 sky130_fd_sc_hd__inv_2 _202_ (.A(_105_),
    .Y(_112_));
 sky130_fd_sc_hd__buf_1 _203_ (.A(_099_),
    .X(_000_));
 sky130_fd_sc_hd__inv_2 _204_ (.A(_000_),
    .Y(_111_));
 sky130_fd_sc_hd__inv_2 _205_ (.A(_000_),
    .Y(_110_));
 sky130_fd_sc_hd__inv_2 _206_ (.A(_000_),
    .Y(_109_));
 sky130_fd_sc_hd__inv_2 _207_ (.A(_000_),
    .Y(_108_));
 sky130_fd_sc_hd__inv_2 _208_ (.A(_000_),
    .Y(_107_));
 sky130_fd_sc_hd__inv_2 _209_ (.A(_100_),
    .Y(_106_));
 sky130_fd_sc_hd__buf_1 _210_ (.A(io_in[23]),
    .X(_001_));
 sky130_fd_sc_hd__nand3b_2 _211_ (.A_N(io_in[35]),
    .B(io_in[34]),
    .C(io_in[35]),
    .Y(_002_));
 sky130_fd_sc_hd__o31a_2 _212_ (.A1(io_in[24]),
    .A2(io_in[22]),
    .A3(_001_),
    .B1(_002_),
    .X(_003_));
 sky130_fd_sc_hd__xnor3_2 _213_ (.A(io_in[25]),
    .B(_003_),
    .C(io_in[25]),
    .X(_004_));
 sky130_fd_sc_hd__or3_2 _214_ (.A(io_in[21]),
    .B(_004_),
    .C(io_in[21]),
    .X(_005_));
 sky130_fd_sc_hd__o21a_2 _215_ (.A1(io_in[22]),
    .A2(_001_),
    .B1(_002_),
    .X(_006_));
 sky130_fd_sc_hd__xnor3_2 _216_ (.A(io_in[24]),
    .B(_006_),
    .C(io_in[24]),
    .X(_007_));
 sky130_fd_sc_hd__or3_2 _217_ (.A(io_in[20]),
    .B(_007_),
    .C(io_in[20]),
    .X(_008_));
 sky130_fd_sc_hd__buf_1 _218_ (.A(io_in[22]),
    .X(_009_));
 sky130_fd_sc_hd__nand3b_2 _219_ (.A_N(_001_),
    .B(_002_),
    .C(_009_),
    .Y(_010_));
 sky130_fd_sc_hd__a21bo_2 _220_ (.A1(io_in[22]),
    .A2(_002_),
    .B1_N(io_in[23]),
    .X(_011_));
 sky130_fd_sc_hd__a21o_2 _221_ (.A1(_010_),
    .A2(_011_),
    .B1(io_in[19]),
    .X(_012_));
 sky130_fd_sc_hd__or3b_2 _222_ (.A(io_in[18]),
    .B(io_in[18]),
    .C_N(_009_),
    .X(_013_));
 sky130_fd_sc_hd__and3_2 _223_ (.A(io_in[19]),
    .B(_010_),
    .C(_011_),
    .X(_014_));
 sky130_fd_sc_hd__a21o_2 _224_ (.A1(_012_),
    .A2(_013_),
    .B1(_014_),
    .X(_015_));
 sky130_fd_sc_hd__and3_2 _225_ (.A(io_in[21]),
    .B(_004_),
    .C(io_in[21]),
    .X(_016_));
 sky130_fd_sc_hd__and3_2 _226_ (.A(io_in[20]),
    .B(_007_),
    .C(io_in[20]),
    .X(_017_));
 sky130_fd_sc_hd__a211o_2 _227_ (.A1(_008_),
    .A2(_015_),
    .B1(_016_),
    .C1(_017_),
    .X(_018_));
 sky130_fd_sc_hd__a21oi_2 _228_ (.A1(io_in[25]),
    .A2(_002_),
    .B1(_003_),
    .Y(_019_));
 sky130_fd_sc_hd__a21oi_2 _229_ (.A1(_005_),
    .A2(_018_),
    .B1(_019_),
    .Y(_020_));
 sky130_fd_sc_hd__buf_1 _230_ (.A(io_in[35]),
    .X(_021_));
 sky130_fd_sc_hd__a31o_2 _231_ (.A1(_019_),
    .A2(_005_),
    .A3(_018_),
    .B1(_021_),
    .X(_022_));
 sky130_fd_sc_hd__or3_2 _232_ (.A(_020_),
    .B(_022_),
    .C(_020_),
    .X(_023_));
 sky130_fd_sc_hd__buf_1 _233_ (.A(io_in[31]),
    .X(_024_));
 sky130_fd_sc_hd__nand3b_2 _234_ (.A_N(io_in[37]),
    .B(io_in[36]),
    .C(io_in[37]),
    .Y(_025_));
 sky130_fd_sc_hd__o31a_2 _235_ (.A1(io_in[32]),
    .A2(io_in[30]),
    .A3(_024_),
    .B1(_025_),
    .X(_026_));
 sky130_fd_sc_hd__xnor3_2 _236_ (.A(io_in[33]),
    .B(_026_),
    .C(io_in[33]),
    .X(_027_));
 sky130_fd_sc_hd__or3_2 _237_ (.A(io_in[29]),
    .B(_027_),
    .C(io_in[29]),
    .X(_028_));
 sky130_fd_sc_hd__o21a_2 _238_ (.A1(io_in[30]),
    .A2(_024_),
    .B1(_025_),
    .X(_029_));
 sky130_fd_sc_hd__xnor3_2 _239_ (.A(io_in[32]),
    .B(_029_),
    .C(io_in[32]),
    .X(_030_));
 sky130_fd_sc_hd__or3_2 _240_ (.A(io_in[28]),
    .B(_030_),
    .C(io_in[28]),
    .X(_031_));
 sky130_fd_sc_hd__buf_1 _241_ (.A(io_in[30]),
    .X(_032_));
 sky130_fd_sc_hd__nand3b_2 _242_ (.A_N(_024_),
    .B(_025_),
    .C(_032_),
    .Y(_033_));
 sky130_fd_sc_hd__a21bo_2 _243_ (.A1(io_in[30]),
    .A2(_025_),
    .B1_N(io_in[31]),
    .X(_034_));
 sky130_fd_sc_hd__a21o_2 _244_ (.A1(_033_),
    .A2(_034_),
    .B1(io_in[27]),
    .X(_035_));
 sky130_fd_sc_hd__or3b_2 _245_ (.A(io_in[26]),
    .B(io_in[26]),
    .C_N(_032_),
    .X(_036_));
 sky130_fd_sc_hd__and3_2 _246_ (.A(io_in[27]),
    .B(_033_),
    .C(_034_),
    .X(_037_));
 sky130_fd_sc_hd__a21o_2 _247_ (.A1(_035_),
    .A2(_036_),
    .B1(_037_),
    .X(_038_));
 sky130_fd_sc_hd__and3_2 _248_ (.A(io_in[29]),
    .B(_027_),
    .C(io_in[29]),
    .X(_039_));
 sky130_fd_sc_hd__and3_2 _249_ (.A(io_in[28]),
    .B(_030_),
    .C(io_in[28]),
    .X(_040_));
 sky130_fd_sc_hd__a211o_2 _250_ (.A1(_031_),
    .A2(_038_),
    .B1(_039_),
    .C1(_040_),
    .X(_041_));
 sky130_fd_sc_hd__a21oi_2 _251_ (.A1(io_in[33]),
    .A2(_025_),
    .B1(_026_),
    .Y(_042_));
 sky130_fd_sc_hd__a21oi_2 _252_ (.A1(_028_),
    .A2(_041_),
    .B1(_042_),
    .Y(_043_));
 sky130_fd_sc_hd__buf_1 _253_ (.A(io_in[37]),
    .X(_044_));
 sky130_fd_sc_hd__a31o_2 _254_ (.A1(_042_),
    .A2(_028_),
    .A3(_041_),
    .B1(_044_),
    .X(_045_));
 sky130_fd_sc_hd__or3_2 _255_ (.A(_043_),
    .B(_045_),
    .C(_043_),
    .X(_046_));
 sky130_fd_sc_hd__nor3_2 _256_ (.A(_137_),
    .B(_043_),
    .C(_045_),
    .Y(io_out[4]));
 sky130_fd_sc_hd__nor3_2 _257_ (.A(_137_),
    .B(_020_),
    .C(_022_),
    .Y(io_out[5]));
 sky130_fd_sc_hd__o22a_2 _258_ (.A1(_023_),
    .A2(_046_),
    .B1(io_out[4]),
    .B2(io_out[5]),
    .X(io_out[0]));
 sky130_fd_sc_hd__inv_2 _259_ (.A(io_in[35]),
    .Y(_047_));
 sky130_fd_sc_hd__o2bb2a_2 _260_ (.A1_N(_009_),
    .A2_N(io_in[18]),
    .B1(_047_),
    .B2(io_in[34]),
    .X(_048_));
 sky130_fd_sc_hd__o21a_2 _261_ (.A1(_009_),
    .A2(io_in[18]),
    .B1(_048_),
    .X(_049_));
 sky130_fd_sc_hd__a31o_2 _262_ (.A1(_009_),
    .A2(_021_),
    .A3(io_in[18]),
    .B1(_049_),
    .X(_050_));
 sky130_fd_sc_hd__inv_2 _263_ (.A(io_in[37]),
    .Y(_051_));
 sky130_fd_sc_hd__o2bb2a_2 _264_ (.A1_N(_032_),
    .A2_N(io_in[26]),
    .B1(_051_),
    .B2(io_in[36]),
    .X(_052_));
 sky130_fd_sc_hd__o21a_2 _265_ (.A1(_032_),
    .A2(io_in[26]),
    .B1(_052_),
    .X(_053_));
 sky130_fd_sc_hd__a31o_2 _266_ (.A1(_032_),
    .A2(_044_),
    .A3(io_in[26]),
    .B1(_053_),
    .X(_054_));
 sky130_fd_sc_hd__buf_1 _267_ (.A(active),
    .X(_055_));
 sky130_fd_sc_hd__and3_2 _268_ (.A(_055_),
    .B(_054_),
    .C(_055_),
    .X(_056_));
 sky130_fd_sc_hd__buf_1 _269_ (.A(_056_),
    .X(io_out[10]));
 sky130_fd_sc_hd__and3_2 _270_ (.A(_099_),
    .B(_050_),
    .C(_099_),
    .X(_057_));
 sky130_fd_sc_hd__buf_1 _271_ (.A(_057_),
    .X(io_out[14]));
 sky130_fd_sc_hd__o2bb2a_2 _272_ (.A1_N(_050_),
    .A2_N(_054_),
    .B1(io_out[10]),
    .B2(io_out[14]),
    .X(io_out[6]));
 sky130_fd_sc_hd__or3b_2 _273_ (.A(_014_),
    .B(_014_),
    .C_N(_012_),
    .X(_058_));
 sky130_fd_sc_hd__xnor3_2 _274_ (.A(_058_),
    .B(_013_),
    .C(_058_),
    .X(_059_));
 sky130_fd_sc_hd__buf_1 _275_ (.A(io_in[34]),
    .X(_060_));
 sky130_fd_sc_hd__o21a_2 _276_ (.A1(_001_),
    .A2(io_in[34]),
    .B1(io_in[19]),
    .X(_061_));
 sky130_fd_sc_hd__a211o_2 _277_ (.A1(_001_),
    .A2(_060_),
    .B1(_047_),
    .C1(_061_),
    .X(_062_));
 sky130_fd_sc_hd__o21a_2 _278_ (.A1(_021_),
    .A2(_059_),
    .B1(_062_),
    .X(_063_));
 sky130_fd_sc_hd__or3b_2 _279_ (.A(_037_),
    .B(_037_),
    .C_N(_035_),
    .X(_064_));
 sky130_fd_sc_hd__xnor3_2 _280_ (.A(_064_),
    .B(_036_),
    .C(_064_),
    .X(_065_));
 sky130_fd_sc_hd__buf_1 _281_ (.A(io_in[36]),
    .X(_066_));
 sky130_fd_sc_hd__o21a_2 _282_ (.A1(_024_),
    .A2(io_in[36]),
    .B1(io_in[27]),
    .X(_067_));
 sky130_fd_sc_hd__a211o_2 _283_ (.A1(_024_),
    .A2(_066_),
    .B1(_051_),
    .C1(_067_),
    .X(_068_));
 sky130_fd_sc_hd__o21a_2 _284_ (.A1(_044_),
    .A2(_065_),
    .B1(_068_),
    .X(_069_));
 sky130_fd_sc_hd__and3_2 _285_ (.A(_055_),
    .B(_069_),
    .C(_055_),
    .X(_070_));
 sky130_fd_sc_hd__buf_1 _286_ (.A(_070_),
    .X(io_out[11]));
 sky130_fd_sc_hd__and3_2 _287_ (.A(_055_),
    .B(_063_),
    .C(_055_),
    .X(_071_));
 sky130_fd_sc_hd__buf_1 _288_ (.A(_071_),
    .X(io_out[15]));
 sky130_fd_sc_hd__o2bb2a_2 _289_ (.A1_N(_063_),
    .A2_N(_069_),
    .B1(io_out[11]),
    .B2(io_out[15]),
    .X(io_out[7]));
 sky130_fd_sc_hd__a21o_2 _290_ (.A1(_060_),
    .A2(io_in[20]),
    .B1(io_in[24]),
    .X(_072_));
 sky130_fd_sc_hd__or3_2 _291_ (.A(_060_),
    .B(io_in[20]),
    .C(_060_),
    .X(_073_));
 sky130_fd_sc_hd__xor3_2 _292_ (.A(io_in[20]),
    .B(_007_),
    .C(io_in[20]),
    .X(_074_));
 sky130_fd_sc_hd__or3_2 _293_ (.A(_074_),
    .B(_015_),
    .C(_074_),
    .X(_075_));
 sky130_fd_sc_hd__a21oi_2 _294_ (.A1(_074_),
    .A2(_015_),
    .B1(io_in[35]),
    .Y(_076_));
 sky130_fd_sc_hd__a32o_2 _295_ (.A1(io_in[35]),
    .A2(_072_),
    .A3(_073_),
    .B1(_075_),
    .B2(_076_),
    .X(_077_));
 sky130_fd_sc_hd__a21o_2 _296_ (.A1(_066_),
    .A2(io_in[28]),
    .B1(io_in[32]),
    .X(_078_));
 sky130_fd_sc_hd__or3_2 _297_ (.A(_066_),
    .B(io_in[28]),
    .C(_066_),
    .X(_079_));
 sky130_fd_sc_hd__xor3_2 _298_ (.A(io_in[28]),
    .B(_030_),
    .C(io_in[28]),
    .X(_080_));
 sky130_fd_sc_hd__or3_2 _299_ (.A(_080_),
    .B(_038_),
    .C(_080_),
    .X(_081_));
 sky130_fd_sc_hd__a21oi_2 _300_ (.A1(_080_),
    .A2(_038_),
    .B1(_044_),
    .Y(_082_));
 sky130_fd_sc_hd__a32o_2 _301_ (.A1(_044_),
    .A2(_078_),
    .A3(_079_),
    .B1(_081_),
    .B2(_082_),
    .X(_083_));
 sky130_fd_sc_hd__and3_2 _302_ (.A(_055_),
    .B(_083_),
    .C(_055_),
    .X(_084_));
 sky130_fd_sc_hd__buf_1 _303_ (.A(_084_),
    .X(io_out[12]));
 sky130_fd_sc_hd__and3_2 _304_ (.A(_055_),
    .B(_077_),
    .C(_055_),
    .X(_085_));
 sky130_fd_sc_hd__buf_1 _305_ (.A(_085_),
    .X(io_out[16]));
 sky130_fd_sc_hd__o2bb2a_2 _306_ (.A1_N(_077_),
    .A2_N(_083_),
    .B1(io_out[12]),
    .B2(io_out[16]),
    .X(io_out[8]));
 sky130_fd_sc_hd__a21oi_2 _307_ (.A1(_008_),
    .A2(_015_),
    .B1(_017_),
    .Y(_086_));
 sky130_fd_sc_hd__and3b_2 _308_ (.A_N(_016_),
    .B(_005_),
    .C(_016_),
    .X(_087_));
 sky130_fd_sc_hd__xnor3_2 _309_ (.A(_086_),
    .B(_087_),
    .C(_086_),
    .X(_088_));
 sky130_fd_sc_hd__nor3_2 _310_ (.A(_021_),
    .B(_088_),
    .C(_021_),
    .Y(_089_));
 sky130_fd_sc_hd__o21a_2 _311_ (.A1(io_in[25]),
    .A2(_060_),
    .B1(io_in[21]),
    .X(_090_));
 sky130_fd_sc_hd__a21o_2 _312_ (.A1(io_in[25]),
    .A2(_060_),
    .B1(_047_),
    .X(_091_));
 sky130_fd_sc_hd__nor3_2 _313_ (.A(_090_),
    .B(_091_),
    .C(_090_),
    .Y(_092_));
 sky130_fd_sc_hd__a21o_2 _314_ (.A1(_031_),
    .A2(_038_),
    .B1(_040_),
    .X(_093_));
 sky130_fd_sc_hd__and3b_2 _315_ (.A_N(_039_),
    .B(_028_),
    .C(_039_),
    .X(_094_));
 sky130_fd_sc_hd__xnor3_2 _316_ (.A(_093_),
    .B(_094_),
    .C(_093_),
    .X(_095_));
 sky130_fd_sc_hd__o21a_2 _317_ (.A1(io_in[33]),
    .A2(_066_),
    .B1(io_in[29]),
    .X(_096_));
 sky130_fd_sc_hd__a211oi_2 _318_ (.A1(io_in[33]),
    .A2(_066_),
    .B1(_051_),
    .C1(_096_),
    .Y(_097_));
 sky130_fd_sc_hd__a21o_2 _319_ (.A1(_051_),
    .A2(_095_),
    .B1(_097_),
    .X(_098_));
 sky130_fd_sc_hd__a211oi_2 _320_ (.A1(_051_),
    .A2(_095_),
    .B1(_097_),
    .C1(_137_),
    .Y(io_out[13]));
 sky130_fd_sc_hd__o221a_2 _321_ (.A1(_021_),
    .A2(_088_),
    .B1(_090_),
    .B2(_091_),
    .C1(_099_),
    .X(io_out[17]));
 sky130_fd_sc_hd__o32a_2 _322_ (.A1(_089_),
    .A2(_092_),
    .A3(_098_),
    .B1(io_out[13]),
    .B2(io_out[17]),
    .X(io_out[9]));
 sky130_fd_sc_hd__conb_1 _323_ (.LO(io_oeb[28]));
 sky130_fd_sc_hd__conb_1 _324_ (.LO(io_oeb[29]));
 sky130_fd_sc_hd__conb_1 _325_ (.LO(io_oeb[30]));
 sky130_fd_sc_hd__conb_1 _326_ (.LO(io_oeb[31]));
 sky130_fd_sc_hd__conb_1 _327_ (.LO(io_oeb[32]));
 sky130_fd_sc_hd__conb_1 _328_ (.LO(io_oeb[33]));
 sky130_fd_sc_hd__conb_1 _329_ (.LO(io_oeb[34]));
 sky130_fd_sc_hd__conb_1 _330_ (.LO(io_oeb[35]));
 sky130_fd_sc_hd__conb_1 _331_ (.LO(io_oeb[36]));
 sky130_fd_sc_hd__conb_1 _332_ (.LO(io_oeb[37]));
 sky130_fd_sc_hd__conb_1 _333_ (.LO(io_out[1]));
 sky130_fd_sc_hd__conb_1 _334_ (.LO(io_out[2]));
 sky130_fd_sc_hd__conb_1 _335_ (.LO(io_out[3]));
 sky130_fd_sc_hd__conb_1 _336_ (.LO(io_out[18]));
 sky130_fd_sc_hd__conb_1 _337_ (.LO(io_out[19]));
 sky130_fd_sc_hd__conb_1 _338_ (.LO(io_out[20]));
 sky130_fd_sc_hd__conb_1 _339_ (.LO(io_out[21]));
 sky130_fd_sc_hd__conb_1 _340_ (.LO(io_out[22]));
 sky130_fd_sc_hd__conb_1 _341_ (.LO(io_out[23]));
 sky130_fd_sc_hd__conb_1 _342_ (.LO(io_out[24]));
 sky130_fd_sc_hd__conb_1 _343_ (.LO(io_out[25]));
 sky130_fd_sc_hd__conb_1 _344_ (.LO(io_out[26]));
 sky130_fd_sc_hd__conb_1 _345_ (.LO(io_out[27]));
 sky130_fd_sc_hd__conb_1 _346_ (.LO(io_out[28]));
 sky130_fd_sc_hd__conb_1 _347_ (.LO(io_out[29]));
 sky130_fd_sc_hd__conb_1 _348_ (.LO(io_out[30]));
 sky130_fd_sc_hd__conb_1 _349_ (.LO(io_out[31]));
 sky130_fd_sc_hd__conb_1 _350_ (.LO(io_out[32]));
 sky130_fd_sc_hd__conb_1 _351_ (.LO(io_out[33]));
 sky130_fd_sc_hd__conb_1 _352_ (.LO(io_out[34]));
 sky130_fd_sc_hd__conb_1 _353_ (.LO(io_out[35]));
 sky130_fd_sc_hd__conb_1 _354_ (.LO(io_out[36]));
 sky130_fd_sc_hd__conb_1 _355_ (.LO(io_out[37]));
 sky130_fd_sc_hd__conb_1 _356_ (.LO(la_data_out[0]));
 sky130_fd_sc_hd__conb_1 _357_ (.LO(la_data_out[1]));
 sky130_fd_sc_hd__conb_1 _358_ (.LO(la_data_out[2]));
 sky130_fd_sc_hd__conb_1 _359_ (.LO(la_data_out[3]));
 sky130_fd_sc_hd__conb_1 _360_ (.LO(la_data_out[4]));
 sky130_fd_sc_hd__conb_1 _361_ (.LO(la_data_out[5]));
 sky130_fd_sc_hd__conb_1 _362_ (.LO(la_data_out[6]));
 sky130_fd_sc_hd__conb_1 _363_ (.LO(la_data_out[7]));
 sky130_fd_sc_hd__conb_1 _364_ (.LO(la_data_out[8]));
 sky130_fd_sc_hd__conb_1 _365_ (.LO(la_data_out[9]));
 sky130_fd_sc_hd__conb_1 _366_ (.LO(la_data_out[10]));
 sky130_fd_sc_hd__conb_1 _367_ (.LO(la_data_out[11]));
 sky130_fd_sc_hd__conb_1 _368_ (.LO(la_data_out[12]));
 sky130_fd_sc_hd__conb_1 _369_ (.LO(la_data_out[13]));
 sky130_fd_sc_hd__conb_1 _370_ (.LO(la_data_out[14]));
 sky130_fd_sc_hd__conb_1 _371_ (.LO(la_data_out[15]));
 sky130_fd_sc_hd__conb_1 _372_ (.LO(la_data_out[16]));
 sky130_fd_sc_hd__conb_1 _373_ (.LO(la_data_out[17]));
 sky130_fd_sc_hd__conb_1 _374_ (.LO(la_data_out[18]));
 sky130_fd_sc_hd__conb_1 _375_ (.LO(la_data_out[19]));
 sky130_fd_sc_hd__conb_1 _376_ (.LO(la_data_out[20]));
 sky130_fd_sc_hd__conb_1 _377_ (.LO(la_data_out[21]));
 sky130_fd_sc_hd__conb_1 _378_ (.LO(la_data_out[22]));
 sky130_fd_sc_hd__conb_1 _379_ (.LO(la_data_out[23]));
 sky130_fd_sc_hd__conb_1 _380_ (.LO(la_data_out[24]));
 sky130_fd_sc_hd__conb_1 _381_ (.LO(la_data_out[25]));
 sky130_fd_sc_hd__conb_1 _382_ (.LO(la_data_out[26]));
 sky130_fd_sc_hd__conb_1 _383_ (.LO(la_data_out[27]));
 sky130_fd_sc_hd__conb_1 _384_ (.LO(la_data_out[28]));
 sky130_fd_sc_hd__conb_1 _385_ (.LO(la_data_out[29]));
 sky130_fd_sc_hd__conb_1 _386_ (.LO(la_data_out[30]));
 sky130_fd_sc_hd__conb_1 _387_ (.LO(la_data_out[31]));
 sky130_fd_sc_hd__conb_1 _388_ (.LO(la_data_out[64]));
 sky130_fd_sc_hd__conb_1 _389_ (.LO(la_data_out[65]));
 sky130_fd_sc_hd__conb_1 _390_ (.LO(la_data_out[66]));
 sky130_fd_sc_hd__conb_1 _391_ (.LO(la_data_out[67]));
 sky130_fd_sc_hd__conb_1 _392_ (.LO(la_data_out[68]));
 sky130_fd_sc_hd__conb_1 _393_ (.LO(la_data_out[69]));
 sky130_fd_sc_hd__conb_1 _394_ (.LO(la_data_out[70]));
 sky130_fd_sc_hd__conb_1 _395_ (.LO(la_data_out[71]));
 sky130_fd_sc_hd__conb_1 _396_ (.LO(la_data_out[72]));
 sky130_fd_sc_hd__conb_1 _397_ (.LO(la_data_out[73]));
 sky130_fd_sc_hd__conb_1 _398_ (.LO(la_data_out[74]));
 sky130_fd_sc_hd__conb_1 _399_ (.LO(la_data_out[75]));
 sky130_fd_sc_hd__conb_1 _400_ (.LO(la_data_out[76]));
 sky130_fd_sc_hd__conb_1 _401_ (.LO(la_data_out[77]));
 sky130_fd_sc_hd__conb_1 _402_ (.LO(la_data_out[78]));
 sky130_fd_sc_hd__conb_1 _403_ (.LO(la_data_out[79]));
 sky130_fd_sc_hd__conb_1 _404_ (.LO(la_data_out[80]));
 sky130_fd_sc_hd__conb_1 _405_ (.LO(la_data_out[81]));
 sky130_fd_sc_hd__conb_1 _406_ (.LO(la_data_out[82]));
 sky130_fd_sc_hd__conb_1 _407_ (.LO(la_data_out[83]));
 sky130_fd_sc_hd__conb_1 _408_ (.LO(la_data_out[84]));
 sky130_fd_sc_hd__conb_1 _409_ (.LO(la_data_out[85]));
 sky130_fd_sc_hd__conb_1 _410_ (.LO(la_data_out[86]));
 sky130_fd_sc_hd__conb_1 _411_ (.LO(la_data_out[87]));
 sky130_fd_sc_hd__conb_1 _412_ (.LO(la_data_out[88]));
 sky130_fd_sc_hd__conb_1 _413_ (.LO(la_data_out[89]));
 sky130_fd_sc_hd__conb_1 _414_ (.LO(la_data_out[90]));
 sky130_fd_sc_hd__conb_1 _415_ (.LO(la_data_out[91]));
 sky130_fd_sc_hd__conb_1 _416_ (.LO(la_data_out[92]));
 sky130_fd_sc_hd__conb_1 _417_ (.LO(la_data_out[93]));
 sky130_fd_sc_hd__conb_1 _418_ (.LO(la_data_out[94]));
 sky130_fd_sc_hd__conb_1 _419_ (.LO(la_data_out[95]));
 sky130_fd_sc_hd__conb_1 _420_ (.LO(la_data_out[96]));
 sky130_fd_sc_hd__conb_1 _421_ (.LO(la_data_out[97]));
 sky130_fd_sc_hd__conb_1 _422_ (.LO(la_data_out[98]));
 sky130_fd_sc_hd__conb_1 _423_ (.LO(la_data_out[99]));
 sky130_fd_sc_hd__conb_1 _424_ (.LO(la_data_out[100]));
 sky130_fd_sc_hd__conb_1 _425_ (.LO(la_data_out[101]));
 sky130_fd_sc_hd__conb_1 _426_ (.LO(la_data_out[102]));
 sky130_fd_sc_hd__conb_1 _427_ (.LO(la_data_out[103]));
 sky130_fd_sc_hd__conb_1 _428_ (.LO(la_data_out[104]));
 sky130_fd_sc_hd__conb_1 _429_ (.LO(la_data_out[105]));
 sky130_fd_sc_hd__conb_1 _430_ (.LO(la_data_out[106]));
 sky130_fd_sc_hd__conb_1 _431_ (.LO(la_data_out[107]));
 sky130_fd_sc_hd__conb_1 _432_ (.LO(la_data_out[108]));
 sky130_fd_sc_hd__conb_1 _433_ (.LO(la_data_out[109]));
 sky130_fd_sc_hd__conb_1 _434_ (.LO(la_data_out[110]));
 sky130_fd_sc_hd__conb_1 _435_ (.LO(la_data_out[111]));
 sky130_fd_sc_hd__conb_1 _436_ (.LO(la_data_out[112]));
 sky130_fd_sc_hd__conb_1 _437_ (.LO(la_data_out[113]));
 sky130_fd_sc_hd__conb_1 _438_ (.LO(la_data_out[114]));
 sky130_fd_sc_hd__conb_1 _439_ (.LO(la_data_out[115]));
 sky130_fd_sc_hd__conb_1 _440_ (.LO(la_data_out[116]));
 sky130_fd_sc_hd__conb_1 _441_ (.LO(la_data_out[117]));
 sky130_fd_sc_hd__conb_1 _442_ (.LO(la_data_out[118]));
 sky130_fd_sc_hd__conb_1 _443_ (.LO(la_data_out[119]));
 sky130_fd_sc_hd__conb_1 _444_ (.LO(la_data_out[120]));
 sky130_fd_sc_hd__conb_1 _445_ (.LO(la_data_out[121]));
 sky130_fd_sc_hd__conb_1 _446_ (.LO(la_data_out[122]));
 sky130_fd_sc_hd__conb_1 _447_ (.LO(la_data_out[123]));
 sky130_fd_sc_hd__conb_1 _448_ (.LO(la_data_out[124]));
 sky130_fd_sc_hd__conb_1 _449_ (.LO(la_data_out[125]));
 sky130_fd_sc_hd__conb_1 _450_ (.LO(la_data_out[126]));
 sky130_fd_sc_hd__conb_1 _451_ (.LO(la_data_out[127]));
 sky130_fd_sc_hd__conb_1 _455_ (.LO(wbs_ack_o));
 sky130_fd_sc_hd__conb_1 _456_ (.LO(wbs_dat_o[0]));
 sky130_fd_sc_hd__conb_1 _457_ (.LO(wbs_dat_o[1]));
 sky130_fd_sc_hd__conb_1 _458_ (.LO(wbs_dat_o[2]));
 sky130_fd_sc_hd__conb_1 _459_ (.LO(wbs_dat_o[3]));
 sky130_fd_sc_hd__conb_1 _460_ (.LO(wbs_dat_o[4]));
 sky130_fd_sc_hd__conb_1 _461_ (.LO(wbs_dat_o[5]));
 sky130_fd_sc_hd__conb_1 _462_ (.LO(wbs_dat_o[6]));
 sky130_fd_sc_hd__conb_1 _463_ (.LO(wbs_dat_o[7]));
 sky130_fd_sc_hd__conb_1 _464_ (.LO(wbs_dat_o[8]));
 sky130_fd_sc_hd__conb_1 _465_ (.LO(wbs_dat_o[9]));
 sky130_fd_sc_hd__conb_1 _466_ (.LO(wbs_dat_o[10]));
 sky130_fd_sc_hd__conb_1 _467_ (.LO(wbs_dat_o[11]));
 sky130_fd_sc_hd__conb_1 _468_ (.LO(wbs_dat_o[12]));
 sky130_fd_sc_hd__conb_1 _469_ (.LO(wbs_dat_o[13]));
 sky130_fd_sc_hd__conb_1 _470_ (.LO(wbs_dat_o[14]));
 sky130_fd_sc_hd__conb_1 _471_ (.LO(wbs_dat_o[15]));
 sky130_fd_sc_hd__conb_1 _472_ (.LO(wbs_dat_o[16]));
 sky130_fd_sc_hd__conb_1 _473_ (.LO(wbs_dat_o[17]));
 sky130_fd_sc_hd__conb_1 _474_ (.LO(wbs_dat_o[18]));
 sky130_fd_sc_hd__conb_1 _475_ (.LO(wbs_dat_o[19]));
 sky130_fd_sc_hd__conb_1 _476_ (.LO(wbs_dat_o[20]));
 sky130_fd_sc_hd__conb_1 _477_ (.LO(wbs_dat_o[21]));
 sky130_fd_sc_hd__conb_1 _478_ (.LO(wbs_dat_o[22]));
 sky130_fd_sc_hd__conb_1 _479_ (.LO(wbs_dat_o[23]));
 sky130_fd_sc_hd__conb_1 _480_ (.LO(wbs_dat_o[24]));
 sky130_fd_sc_hd__conb_1 _481_ (.LO(wbs_dat_o[25]));
 sky130_fd_sc_hd__conb_1 _482_ (.LO(wbs_dat_o[26]));
 sky130_fd_sc_hd__conb_1 _483_ (.LO(wbs_dat_o[27]));
 sky130_fd_sc_hd__conb_1 _484_ (.LO(wbs_dat_o[28]));
 sky130_fd_sc_hd__conb_1 _485_ (.LO(wbs_dat_o[29]));
 sky130_fd_sc_hd__conb_1 _486_ (.LO(wbs_dat_o[30]));
 sky130_fd_sc_hd__conb_1 _487_ (.LO(wbs_dat_o[31]));
 sky130_fd_sc_hd__conb_1 _488_ (.LO(_138_));
 sky130_fd_sc_hd__conb_1 _489_ (.LO(_139_));
 sky130_fd_sc_hd__conb_1 _490_ (.LO(_140_));
 sky130_fd_sc_hd__conb_1 _491_ (.LO(_141_));
 sky130_fd_sc_hd__conb_1 _492_ (.LO(_142_));
 sky130_fd_sc_hd__conb_1 _493_ (.LO(_143_));
 sky130_fd_sc_hd__conb_1 _494_ (.LO(_144_));
 sky130_fd_sc_hd__conb_1 _495_ (.LO(_145_));
 sky130_fd_sc_hd__conb_1 _496_ (.LO(_146_));
 sky130_fd_sc_hd__conb_1 _497_ (.LO(_147_));
 sky130_fd_sc_hd__conb_1 _498_ (.LO(_148_));
 sky130_fd_sc_hd__conb_1 _499_ (.LO(_149_));
 sky130_fd_sc_hd__conb_1 _500_ (.LO(_150_));
 sky130_fd_sc_hd__conb_1 _501_ (.LO(_151_));
 sky130_fd_sc_hd__conb_1 _502_ (.LO(_152_));
 sky130_fd_sc_hd__conb_1 _503_ (.LO(_153_));
 sky130_fd_sc_hd__conb_1 _504_ (.LO(_154_));
 sky130_fd_sc_hd__conb_1 _505_ (.LO(_155_));
 sky130_fd_sc_hd__conb_1 _506_ (.LO(_156_));
 sky130_fd_sc_hd__conb_1 _507_ (.LO(_157_));
 sky130_fd_sc_hd__conb_1 _508_ (.LO(_158_));
 sky130_fd_sc_hd__conb_1 _509_ (.LO(_159_));
 sky130_fd_sc_hd__conb_1 _510_ (.LO(_160_));
 sky130_fd_sc_hd__conb_1 _511_ (.LO(_161_));
 sky130_fd_sc_hd__conb_1 _512_ (.LO(_162_));
 sky130_fd_sc_hd__conb_1 _513_ (.LO(_163_));
 sky130_fd_sc_hd__conb_1 _514_ (.LO(_164_));
 sky130_fd_sc_hd__conb_1 _515_ (.LO(_165_));
 sky130_fd_sc_hd__conb_1 _516_ (.LO(_166_));
 sky130_fd_sc_hd__conb_1 _517_ (.LO(_167_));
 sky130_fd_sc_hd__conb_1 _518_ (.LO(_168_));
 sky130_fd_sc_hd__conb_1 _519_ (.LO(_169_));
 sky130_fd_sc_hd__conb_1 _520_ (.LO(io_oeb[0]));
 sky130_fd_sc_hd__conb_1 _521_ (.LO(io_oeb[1]));
 sky130_fd_sc_hd__conb_1 _522_ (.LO(io_oeb[2]));
 sky130_fd_sc_hd__conb_1 _523_ (.LO(io_oeb[3]));
 sky130_fd_sc_hd__conb_1 _524_ (.LO(io_oeb[4]));
 sky130_fd_sc_hd__conb_1 _525_ (.LO(io_oeb[5]));
 sky130_fd_sc_hd__conb_1 _526_ (.LO(io_oeb[6]));
 sky130_fd_sc_hd__conb_1 _527_ (.LO(io_oeb[7]));
 sky130_fd_sc_hd__conb_1 _528_ (.LO(io_oeb[8]));
 sky130_fd_sc_hd__conb_1 _529_ (.LO(io_oeb[9]));
 sky130_fd_sc_hd__conb_1 _530_ (.LO(io_oeb[10]));
 sky130_fd_sc_hd__conb_1 _531_ (.LO(io_oeb[11]));
 sky130_fd_sc_hd__conb_1 _532_ (.LO(io_oeb[12]));
 sky130_fd_sc_hd__conb_1 _533_ (.LO(io_oeb[13]));
 sky130_fd_sc_hd__conb_1 _534_ (.LO(io_oeb[14]));
 sky130_fd_sc_hd__conb_1 _535_ (.LO(io_oeb[15]));
 sky130_fd_sc_hd__conb_1 _536_ (.LO(io_oeb[16]));
 sky130_fd_sc_hd__conb_1 _537_ (.LO(io_oeb[17]));
 sky130_fd_sc_hd__conb_1 _538_ (.LO(io_oeb[18]));
 sky130_fd_sc_hd__conb_1 _539_ (.LO(io_oeb[19]));
 sky130_fd_sc_hd__conb_1 _540_ (.LO(io_oeb[20]));
 sky130_fd_sc_hd__conb_1 _541_ (.LO(io_oeb[21]));
 sky130_fd_sc_hd__conb_1 _542_ (.LO(io_oeb[22]));
 sky130_fd_sc_hd__conb_1 _543_ (.LO(io_oeb[23]));
 sky130_fd_sc_hd__conb_1 _544_ (.LO(io_oeb[24]));
 sky130_fd_sc_hd__conb_1 _545_ (.LO(io_oeb[25]));
 sky130_fd_sc_hd__conb_1 _546_ (.LO(io_oeb[26]));
 sky130_fd_sc_hd__conb_1 _547_ (.LO(io_oeb[27]));
 sky130_fd_sc_hd__ebufn_2 _548_ (.A(_138_),
    .TE_B(_106_),
    .Z(la_data_out[32]));
 sky130_fd_sc_hd__ebufn_2 _549_ (.A(_139_),
    .TE_B(_107_),
    .Z(la_data_out[33]));
 sky130_fd_sc_hd__ebufn_2 _550_ (.A(_140_),
    .TE_B(_108_),
    .Z(la_data_out[34]));
 sky130_fd_sc_hd__ebufn_2 _551_ (.A(_141_),
    .TE_B(_109_),
    .Z(la_data_out[35]));
 sky130_fd_sc_hd__ebufn_2 _552_ (.A(_142_),
    .TE_B(_110_),
    .Z(la_data_out[36]));
 sky130_fd_sc_hd__ebufn_2 _553_ (.A(_143_),
    .TE_B(_111_),
    .Z(la_data_out[37]));
 sky130_fd_sc_hd__ebufn_2 _554_ (.A(_144_),
    .TE_B(_112_),
    .Z(la_data_out[38]));
 sky130_fd_sc_hd__ebufn_2 _555_ (.A(_145_),
    .TE_B(_113_),
    .Z(la_data_out[39]));
 sky130_fd_sc_hd__ebufn_2 _556_ (.A(_146_),
    .TE_B(_114_),
    .Z(la_data_out[40]));
 sky130_fd_sc_hd__ebufn_2 _557_ (.A(_147_),
    .TE_B(_115_),
    .Z(la_data_out[41]));
 sky130_fd_sc_hd__ebufn_2 _558_ (.A(_148_),
    .TE_B(_116_),
    .Z(la_data_out[42]));
 sky130_fd_sc_hd__ebufn_2 _559_ (.A(_149_),
    .TE_B(_117_),
    .Z(la_data_out[43]));
 sky130_fd_sc_hd__ebufn_2 _560_ (.A(_150_),
    .TE_B(_118_),
    .Z(la_data_out[44]));
 sky130_fd_sc_hd__ebufn_2 _561_ (.A(_151_),
    .TE_B(_119_),
    .Z(la_data_out[45]));
 sky130_fd_sc_hd__ebufn_2 _562_ (.A(_152_),
    .TE_B(_120_),
    .Z(la_data_out[46]));
 sky130_fd_sc_hd__ebufn_2 _563_ (.A(_153_),
    .TE_B(_121_),
    .Z(la_data_out[47]));
 sky130_fd_sc_hd__ebufn_2 _564_ (.A(_154_),
    .TE_B(_122_),
    .Z(la_data_out[48]));
 sky130_fd_sc_hd__ebufn_2 _565_ (.A(_155_),
    .TE_B(_123_),
    .Z(la_data_out[49]));
 sky130_fd_sc_hd__ebufn_2 _566_ (.A(_156_),
    .TE_B(_124_),
    .Z(la_data_out[50]));
 sky130_fd_sc_hd__ebufn_2 _567_ (.A(_157_),
    .TE_B(_125_),
    .Z(la_data_out[51]));
 sky130_fd_sc_hd__ebufn_2 _568_ (.A(_158_),
    .TE_B(_126_),
    .Z(la_data_out[52]));
 sky130_fd_sc_hd__ebufn_2 _569_ (.A(_159_),
    .TE_B(_127_),
    .Z(la_data_out[53]));
 sky130_fd_sc_hd__ebufn_2 _570_ (.A(_160_),
    .TE_B(_128_),
    .Z(la_data_out[54]));
 sky130_fd_sc_hd__ebufn_2 _571_ (.A(_161_),
    .TE_B(_129_),
    .Z(la_data_out[55]));
 sky130_fd_sc_hd__ebufn_2 _572_ (.A(_162_),
    .TE_B(_130_),
    .Z(la_data_out[56]));
 sky130_fd_sc_hd__ebufn_2 _573_ (.A(_163_),
    .TE_B(_131_),
    .Z(la_data_out[57]));
 sky130_fd_sc_hd__ebufn_2 _574_ (.A(_164_),
    .TE_B(_132_),
    .Z(la_data_out[58]));
 sky130_fd_sc_hd__ebufn_2 _575_ (.A(_165_),
    .TE_B(_133_),
    .Z(la_data_out[59]));
 sky130_fd_sc_hd__ebufn_2 _576_ (.A(_166_),
    .TE_B(_134_),
    .Z(la_data_out[60]));
 sky130_fd_sc_hd__ebufn_2 _577_ (.A(_167_),
    .TE_B(_135_),
    .Z(la_data_out[61]));
 sky130_fd_sc_hd__ebufn_2 _578_ (.A(_168_),
    .TE_B(_136_),
    .Z(la_data_out[62]));
 sky130_fd_sc_hd__ebufn_2 _579_ (.A(_169_),
    .TE_B(_137_),
    .Z(la_data_out[63]));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__diode_2 ANTENNA__272__A2_N (.DIODE(_054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__268__B (.DIODE(_054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__321__C1 (.DIODE(_099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__270__C (.DIODE(_099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__270__A (.DIODE(_099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__203__A (.DIODE(_099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__197__A (.DIODE(_099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__172__A (.DIODE(_099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__262__A3 (.DIODE(io_in[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA__261__A2 (.DIODE(io_in[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA__260__A2_N (.DIODE(io_in[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA__222__B (.DIODE(io_in[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA__222__A (.DIODE(io_in[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA__276__B1 (.DIODE(io_in[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA__223__A (.DIODE(io_in[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA__221__B1 (.DIODE(io_in[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA__292__C (.DIODE(io_in[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA__292__A (.DIODE(io_in[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA__291__B (.DIODE(io_in[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA__290__A2 (.DIODE(io_in[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA__226__C (.DIODE(io_in[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA__226__A (.DIODE(io_in[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA__217__C (.DIODE(io_in[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA__217__A (.DIODE(io_in[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA__311__B1 (.DIODE(io_in[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA__225__C (.DIODE(io_in[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA__225__A (.DIODE(io_in[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA__214__C (.DIODE(io_in[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA__214__A (.DIODE(io_in[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA__220__A1 (.DIODE(io_in[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA__218__A (.DIODE(io_in[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA__215__A1 (.DIODE(io_in[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA__212__A2 (.DIODE(io_in[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA__220__B1_N (.DIODE(io_in[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA__210__A (.DIODE(io_in[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA__290__B1 (.DIODE(io_in[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA__216__C (.DIODE(io_in[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA__216__A (.DIODE(io_in[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA__212__A1 (.DIODE(io_in[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA__312__A1 (.DIODE(io_in[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA__311__A1 (.DIODE(io_in[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA__228__A1 (.DIODE(io_in[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA__213__C (.DIODE(io_in[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA__213__A (.DIODE(io_in[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA__266__A3 (.DIODE(io_in[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA__265__A2 (.DIODE(io_in[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA__264__A2_N (.DIODE(io_in[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA__245__B (.DIODE(io_in[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA__245__A (.DIODE(io_in[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA__282__B1 (.DIODE(io_in[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA__246__A (.DIODE(io_in[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA__244__B1 (.DIODE(io_in[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA__298__C (.DIODE(io_in[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA__298__A (.DIODE(io_in[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA__297__B (.DIODE(io_in[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA__296__A2 (.DIODE(io_in[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA__249__C (.DIODE(io_in[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA__249__A (.DIODE(io_in[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA__240__C (.DIODE(io_in[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA__240__A (.DIODE(io_in[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA__317__B1 (.DIODE(io_in[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA__248__C (.DIODE(io_in[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA__248__A (.DIODE(io_in[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA__237__C (.DIODE(io_in[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA__237__A (.DIODE(io_in[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA__243__A1 (.DIODE(io_in[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA__241__A (.DIODE(io_in[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA__238__A1 (.DIODE(io_in[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA__235__A2 (.DIODE(io_in[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA__243__B1_N (.DIODE(io_in[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA__233__A (.DIODE(io_in[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA__296__B1 (.DIODE(io_in[32]));
 sky130_fd_sc_hd__diode_2 ANTENNA__239__C (.DIODE(io_in[32]));
 sky130_fd_sc_hd__diode_2 ANTENNA__239__A (.DIODE(io_in[32]));
 sky130_fd_sc_hd__diode_2 ANTENNA__235__A1 (.DIODE(io_in[32]));
 sky130_fd_sc_hd__diode_2 ANTENNA__318__A1 (.DIODE(io_in[33]));
 sky130_fd_sc_hd__diode_2 ANTENNA__317__A1 (.DIODE(io_in[33]));
 sky130_fd_sc_hd__diode_2 ANTENNA__251__A1 (.DIODE(io_in[33]));
 sky130_fd_sc_hd__diode_2 ANTENNA__236__C (.DIODE(io_in[33]));
 sky130_fd_sc_hd__diode_2 ANTENNA__236__A (.DIODE(io_in[33]));
 sky130_fd_sc_hd__diode_2 ANTENNA__276__A2 (.DIODE(io_in[34]));
 sky130_fd_sc_hd__diode_2 ANTENNA__275__A (.DIODE(io_in[34]));
 sky130_fd_sc_hd__diode_2 ANTENNA__260__B2 (.DIODE(io_in[34]));
 sky130_fd_sc_hd__diode_2 ANTENNA__211__B (.DIODE(io_in[34]));
 sky130_fd_sc_hd__diode_2 ANTENNA__295__A1 (.DIODE(io_in[35]));
 sky130_fd_sc_hd__diode_2 ANTENNA__294__B1 (.DIODE(io_in[35]));
 sky130_fd_sc_hd__diode_2 ANTENNA__259__A (.DIODE(io_in[35]));
 sky130_fd_sc_hd__diode_2 ANTENNA__230__A (.DIODE(io_in[35]));
 sky130_fd_sc_hd__diode_2 ANTENNA__211__C (.DIODE(io_in[35]));
 sky130_fd_sc_hd__diode_2 ANTENNA__211__A_N (.DIODE(io_in[35]));
 sky130_fd_sc_hd__diode_2 ANTENNA__282__A2 (.DIODE(io_in[36]));
 sky130_fd_sc_hd__diode_2 ANTENNA__281__A (.DIODE(io_in[36]));
 sky130_fd_sc_hd__diode_2 ANTENNA__264__B2 (.DIODE(io_in[36]));
 sky130_fd_sc_hd__diode_2 ANTENNA__234__B (.DIODE(io_in[36]));
 sky130_fd_sc_hd__diode_2 ANTENNA__263__A (.DIODE(io_in[37]));
 sky130_fd_sc_hd__diode_2 ANTENNA__253__A (.DIODE(io_in[37]));
 sky130_fd_sc_hd__diode_2 ANTENNA__234__C (.DIODE(io_in[37]));
 sky130_fd_sc_hd__diode_2 ANTENNA__234__A_N (.DIODE(io_in[37]));
 sky130_fd_sc_hd__diode_2 ANTENNA__258__B1 (.DIODE(io_out[4]));
 sky130_fd_sc_hd__decap_6 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_513 ();
endmodule

