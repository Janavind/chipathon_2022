magic
tech sky130A
magscale 1 2
timestamp 1666199351
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 107 157 524 203
rect 1 21 827 157
rect 30 -17 64 21
<< scnmos >>
rect 81 47 111 131
rect 198 47 228 177
rect 415 47 445 177
rect 587 47 617 131
rect 673 47 703 131
<< scpmoshvt >>
rect 81 297 111 497
rect 198 333 228 497
rect 415 333 445 497
rect 587 297 617 497
rect 673 297 703 497
<< ndiff >>
rect 133 131 198 177
rect 27 101 81 131
rect 27 67 36 101
rect 70 67 81 101
rect 27 47 81 67
rect 111 101 198 131
rect 111 67 133 101
rect 167 67 198 101
rect 111 47 198 67
rect 228 101 309 177
rect 228 67 267 101
rect 301 67 309 101
rect 228 47 309 67
rect 363 101 415 177
rect 363 67 371 101
rect 405 67 415 101
rect 363 47 415 67
rect 445 131 498 177
rect 445 97 587 131
rect 445 63 526 97
rect 560 63 587 97
rect 445 47 587 63
rect 617 101 673 131
rect 617 67 628 101
rect 662 67 673 101
rect 617 47 673 67
rect 703 101 801 131
rect 703 67 759 101
rect 793 67 801 101
rect 703 47 801 67
<< pdiff >>
rect 27 477 81 497
rect 27 443 36 477
rect 70 443 81 477
rect 27 409 81 443
rect 27 375 36 409
rect 70 375 81 409
rect 27 297 81 375
rect 111 477 198 497
rect 111 443 136 477
rect 170 443 198 477
rect 111 333 198 443
rect 228 477 304 497
rect 228 443 262 477
rect 296 443 304 477
rect 228 409 304 443
rect 228 375 262 409
rect 296 375 304 409
rect 228 333 304 375
rect 362 477 415 497
rect 362 443 370 477
rect 404 443 415 477
rect 362 409 415 443
rect 362 375 370 409
rect 404 375 415 409
rect 362 333 415 375
rect 445 477 587 497
rect 445 443 526 477
rect 560 443 587 477
rect 445 333 587 443
rect 111 297 161 333
rect 537 297 587 333
rect 617 477 673 497
rect 617 443 628 477
rect 662 443 673 477
rect 617 388 673 443
rect 617 354 628 388
rect 662 354 673 388
rect 617 297 673 354
rect 703 477 801 497
rect 703 443 759 477
rect 793 443 801 477
rect 703 388 801 443
rect 703 354 759 388
rect 793 354 801 388
rect 703 297 801 354
<< ndiffc >>
rect 36 67 70 101
rect 133 67 167 101
rect 267 67 301 101
rect 371 67 405 101
rect 526 63 560 97
rect 628 67 662 101
rect 759 67 793 101
<< pdiffc >>
rect 36 443 70 477
rect 36 375 70 409
rect 136 443 170 477
rect 262 443 296 477
rect 262 375 296 409
rect 370 443 404 477
rect 370 375 404 409
rect 526 443 560 477
rect 628 443 662 477
rect 628 354 662 388
rect 759 443 793 477
rect 759 354 793 388
<< poly >>
rect 81 497 111 523
rect 198 497 228 523
rect 415 497 445 523
rect 587 497 617 523
rect 673 497 703 523
rect 81 259 111 297
rect 44 249 111 259
rect 44 215 60 249
rect 94 215 111 249
rect 44 205 111 215
rect 81 131 111 205
rect 198 259 228 333
rect 415 259 445 333
rect 587 259 617 297
rect 673 259 703 297
rect 198 249 264 259
rect 198 215 214 249
rect 248 215 264 249
rect 198 205 264 215
rect 349 249 483 259
rect 349 215 365 249
rect 399 215 433 249
rect 467 215 483 249
rect 349 205 483 215
rect 571 249 703 259
rect 571 215 587 249
rect 621 215 703 249
rect 571 205 703 215
rect 198 177 228 205
rect 415 177 445 205
rect 587 131 617 205
rect 673 131 703 205
rect 81 21 111 47
rect 198 21 228 47
rect 415 21 445 47
rect 587 21 617 47
rect 673 21 703 47
<< polycont >>
rect 60 215 94 249
rect 214 215 248 249
rect 365 215 399 249
rect 433 215 467 249
rect 587 215 621 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 17 477 86 493
rect 17 443 36 477
rect 70 443 86 477
rect 17 409 86 443
rect 120 477 186 527
rect 120 443 136 477
rect 170 443 186 477
rect 120 427 186 443
rect 246 477 332 493
rect 246 443 262 477
rect 296 443 332 477
rect 17 375 36 409
rect 70 393 86 409
rect 246 409 332 443
rect 70 375 212 393
rect 17 359 212 375
rect 17 249 111 325
rect 17 215 60 249
rect 94 215 111 249
rect 17 212 111 215
rect 178 249 212 359
rect 246 375 262 409
rect 296 375 332 409
rect 246 357 332 375
rect 366 477 420 493
rect 366 443 370 477
rect 404 443 420 477
rect 366 409 420 443
rect 510 477 576 527
rect 510 443 526 477
rect 560 443 576 477
rect 510 427 576 443
rect 614 477 710 493
rect 614 443 628 477
rect 662 443 710 477
rect 366 375 370 409
rect 404 393 420 409
rect 404 375 580 393
rect 366 358 580 375
rect 298 297 332 357
rect 298 249 483 297
rect 178 215 214 249
rect 248 215 264 249
rect 298 215 365 249
rect 399 215 433 249
rect 467 215 483 249
rect 546 249 580 358
rect 614 388 710 443
rect 614 354 628 388
rect 662 354 710 388
rect 614 297 710 354
rect 744 477 811 527
rect 744 443 759 477
rect 793 443 811 477
rect 744 388 811 443
rect 744 354 759 388
rect 793 354 811 388
rect 744 297 811 354
rect 546 215 587 249
rect 621 215 637 249
rect 178 178 212 215
rect 298 181 332 215
rect 546 181 580 215
rect 17 144 212 178
rect 17 101 83 144
rect 17 67 36 101
rect 70 67 83 101
rect 17 51 83 67
rect 117 101 183 110
rect 117 67 133 101
rect 167 67 183 101
rect 117 17 183 67
rect 256 101 332 181
rect 256 67 267 101
rect 301 67 332 101
rect 256 51 332 67
rect 366 147 580 181
rect 366 101 420 147
rect 671 128 710 297
rect 366 67 371 101
rect 405 67 420 101
rect 366 51 420 67
rect 510 97 576 113
rect 510 63 526 97
rect 560 63 576 97
rect 510 17 576 63
rect 610 101 710 128
rect 610 67 628 101
rect 662 67 710 101
rect 610 51 710 67
rect 744 101 811 129
rect 744 67 759 101
rect 793 67 811 101
rect 744 17 811 67
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
flabel locali s 30 289 64 323 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 673 425 707 459 0 FreeSans 400 0 0 0 X
port 6 nsew signal output
flabel locali s 673 357 707 391 0 FreeSans 400 0 0 0 X
port 6 nsew signal output
flabel locali s 673 289 707 323 0 FreeSans 400 0 0 0 X
port 6 nsew signal output
flabel locali s 673 221 707 255 0 FreeSans 400 0 0 0 X
port 6 nsew signal output
flabel locali s 673 153 707 187 0 FreeSans 400 0 0 0 X
port 6 nsew signal output
flabel locali s 673 85 707 119 0 FreeSans 400 0 0 0 X
port 6 nsew signal output
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power bidirectional abutment
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground bidirectional abutment
rlabel comment s 0 0 0 0 4 clkdlybuf4s15_2
rlabel metal1 s 0 -48 828 48 1 VGND
port 2 nsew ground bidirectional abutment
rlabel metal1 s 0 496 828 592 1 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 828 544
string GDS_END 3265580
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3259014
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 20.700 0.000 
<< end >>
