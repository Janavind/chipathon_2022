magic
tech sky130A
magscale 1 2
timestamp 1666464484
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 188 157 641 203
rect 1 21 641 157
rect 29 -17 63 21
<< locali >>
rect 17 199 65 277
rect 557 339 627 493
rect 389 289 627 339
rect 473 169 523 289
rect 557 215 627 255
rect 473 119 539 169
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 17 345 69 493
rect 103 379 179 527
rect 214 417 248 493
rect 282 451 455 527
rect 489 417 523 493
rect 214 373 523 417
rect 17 311 179 345
rect 99 255 179 311
rect 214 289 355 373
rect 99 199 407 255
rect 99 165 168 199
rect 17 131 168 165
rect 203 131 439 165
rect 17 51 69 131
rect 103 17 169 97
rect 203 51 256 131
rect 290 17 356 97
rect 390 85 439 131
rect 573 85 627 155
rect 390 51 627 85
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel locali s 557 215 627 255 6 A
port 1 nsew signal input
rlabel locali s 17 199 65 277 6 TE_B
port 2 nsew signal input
rlabel metal1 s 0 -48 644 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 1 21 641 157 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 188 157 641 203 6 VNB
port 4 nsew ground bidirectional
rlabel nwell s -38 261 682 582 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 496 644 592 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 473 119 539 169 6 Z
port 7 nsew signal output
rlabel locali s 473 169 523 289 6 Z
port 7 nsew signal output
rlabel locali s 389 289 627 339 6 Z
port 7 nsew signal output
rlabel locali s 557 339 627 493 6 Z
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 644 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2972072
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2965786
<< end >>
