magic
tech sky130B
magscale 1 2
timestamp 1666199351
<< metal1 >>
rect 4549 3491 4555 3543
rect 4607 3491 4613 3543
rect 4425 2153 4431 2205
rect 4483 2153 4489 2205
rect 4301 663 4307 715
rect 4359 663 4365 715
rect 3251 -2014 3257 -1962
rect 3309 -1974 3315 -1962
rect 4425 -1974 4431 -1962
rect 3309 -2002 4431 -1974
rect 3309 -2014 3315 -2002
rect 4425 -2014 4431 -2002
rect 4483 -2014 4489 -1962
rect 4419 -2116 4425 -2064
rect 4477 -2076 4483 -2064
rect 4549 -2076 4555 -2064
rect 4477 -2104 4555 -2076
rect 4477 -2116 4483 -2104
rect 4549 -2116 4555 -2104
rect 4607 -2116 4613 -2064
rect 2083 -2218 2089 -2166
rect 2141 -2178 2147 -2166
rect 4301 -2178 4307 -2166
rect 2141 -2206 4307 -2178
rect 2141 -2218 2147 -2206
rect 4301 -2218 4307 -2206
rect 4359 -2218 4365 -2166
<< via1 >>
rect 4555 3491 4607 3543
rect 4431 2153 4483 2205
rect 4307 663 4359 715
rect 3257 -2014 3309 -1962
rect 4431 -2014 4483 -1962
rect 4425 -2116 4477 -2064
rect 4555 -2116 4607 -2064
rect 2089 -2218 2141 -2166
rect 4307 -2218 4359 -2166
<< metal2 >>
rect 4555 3543 4607 3549
rect 4555 3485 4607 3491
rect 4431 2205 4483 2211
rect 4431 2147 4483 2153
rect 4307 715 4359 721
rect 4307 657 4359 663
rect 3257 -1962 3309 -1956
rect 3257 -2020 3309 -2014
rect 2089 -2166 2141 -2160
rect 2089 -2224 2141 -2218
rect 2101 -3207 2129 -2224
rect 3269 -3207 3297 -2020
rect 4319 -2160 4347 657
rect 4443 -1956 4471 2147
rect 4431 -1962 4483 -1956
rect 4431 -2020 4483 -2014
rect 4567 -2058 4595 3485
rect 4425 -2064 4477 -2058
rect 4425 -2122 4477 -2116
rect 4555 -2064 4607 -2058
rect 4555 -2122 4607 -2116
rect 4307 -2166 4359 -2160
rect 4307 -2224 4359 -2218
rect 4437 -3207 4465 -2122
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_0
timestamp 1666199351
transform 1 0 3251 0 1 -2020
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_1
timestamp 1666199351
transform 1 0 4425 0 1 2147
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_2
timestamp 1666199351
transform 1 0 4425 0 1 -2020
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_3
timestamp 1666199351
transform 1 0 4419 0 1 -2122
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_4
timestamp 1666199351
transform 1 0 4549 0 1 3485
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_5
timestamp 1666199351
transform 1 0 4549 0 1 -2122
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_6
timestamp 1666199351
transform 1 0 2083 0 1 -2224
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_7
timestamp 1666199351
transform 1 0 4301 0 1 657
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_8
timestamp 1666199351
transform 1 0 4301 0 1 -2224
box 0 0 1 1
<< properties >>
string FIXED_BBOX 2083 -3207 4613 3549
string GDS_END 7033170
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_8x1024_8.gds
string GDS_START 7031604
<< end >>
