magic
tech sky130B
magscale 1 2
timestamp 1666199351
<< nwell >>
rect -38 261 2246 582
<< pwell >>
rect 1165 157 1347 201
rect 1650 157 2205 203
rect 1 145 817 157
rect 1019 145 2205 157
rect 1 21 2205 145
rect 29 -17 63 21
<< locali >>
rect 19 195 89 325
rect 352 176 386 337
rect 488 271 555 337
rect 352 175 388 176
rect 352 174 389 175
rect 352 172 390 174
rect 352 171 391 172
rect 352 170 392 171
rect 352 168 393 170
rect 352 167 394 168
rect 352 164 395 167
rect 352 162 398 164
rect 352 157 402 162
rect 613 157 647 223
rect 703 211 799 331
rect 352 150 647 157
rect 358 147 647 150
rect 361 145 647 147
rect 364 143 647 145
rect 366 141 647 143
rect 368 138 647 141
rect 372 131 647 138
rect 375 123 647 131
rect 491 61 526 123
rect 1840 308 1906 493
rect 1840 301 1922 308
rect 1871 286 1922 301
rect 1878 165 1922 286
rect 1836 158 1922 165
rect 2137 289 2188 465
rect 1836 145 1912 158
rect 1836 61 1906 145
rect 2146 159 2188 289
rect 2137 53 2188 159
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2208 561
rect 35 393 69 493
rect 103 427 169 527
rect 35 359 169 393
rect 123 194 169 359
rect 123 161 162 194
rect 35 127 162 161
rect 35 69 69 127
rect 103 17 169 93
rect 203 69 237 493
rect 284 415 341 489
rect 375 449 441 527
rect 535 449 714 483
rect 284 372 646 415
rect 284 117 318 372
rect 420 225 454 372
rect 612 337 646 372
rect 680 399 714 449
rect 748 433 782 527
rect 833 414 890 488
rect 929 438 1143 472
rect 833 399 867 414
rect 680 365 867 399
rect 612 271 651 337
rect 420 191 489 225
rect 833 177 867 365
rect 681 143 867 177
rect 284 51 341 117
rect 391 17 457 89
rect 681 89 715 143
rect 560 55 715 89
rect 749 17 789 109
rect 833 107 867 143
rect 901 207 949 381
rect 987 331 1075 402
rect 1109 315 1143 438
rect 1177 367 1211 527
rect 1245 427 1295 493
rect 1340 433 1517 467
rect 1109 297 1211 315
rect 1051 263 1211 297
rect 901 141 1017 207
rect 1051 107 1085 263
rect 1177 249 1211 263
rect 1119 213 1153 219
rect 1245 213 1279 427
rect 1313 249 1351 393
rect 1385 315 1449 381
rect 1119 153 1279 213
rect 1385 207 1423 315
rect 1483 281 1517 433
rect 1553 427 1614 527
rect 1676 381 1734 491
rect 1551 315 1734 381
rect 1768 325 1802 527
rect 833 73 903 107
rect 937 73 1085 107
rect 1135 17 1209 117
rect 1245 107 1279 153
rect 1313 141 1423 207
rect 1457 265 1517 281
rect 1697 265 1734 315
rect 1940 337 2006 485
rect 1457 199 1663 265
rect 1697 199 1844 265
rect 1457 107 1491 199
rect 1697 165 1734 199
rect 1245 73 1337 107
rect 1383 73 1491 107
rect 1540 17 1614 123
rect 1668 60 1734 165
rect 1956 265 2006 337
rect 2042 299 2103 527
rect 1956 199 2112 265
rect 1768 17 1802 139
rect 1956 124 1990 199
rect 1940 69 1990 124
rect 2037 17 2103 161
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2208 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
<< metal1 >>
rect 0 561 2208 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2208 561
rect 0 496 2208 527
rect 0 17 2208 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2208 17
rect 0 -48 2208 -17
<< obsm1 >>
rect 117 388 175 397
rect 1021 388 1079 397
rect 1303 388 1361 397
rect 117 360 1361 388
rect 117 351 175 360
rect 1021 351 1079 360
rect 1303 351 1361 360
rect 191 184 249 193
rect 937 184 995 193
rect 1305 184 1363 193
rect 191 156 1363 184
rect 191 147 249 156
rect 937 147 995 156
rect 1305 147 1363 156
<< labels >>
rlabel locali s 19 195 89 325 6 CLK
port 1 nsew clock input
rlabel locali s 488 271 555 337 6 D
port 2 nsew signal input
rlabel locali s 703 211 799 331 6 SCD
port 3 nsew signal input
rlabel locali s 491 61 526 123 6 SCE
port 4 nsew signal input
rlabel locali s 375 123 647 131 6 SCE
port 4 nsew signal input
rlabel locali s 372 131 647 138 6 SCE
port 4 nsew signal input
rlabel locali s 368 138 647 141 6 SCE
port 4 nsew signal input
rlabel locali s 366 141 647 143 6 SCE
port 4 nsew signal input
rlabel locali s 364 143 647 145 6 SCE
port 4 nsew signal input
rlabel locali s 361 145 647 147 6 SCE
port 4 nsew signal input
rlabel locali s 358 147 647 150 6 SCE
port 4 nsew signal input
rlabel locali s 352 150 647 157 6 SCE
port 4 nsew signal input
rlabel locali s 613 157 647 223 6 SCE
port 4 nsew signal input
rlabel locali s 352 157 402 162 6 SCE
port 4 nsew signal input
rlabel locali s 352 162 398 164 6 SCE
port 4 nsew signal input
rlabel locali s 352 164 395 167 6 SCE
port 4 nsew signal input
rlabel locali s 352 167 394 168 6 SCE
port 4 nsew signal input
rlabel locali s 352 168 393 170 6 SCE
port 4 nsew signal input
rlabel locali s 352 170 392 171 6 SCE
port 4 nsew signal input
rlabel locali s 352 171 391 172 6 SCE
port 4 nsew signal input
rlabel locali s 352 172 390 174 6 SCE
port 4 nsew signal input
rlabel locali s 352 174 389 175 6 SCE
port 4 nsew signal input
rlabel locali s 352 175 388 176 6 SCE
port 4 nsew signal input
rlabel locali s 352 176 386 337 6 SCE
port 4 nsew signal input
rlabel metal1 s 0 -48 2208 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 21 2205 145 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1019 145 2205 157 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 145 817 157 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1650 157 2205 203 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1165 157 1347 201 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 2246 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 2208 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1836 61 1906 145 6 Q
port 9 nsew signal output
rlabel locali s 1836 145 1912 158 6 Q
port 9 nsew signal output
rlabel locali s 1836 158 1922 165 6 Q
port 9 nsew signal output
rlabel locali s 1878 165 1922 286 6 Q
port 9 nsew signal output
rlabel locali s 1871 286 1922 301 6 Q
port 9 nsew signal output
rlabel locali s 1840 301 1922 308 6 Q
port 9 nsew signal output
rlabel locali s 1840 308 1906 493 6 Q
port 9 nsew signal output
rlabel locali s 2137 53 2188 159 6 Q_N
port 10 nsew signal output
rlabel locali s 2146 159 2188 289 6 Q_N
port 10 nsew signal output
rlabel locali s 2137 289 2188 465 6 Q_N
port 10 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2208 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 343100
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 326098
<< end >>
