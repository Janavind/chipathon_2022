magic
tech sky130A
magscale 1 2
timestamp 1666199351
use sky130_fd_pr__hvdfl1sd2__example_55959141808491  sky130_fd_pr__hvdfl1sd2__example_55959141808491_0
timestamp 1666199351
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808491  sky130_fd_pr__hvdfl1sd2__example_55959141808491_1
timestamp 1666199351
transform 1 0 256 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808476  sky130_fd_pr__hvdfl1sd__example_55959141808476_0
timestamp 1666199351
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808476  sky130_fd_pr__hvdfl1sd__example_55959141808476_1
timestamp 1666199351
transform 1 0 412 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 29505478
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 29503388
<< end >>
