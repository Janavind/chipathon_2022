magic
tech sky130B
magscale 1 2
timestamp 1666199351
<< pwell >>
rect 15 163 627 817
<< nmoslvt >>
rect 171 189 201 791
rect 257 189 293 791
rect 349 189 385 791
rect 441 189 471 791
<< ndiff >>
rect 111 779 171 791
rect 111 745 126 779
rect 160 745 171 779
rect 111 711 171 745
rect 111 677 126 711
rect 160 677 171 711
rect 111 643 171 677
rect 111 609 126 643
rect 160 609 171 643
rect 111 575 171 609
rect 111 541 126 575
rect 160 541 171 575
rect 111 507 171 541
rect 111 473 126 507
rect 160 473 171 507
rect 111 439 171 473
rect 111 405 126 439
rect 160 405 171 439
rect 111 371 171 405
rect 111 337 126 371
rect 160 337 171 371
rect 111 303 171 337
rect 111 269 126 303
rect 160 269 171 303
rect 111 235 171 269
rect 111 201 126 235
rect 160 201 171 235
rect 111 189 171 201
rect 201 779 257 791
rect 201 513 212 779
rect 246 513 257 779
rect 201 467 257 513
rect 201 201 212 467
rect 246 201 257 467
rect 201 189 257 201
rect 293 779 349 791
rect 293 513 304 779
rect 338 513 349 779
rect 293 467 349 513
rect 293 201 304 467
rect 338 201 349 467
rect 293 189 349 201
rect 385 779 441 791
rect 385 513 396 779
rect 430 513 441 779
rect 385 467 441 513
rect 385 201 396 467
rect 430 201 441 467
rect 385 189 441 201
rect 471 779 531 791
rect 471 745 482 779
rect 516 745 531 779
rect 471 711 531 745
rect 471 677 482 711
rect 516 677 531 711
rect 471 643 531 677
rect 471 609 482 643
rect 516 609 531 643
rect 471 575 531 609
rect 471 541 482 575
rect 516 541 531 575
rect 471 507 531 541
rect 471 473 482 507
rect 516 473 531 507
rect 471 439 531 473
rect 471 405 482 439
rect 516 405 531 439
rect 471 371 531 405
rect 471 337 482 371
rect 516 337 531 371
rect 471 303 531 337
rect 471 269 482 303
rect 516 269 531 303
rect 471 235 531 269
rect 471 201 482 235
rect 516 201 531 235
rect 471 189 531 201
<< ndiffc >>
rect 126 745 160 779
rect 126 677 160 711
rect 126 609 160 643
rect 126 541 160 575
rect 126 473 160 507
rect 126 405 160 439
rect 126 337 160 371
rect 126 269 160 303
rect 126 201 160 235
rect 212 513 246 779
rect 212 201 246 467
rect 304 513 338 779
rect 304 201 338 467
rect 396 513 430 779
rect 396 201 430 467
rect 482 745 516 779
rect 482 677 516 711
rect 482 609 516 643
rect 482 541 516 575
rect 482 473 516 507
rect 482 405 516 439
rect 482 337 516 371
rect 482 269 516 303
rect 482 201 516 235
<< psubdiff >>
rect 41 779 111 791
rect 41 745 58 779
rect 92 745 111 779
rect 41 711 111 745
rect 41 677 58 711
rect 92 677 111 711
rect 41 643 111 677
rect 41 609 58 643
rect 92 609 111 643
rect 41 575 111 609
rect 41 541 58 575
rect 92 541 111 575
rect 41 507 111 541
rect 41 473 58 507
rect 92 473 111 507
rect 41 439 111 473
rect 41 405 58 439
rect 92 405 111 439
rect 41 371 111 405
rect 41 337 58 371
rect 92 337 111 371
rect 41 303 111 337
rect 41 269 58 303
rect 92 269 111 303
rect 41 235 111 269
rect 41 201 58 235
rect 92 201 111 235
rect 41 189 111 201
rect 531 779 601 791
rect 531 745 550 779
rect 584 745 601 779
rect 531 711 601 745
rect 531 677 550 711
rect 584 677 601 711
rect 531 643 601 677
rect 531 609 550 643
rect 584 609 601 643
rect 531 575 601 609
rect 531 541 550 575
rect 584 541 601 575
rect 531 507 601 541
rect 531 473 550 507
rect 584 473 601 507
rect 531 439 601 473
rect 531 405 550 439
rect 584 405 601 439
rect 531 371 601 405
rect 531 337 550 371
rect 584 337 601 371
rect 531 303 601 337
rect 531 269 550 303
rect 584 269 601 303
rect 531 235 601 269
rect 531 201 550 235
rect 584 201 601 235
rect 531 189 601 201
<< psubdiffcont >>
rect 58 745 92 779
rect 58 677 92 711
rect 58 609 92 643
rect 58 541 92 575
rect 58 473 92 507
rect 58 405 92 439
rect 58 337 92 371
rect 58 269 92 303
rect 58 201 92 235
rect 550 745 584 779
rect 550 677 584 711
rect 550 609 584 643
rect 550 541 584 575
rect 550 473 584 507
rect 550 405 584 439
rect 550 337 584 371
rect 550 269 584 303
rect 550 201 584 235
<< poly >>
rect 243 891 399 907
rect 120 867 201 883
rect 120 833 136 867
rect 170 833 201 867
rect 243 857 264 891
rect 378 857 399 891
rect 243 841 399 857
rect 441 867 522 883
rect 120 817 201 833
rect 171 791 201 817
rect 257 791 293 841
rect 349 791 385 841
rect 441 833 472 867
rect 506 833 522 867
rect 441 817 522 833
rect 441 791 471 817
rect 171 163 201 189
rect 120 147 201 163
rect 120 113 136 147
rect 170 113 201 147
rect 257 139 293 189
rect 349 139 385 189
rect 441 163 471 189
rect 441 147 522 163
rect 120 97 201 113
rect 243 123 399 139
rect 243 89 264 123
rect 378 89 399 123
rect 441 113 472 147
rect 506 113 522 147
rect 441 97 522 113
rect 243 73 399 89
<< polycont >>
rect 136 833 170 867
rect 264 857 378 891
rect 472 833 506 867
rect 136 113 170 147
rect 264 89 378 123
rect 472 113 506 147
<< locali >>
rect 248 961 394 980
rect 248 927 262 961
rect 296 927 346 961
rect 380 927 394 961
rect 248 891 394 927
rect 248 889 264 891
rect 378 889 394 891
rect 120 867 186 883
rect 120 833 136 867
rect 170 833 186 867
rect 248 855 262 889
rect 296 855 346 857
rect 380 855 394 889
rect 248 841 394 855
rect 456 867 522 883
rect 120 817 186 833
rect 456 833 472 867
rect 506 833 522 867
rect 456 817 522 833
rect 120 795 160 817
rect 482 795 522 817
rect 41 779 160 795
rect 41 745 58 779
rect 92 759 126 779
rect 94 745 126 759
rect 41 725 60 745
rect 94 725 160 745
rect 41 711 160 725
rect 41 677 58 711
rect 92 687 126 711
rect 94 677 126 687
rect 41 653 60 677
rect 94 653 160 677
rect 41 643 160 653
rect 41 609 58 643
rect 92 615 126 643
rect 94 609 126 615
rect 41 581 60 609
rect 94 581 160 609
rect 41 575 160 581
rect 41 541 58 575
rect 92 543 126 575
rect 94 541 126 543
rect 41 509 60 541
rect 94 509 160 541
rect 41 507 160 509
rect 41 473 58 507
rect 92 473 126 507
rect 41 471 160 473
rect 41 439 60 471
rect 94 439 160 471
rect 41 405 58 439
rect 94 437 126 439
rect 92 405 126 437
rect 41 399 160 405
rect 41 371 60 399
rect 94 371 160 399
rect 41 337 58 371
rect 94 365 126 371
rect 92 337 126 365
rect 41 327 160 337
rect 41 303 60 327
rect 94 303 160 327
rect 41 269 58 303
rect 94 293 126 303
rect 92 269 126 293
rect 41 255 160 269
rect 41 235 60 255
rect 94 235 160 255
rect 41 201 58 235
rect 94 221 126 235
rect 92 201 126 221
rect 41 185 160 201
rect 212 779 246 795
rect 212 471 246 509
rect 212 185 246 201
rect 304 779 338 795
rect 304 471 338 509
rect 304 185 338 201
rect 396 779 430 795
rect 396 471 430 509
rect 396 185 430 201
rect 482 779 601 795
rect 516 759 550 779
rect 516 745 548 759
rect 584 745 601 779
rect 482 725 548 745
rect 582 725 601 745
rect 482 711 601 725
rect 516 687 550 711
rect 516 677 548 687
rect 584 677 601 711
rect 482 653 548 677
rect 582 653 601 677
rect 482 643 601 653
rect 516 615 550 643
rect 516 609 548 615
rect 584 609 601 643
rect 482 581 548 609
rect 582 581 601 609
rect 482 575 601 581
rect 516 543 550 575
rect 516 541 548 543
rect 584 541 601 575
rect 482 509 548 541
rect 582 509 601 541
rect 482 507 601 509
rect 516 473 550 507
rect 584 473 601 507
rect 482 471 601 473
rect 482 439 548 471
rect 582 439 601 471
rect 516 437 548 439
rect 516 405 550 437
rect 584 405 601 439
rect 482 399 601 405
rect 482 371 548 399
rect 582 371 601 399
rect 516 365 548 371
rect 516 337 550 365
rect 584 337 601 371
rect 482 327 601 337
rect 482 303 548 327
rect 582 303 601 327
rect 516 293 548 303
rect 516 269 550 293
rect 584 269 601 303
rect 482 255 601 269
rect 482 235 548 255
rect 582 235 601 255
rect 516 221 548 235
rect 516 201 550 221
rect 584 201 601 235
rect 482 185 601 201
rect 120 163 160 185
rect 482 163 522 185
rect 120 147 186 163
rect 120 113 136 147
rect 170 113 186 147
rect 456 147 522 163
rect 120 97 186 113
rect 248 125 394 139
rect 248 91 262 125
rect 296 123 346 125
rect 380 91 394 125
rect 456 113 472 147
rect 506 113 522 147
rect 456 97 522 113
rect 248 89 264 91
rect 378 89 394 91
rect 248 53 394 89
rect 248 19 262 53
rect 296 19 346 53
rect 380 19 394 53
rect 248 0 394 19
<< viali >>
rect 262 927 296 961
rect 346 927 380 961
rect 262 857 264 889
rect 264 857 296 889
rect 346 857 378 889
rect 378 857 380 889
rect 262 855 296 857
rect 346 855 380 857
rect 60 745 92 759
rect 92 745 94 759
rect 60 725 94 745
rect 60 677 92 687
rect 92 677 94 687
rect 60 653 94 677
rect 60 609 92 615
rect 92 609 94 615
rect 60 581 94 609
rect 60 541 92 543
rect 92 541 94 543
rect 60 509 94 541
rect 60 439 94 471
rect 60 437 92 439
rect 92 437 94 439
rect 60 371 94 399
rect 60 365 92 371
rect 92 365 94 371
rect 60 303 94 327
rect 60 293 92 303
rect 92 293 94 303
rect 60 235 94 255
rect 60 221 92 235
rect 92 221 94 235
rect 212 725 246 759
rect 212 653 246 687
rect 212 581 246 615
rect 212 513 246 543
rect 212 509 246 513
rect 212 467 246 471
rect 212 437 246 467
rect 212 365 246 399
rect 212 293 246 327
rect 212 221 246 255
rect 304 725 338 759
rect 304 653 338 687
rect 304 581 338 615
rect 304 513 338 543
rect 304 509 338 513
rect 304 467 338 471
rect 304 437 338 467
rect 304 365 338 399
rect 304 293 338 327
rect 304 221 338 255
rect 396 725 430 759
rect 396 653 430 687
rect 396 581 430 615
rect 396 513 430 543
rect 396 509 430 513
rect 396 467 430 471
rect 396 437 430 467
rect 396 365 430 399
rect 396 293 430 327
rect 396 221 430 255
rect 548 745 550 759
rect 550 745 582 759
rect 548 725 582 745
rect 548 677 550 687
rect 550 677 582 687
rect 548 653 582 677
rect 548 609 550 615
rect 550 609 582 615
rect 548 581 582 609
rect 548 541 550 543
rect 550 541 582 543
rect 548 509 582 541
rect 548 439 582 471
rect 548 437 550 439
rect 550 437 582 439
rect 548 371 582 399
rect 548 365 550 371
rect 550 365 582 371
rect 548 303 582 327
rect 548 293 550 303
rect 550 293 582 303
rect 548 235 582 255
rect 548 221 550 235
rect 550 221 582 235
rect 262 123 296 125
rect 346 123 380 125
rect 262 91 264 123
rect 264 91 296 123
rect 346 91 378 123
rect 378 91 380 123
rect 262 19 296 53
rect 346 19 380 53
<< metal1 >>
rect 250 961 392 980
rect 250 927 262 961
rect 296 927 346 961
rect 380 927 392 961
rect 250 889 392 927
rect 250 855 262 889
rect 296 855 346 889
rect 380 855 392 889
rect 250 843 392 855
rect 41 759 100 771
rect 41 725 60 759
rect 94 725 100 759
rect 41 687 100 725
rect 41 653 60 687
rect 94 653 100 687
rect 41 615 100 653
rect 41 581 60 615
rect 94 581 100 615
rect 41 543 100 581
rect 41 509 60 543
rect 94 509 100 543
rect 41 471 100 509
rect 41 437 60 471
rect 94 437 100 471
rect 41 399 100 437
rect 41 365 60 399
rect 94 365 100 399
rect 41 327 100 365
rect 41 293 60 327
rect 94 293 100 327
rect 41 255 100 293
rect 41 221 60 255
rect 94 221 100 255
rect 41 209 100 221
rect 203 759 255 771
rect 203 725 212 759
rect 246 725 255 759
rect 203 687 255 725
rect 203 653 212 687
rect 246 653 255 687
rect 203 615 255 653
rect 203 581 212 615
rect 246 581 255 615
rect 203 543 255 581
rect 203 509 212 543
rect 246 509 255 543
rect 203 471 255 509
rect 203 459 212 471
rect 246 459 255 471
rect 203 399 255 407
rect 203 395 212 399
rect 246 395 255 399
rect 203 331 255 343
rect 203 267 255 279
rect 203 209 255 215
rect 295 765 347 771
rect 295 701 347 713
rect 295 637 347 649
rect 295 581 304 585
rect 338 581 347 585
rect 295 573 347 581
rect 295 509 304 521
rect 338 509 347 521
rect 295 471 347 509
rect 295 437 304 471
rect 338 437 347 471
rect 295 399 347 437
rect 295 365 304 399
rect 338 365 347 399
rect 295 327 347 365
rect 295 293 304 327
rect 338 293 347 327
rect 295 255 347 293
rect 295 221 304 255
rect 338 221 347 255
rect 295 209 347 221
rect 387 759 439 771
rect 387 725 396 759
rect 430 725 439 759
rect 387 687 439 725
rect 387 653 396 687
rect 430 653 439 687
rect 387 615 439 653
rect 387 581 396 615
rect 430 581 439 615
rect 387 543 439 581
rect 387 509 396 543
rect 430 509 439 543
rect 387 471 439 509
rect 387 459 396 471
rect 430 459 439 471
rect 387 399 439 407
rect 387 395 396 399
rect 430 395 439 399
rect 387 331 439 343
rect 387 267 439 279
rect 387 209 439 215
rect 542 759 601 771
rect 542 725 548 759
rect 582 725 601 759
rect 542 687 601 725
rect 542 653 548 687
rect 582 653 601 687
rect 542 615 601 653
rect 542 581 548 615
rect 582 581 601 615
rect 542 543 601 581
rect 542 509 548 543
rect 582 509 601 543
rect 542 471 601 509
rect 542 437 548 471
rect 582 437 601 471
rect 542 399 601 437
rect 542 365 548 399
rect 582 365 601 399
rect 542 327 601 365
rect 542 293 548 327
rect 582 293 601 327
rect 542 255 601 293
rect 542 221 548 255
rect 582 221 601 255
rect 542 209 601 221
rect 250 125 392 137
rect 250 91 262 125
rect 296 91 346 125
rect 380 91 392 125
rect 250 53 392 91
rect 250 19 262 53
rect 296 19 346 53
rect 380 19 392 53
rect 250 0 392 19
<< via1 >>
rect 203 437 212 459
rect 212 437 246 459
rect 246 437 255 459
rect 203 407 255 437
rect 203 365 212 395
rect 212 365 246 395
rect 246 365 255 395
rect 203 343 255 365
rect 203 327 255 331
rect 203 293 212 327
rect 212 293 246 327
rect 246 293 255 327
rect 203 279 255 293
rect 203 255 255 267
rect 203 221 212 255
rect 212 221 246 255
rect 246 221 255 255
rect 203 215 255 221
rect 295 759 347 765
rect 295 725 304 759
rect 304 725 338 759
rect 338 725 347 759
rect 295 713 347 725
rect 295 687 347 701
rect 295 653 304 687
rect 304 653 338 687
rect 338 653 347 687
rect 295 649 347 653
rect 295 615 347 637
rect 295 585 304 615
rect 304 585 338 615
rect 338 585 347 615
rect 295 543 347 573
rect 295 521 304 543
rect 304 521 338 543
rect 338 521 347 543
rect 387 437 396 459
rect 396 437 430 459
rect 430 437 439 459
rect 387 407 439 437
rect 387 365 396 395
rect 396 365 430 395
rect 430 365 439 395
rect 387 343 439 365
rect 387 327 439 331
rect 387 293 396 327
rect 396 293 430 327
rect 430 293 439 327
rect 387 279 439 293
rect 387 255 439 267
rect 387 221 396 255
rect 396 221 430 255
rect 430 221 439 255
rect 387 215 439 221
<< metal2 >>
rect 14 765 628 771
rect 14 713 295 765
rect 347 713 628 765
rect 14 701 628 713
rect 14 649 295 701
rect 347 649 628 701
rect 14 637 628 649
rect 14 585 295 637
rect 347 585 628 637
rect 14 573 628 585
rect 14 521 295 573
rect 347 521 628 573
rect 14 515 628 521
rect 14 459 628 465
rect 14 407 203 459
rect 255 407 387 459
rect 439 407 628 459
rect 14 395 628 407
rect 14 343 203 395
rect 255 343 387 395
rect 439 343 628 395
rect 14 331 628 343
rect 14 279 203 331
rect 255 279 387 331
rect 439 279 628 331
rect 14 267 628 279
rect 14 215 203 267
rect 255 215 387 267
rect 439 215 628 267
rect 14 209 628 215
<< labels >>
flabel comment s 183 525 183 525 0 FreeSans 180 90 0 0 dummy_poly
flabel comment s 453 516 453 516 0 FreeSans 180 90 0 0 dummy_poly
flabel metal1 s 255 44 386 95 0 FreeSans 200 0 0 0 GATE
port 1 nsew
flabel metal1 s 255 880 386 931 0 FreeSans 200 0 0 0 GATE
port 1 nsew
flabel metal1 s 41 466 100 496 0 FreeSans 200 90 0 0 SUBSTRATE
port 2 nsew
flabel metal1 s 542 469 601 499 0 FreeSans 200 90 0 0 SUBSTRATE
port 2 nsew
flabel metal2 s 14 280 35 408 7 FreeSans 300 180 0 0 SOURCE
port 3 nsew
flabel metal2 s 14 589 35 717 7 FreeSans 300 180 0 0 DRAIN
port 4 nsew
<< properties >>
string GDS_END 4018836
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 4005972
<< end >>
