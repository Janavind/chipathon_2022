magic
tech sky130B
magscale 1 2
timestamp 1666464484
<< nwell >>
rect -38 261 2890 582
<< pwell >>
rect 1411 157 1769 201
rect 2190 157 2850 203
rect 1 21 2850 157
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 131
rect 151 47 181 131
rect 235 47 265 131
rect 328 47 358 131
rect 516 47 546 131
rect 704 47 734 131
rect 788 47 818 131
rect 976 47 1006 131
rect 1060 47 1090 131
rect 1132 47 1162 131
rect 1320 47 1350 131
rect 1392 47 1422 131
rect 1487 47 1517 175
rect 1663 47 1693 175
rect 1783 47 1813 131
rect 1855 47 1885 131
rect 1955 47 1985 131
rect 2052 47 2082 131
rect 2268 47 2298 177
rect 2352 47 2382 177
rect 2553 47 2583 131
rect 2648 47 2678 177
rect 2732 47 2762 177
<< scpmoshvt >>
rect 79 369 109 497
rect 163 369 193 497
rect 235 369 265 497
rect 331 369 361 497
rect 517 369 547 497
rect 705 369 735 497
rect 789 369 819 497
rect 977 413 1007 497
rect 1072 413 1102 497
rect 1162 413 1192 497
rect 1281 413 1311 497
rect 1379 413 1409 497
rect 1495 329 1525 497
rect 1567 329 1597 497
rect 1693 413 1723 497
rect 1781 413 1811 497
rect 1892 413 1922 497
rect 2080 413 2110 497
rect 2268 297 2298 497
rect 2352 297 2382 497
rect 2553 356 2583 484
rect 2648 297 2678 497
rect 2732 297 2762 497
<< ndiff >>
rect 1437 131 1487 175
rect 27 103 79 131
rect 27 69 35 103
rect 69 69 79 103
rect 27 47 79 69
rect 109 47 151 131
rect 181 98 235 131
rect 181 64 191 98
rect 225 64 235 98
rect 181 47 235 64
rect 265 47 328 131
rect 358 93 410 131
rect 358 59 368 93
rect 402 59 410 93
rect 358 47 410 59
rect 464 105 516 131
rect 464 71 472 105
rect 506 71 516 105
rect 464 47 516 71
rect 546 93 598 131
rect 546 59 556 93
rect 590 59 598 93
rect 546 47 598 59
rect 652 105 704 131
rect 652 71 660 105
rect 694 71 704 105
rect 652 47 704 71
rect 734 89 788 131
rect 734 55 744 89
rect 778 55 788 89
rect 734 47 788 55
rect 818 101 870 131
rect 818 67 828 101
rect 862 67 870 101
rect 818 47 870 67
rect 924 101 976 131
rect 924 67 932 101
rect 966 67 976 101
rect 924 47 976 67
rect 1006 101 1060 131
rect 1006 67 1016 101
rect 1050 67 1060 101
rect 1006 47 1060 67
rect 1090 47 1132 131
rect 1162 93 1214 131
rect 1162 59 1172 93
rect 1206 59 1214 93
rect 1162 47 1214 59
rect 1268 119 1320 131
rect 1268 85 1276 119
rect 1310 85 1320 119
rect 1268 47 1320 85
rect 1350 47 1392 131
rect 1422 89 1487 131
rect 1422 55 1432 89
rect 1466 55 1487 89
rect 1422 47 1487 55
rect 1517 47 1663 175
rect 1693 131 1743 175
rect 2216 161 2268 177
rect 1693 89 1783 131
rect 1693 55 1709 89
rect 1743 55 1783 89
rect 1693 47 1783 55
rect 1813 47 1855 131
rect 1885 47 1955 131
rect 1985 89 2052 131
rect 1985 55 2007 89
rect 2041 55 2052 89
rect 1985 47 2052 55
rect 2082 101 2135 131
rect 2082 67 2093 101
rect 2127 67 2135 101
rect 2082 47 2135 67
rect 2216 127 2224 161
rect 2258 127 2268 161
rect 2216 93 2268 127
rect 2216 59 2224 93
rect 2258 59 2268 93
rect 2216 47 2268 59
rect 2298 161 2352 177
rect 2298 127 2308 161
rect 2342 127 2352 161
rect 2298 93 2352 127
rect 2298 59 2308 93
rect 2342 59 2352 93
rect 2298 47 2352 59
rect 2382 161 2447 177
rect 2382 127 2405 161
rect 2439 127 2447 161
rect 2598 131 2648 177
rect 2382 93 2447 127
rect 2382 59 2405 93
rect 2439 59 2447 93
rect 2382 47 2447 59
rect 2501 105 2553 131
rect 2501 71 2509 105
rect 2543 71 2553 105
rect 2501 47 2553 71
rect 2583 89 2648 131
rect 2583 55 2598 89
rect 2632 55 2648 89
rect 2583 47 2648 55
rect 2678 105 2732 177
rect 2678 71 2688 105
rect 2722 71 2732 105
rect 2678 47 2732 71
rect 2762 161 2824 177
rect 2762 127 2782 161
rect 2816 127 2824 161
rect 2762 93 2824 127
rect 2762 59 2782 93
rect 2816 59 2824 93
rect 2762 47 2824 59
<< pdiff >>
rect 27 431 79 497
rect 27 397 35 431
rect 69 397 79 431
rect 27 369 79 397
rect 109 489 163 497
rect 109 455 119 489
rect 153 455 163 489
rect 109 369 163 455
rect 193 369 235 497
rect 265 411 331 497
rect 265 377 287 411
rect 321 377 331 411
rect 265 369 331 377
rect 361 485 413 497
rect 361 451 371 485
rect 405 451 413 485
rect 361 441 413 451
rect 361 440 412 441
rect 361 369 411 440
rect 467 426 517 497
rect 466 425 517 426
rect 465 415 517 425
rect 465 381 473 415
rect 507 381 517 415
rect 465 369 517 381
rect 547 485 599 497
rect 547 451 557 485
rect 591 451 599 485
rect 547 369 599 451
rect 653 449 705 497
rect 653 415 661 449
rect 695 415 705 449
rect 653 369 705 415
rect 735 489 789 497
rect 735 455 745 489
rect 779 455 789 489
rect 735 369 789 455
rect 819 477 871 497
rect 819 443 829 477
rect 863 443 871 477
rect 819 369 871 443
rect 925 477 977 497
rect 925 443 933 477
rect 967 443 977 477
rect 925 413 977 443
rect 1007 477 1072 497
rect 1007 443 1028 477
rect 1062 443 1072 477
rect 1007 413 1072 443
rect 1102 413 1162 497
rect 1192 489 1281 497
rect 1192 455 1216 489
rect 1250 455 1281 489
rect 1192 413 1281 455
rect 1311 474 1379 497
rect 1311 440 1326 474
rect 1360 440 1379 474
rect 1311 413 1379 440
rect 1409 489 1495 497
rect 1409 455 1428 489
rect 1462 455 1495 489
rect 1409 413 1495 455
rect 1445 329 1495 413
rect 1525 329 1567 497
rect 1597 475 1693 497
rect 1597 441 1637 475
rect 1671 441 1693 475
rect 1597 413 1693 441
rect 1723 413 1781 497
rect 1811 489 1892 497
rect 1811 455 1848 489
rect 1882 455 1892 489
rect 1811 413 1892 455
rect 1922 474 1974 497
rect 1922 440 1932 474
rect 1966 440 1974 474
rect 1922 413 1974 440
rect 2028 485 2080 497
rect 2028 451 2036 485
rect 2070 451 2080 485
rect 2028 413 2080 451
rect 2110 474 2162 497
rect 2110 440 2120 474
rect 2154 440 2162 474
rect 2110 413 2162 440
rect 2216 485 2268 497
rect 2216 451 2224 485
rect 2258 451 2268 485
rect 2216 417 2268 451
rect 1597 329 1647 413
rect 2216 383 2224 417
rect 2258 383 2268 417
rect 2216 349 2268 383
rect 2216 315 2224 349
rect 2258 315 2268 349
rect 2216 297 2268 315
rect 2298 484 2352 497
rect 2298 450 2308 484
rect 2342 450 2352 484
rect 2298 416 2352 450
rect 2298 382 2308 416
rect 2342 382 2352 416
rect 2298 348 2352 382
rect 2298 314 2308 348
rect 2342 314 2352 348
rect 2298 297 2352 314
rect 2382 485 2447 497
rect 2382 451 2405 485
rect 2439 451 2447 485
rect 2598 484 2648 497
rect 2382 417 2447 451
rect 2382 383 2405 417
rect 2439 383 2447 417
rect 2382 349 2447 383
rect 2501 472 2553 484
rect 2501 438 2509 472
rect 2543 438 2553 472
rect 2501 404 2553 438
rect 2501 370 2509 404
rect 2543 370 2553 404
rect 2501 356 2553 370
rect 2583 472 2648 484
rect 2583 438 2603 472
rect 2637 438 2648 472
rect 2583 404 2648 438
rect 2583 370 2603 404
rect 2637 370 2648 404
rect 2583 356 2648 370
rect 2382 315 2405 349
rect 2439 315 2447 349
rect 2382 297 2447 315
rect 2598 297 2648 356
rect 2678 474 2732 497
rect 2678 440 2688 474
rect 2722 440 2732 474
rect 2678 406 2732 440
rect 2678 372 2688 406
rect 2722 372 2732 406
rect 2678 297 2732 372
rect 2762 485 2824 497
rect 2762 451 2782 485
rect 2816 451 2824 485
rect 2762 417 2824 451
rect 2762 383 2782 417
rect 2816 383 2824 417
rect 2762 349 2824 383
rect 2762 315 2782 349
rect 2816 315 2824 349
rect 2762 297 2824 315
<< ndiffc >>
rect 35 69 69 103
rect 191 64 225 98
rect 368 59 402 93
rect 472 71 506 105
rect 556 59 590 93
rect 660 71 694 105
rect 744 55 778 89
rect 828 67 862 101
rect 932 67 966 101
rect 1016 67 1050 101
rect 1172 59 1206 93
rect 1276 85 1310 119
rect 1432 55 1466 89
rect 1709 55 1743 89
rect 2007 55 2041 89
rect 2093 67 2127 101
rect 2224 127 2258 161
rect 2224 59 2258 93
rect 2308 127 2342 161
rect 2308 59 2342 93
rect 2405 127 2439 161
rect 2405 59 2439 93
rect 2509 71 2543 105
rect 2598 55 2632 89
rect 2688 71 2722 105
rect 2782 127 2816 161
rect 2782 59 2816 93
<< pdiffc >>
rect 35 397 69 431
rect 119 455 153 489
rect 287 377 321 411
rect 371 451 405 485
rect 473 381 507 415
rect 557 451 591 485
rect 661 415 695 449
rect 745 455 779 489
rect 829 443 863 477
rect 933 443 967 477
rect 1028 443 1062 477
rect 1216 455 1250 489
rect 1326 440 1360 474
rect 1428 455 1462 489
rect 1637 441 1671 475
rect 1848 455 1882 489
rect 1932 440 1966 474
rect 2036 451 2070 485
rect 2120 440 2154 474
rect 2224 451 2258 485
rect 2224 383 2258 417
rect 2224 315 2258 349
rect 2308 450 2342 484
rect 2308 382 2342 416
rect 2308 314 2342 348
rect 2405 451 2439 485
rect 2405 383 2439 417
rect 2509 438 2543 472
rect 2509 370 2543 404
rect 2603 438 2637 472
rect 2603 370 2637 404
rect 2405 315 2439 349
rect 2688 440 2722 474
rect 2688 372 2722 406
rect 2782 451 2816 485
rect 2782 383 2816 417
rect 2782 315 2816 349
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 235 497 265 523
rect 331 497 361 523
rect 517 497 547 523
rect 705 497 735 523
rect 789 497 819 523
rect 977 497 1007 523
rect 1072 497 1102 523
rect 1162 497 1192 523
rect 1281 497 1311 523
rect 1379 497 1409 523
rect 1495 497 1525 523
rect 1567 497 1597 523
rect 1693 497 1723 523
rect 1781 497 1811 523
rect 1892 497 1922 523
rect 2080 497 2110 523
rect 2268 497 2298 523
rect 2352 497 2382 523
rect 977 398 1007 413
rect 79 354 109 369
rect 48 324 109 354
rect 48 265 78 324
rect 163 283 193 369
rect 21 249 78 265
rect 21 215 34 249
rect 68 215 78 249
rect 120 267 193 283
rect 120 233 130 267
rect 164 253 193 267
rect 164 233 181 253
rect 120 217 181 233
rect 235 219 265 369
rect 331 265 361 369
rect 517 265 547 369
rect 705 354 735 369
rect 683 324 735 354
rect 789 336 819 369
rect 683 284 713 324
rect 777 310 819 336
rect 919 368 1007 398
rect 1072 381 1102 413
rect 1162 381 1192 413
rect 777 284 812 310
rect 919 284 949 368
rect 1049 365 1103 381
rect 1049 331 1059 365
rect 1093 331 1103 365
rect 1049 315 1103 331
rect 1162 365 1239 381
rect 1162 331 1195 365
rect 1229 331 1239 365
rect 1162 315 1239 331
rect 328 249 440 265
rect 21 199 78 215
rect 48 176 78 199
rect 48 146 109 176
rect 79 131 109 146
rect 151 131 181 217
rect 223 203 277 219
rect 223 169 233 203
rect 267 169 277 203
rect 223 153 277 169
rect 328 215 396 249
rect 430 215 440 249
rect 328 199 440 215
rect 487 249 547 265
rect 487 215 497 249
rect 531 215 547 249
rect 659 268 713 284
rect 659 234 669 268
rect 703 234 713 268
rect 659 218 713 234
rect 755 268 812 284
rect 755 234 765 268
rect 799 234 812 268
rect 755 218 812 234
rect 854 268 949 284
rect 854 234 864 268
rect 898 248 949 268
rect 898 234 1080 248
rect 854 218 1080 234
rect 1162 219 1192 315
rect 1281 273 1311 413
rect 1379 369 1409 413
rect 1353 353 1409 369
rect 1353 319 1363 353
rect 1397 319 1409 353
rect 1693 381 1723 413
rect 1685 365 1739 381
rect 1685 345 1695 365
rect 1663 331 1695 345
rect 1729 331 1739 365
rect 1353 303 1409 319
rect 1245 263 1311 273
rect 1245 229 1261 263
rect 1295 229 1311 263
rect 1379 273 1409 303
rect 1379 243 1422 273
rect 1495 265 1525 329
rect 1245 219 1311 229
rect 487 199 547 215
rect 235 131 265 153
rect 328 131 358 199
rect 516 131 546 199
rect 683 176 713 218
rect 782 176 812 218
rect 683 146 734 176
rect 782 146 1006 176
rect 1048 172 1080 218
rect 1132 203 1192 219
rect 1048 146 1090 172
rect 704 131 734 146
rect 788 131 818 146
rect 976 131 1006 146
rect 1060 131 1090 146
rect 1132 169 1142 203
rect 1176 169 1192 203
rect 1132 153 1192 169
rect 1281 176 1311 219
rect 1132 131 1162 153
rect 1281 146 1350 176
rect 1320 131 1350 146
rect 1392 131 1422 243
rect 1464 249 1525 265
rect 1464 215 1474 249
rect 1508 215 1525 249
rect 1464 199 1525 215
rect 1567 265 1597 329
rect 1663 315 1739 331
rect 1781 325 1811 413
rect 1892 397 1922 413
rect 1892 367 1985 397
rect 1927 345 1985 367
rect 2080 365 2110 413
rect 1567 249 1621 265
rect 1567 215 1577 249
rect 1611 215 1621 249
rect 1567 199 1621 215
rect 1487 175 1517 199
rect 1663 175 1693 315
rect 1781 295 1885 325
rect 1927 311 1937 345
rect 1971 311 1985 345
rect 2027 355 2110 365
rect 2027 321 2043 355
rect 2077 321 2110 355
rect 2027 311 2110 321
rect 1927 295 1985 311
rect 1759 237 1813 253
rect 1759 203 1769 237
rect 1803 203 1813 237
rect 1759 187 1813 203
rect 1783 131 1813 187
rect 1855 237 1885 295
rect 1855 221 1913 237
rect 1855 187 1869 221
rect 1903 187 1913 221
rect 1855 171 1913 187
rect 1855 131 1885 171
rect 1955 131 1985 295
rect 2052 265 2110 311
rect 2553 484 2583 523
rect 2648 497 2678 523
rect 2732 497 2762 523
rect 2268 265 2298 297
rect 2352 265 2382 297
rect 2553 265 2583 356
rect 2648 265 2678 297
rect 2732 265 2762 297
rect 2052 203 2583 265
rect 2052 169 2062 203
rect 2096 199 2583 203
rect 2625 249 2762 265
rect 2625 215 2635 249
rect 2669 215 2762 249
rect 2625 199 2762 215
rect 2096 169 2106 199
rect 2268 177 2298 199
rect 2352 177 2382 199
rect 2052 153 2106 169
rect 2052 131 2082 153
rect 2553 131 2583 199
rect 2648 177 2678 199
rect 2732 177 2762 199
rect 79 21 109 47
rect 151 21 181 47
rect 235 21 265 47
rect 328 21 358 47
rect 516 21 546 47
rect 704 21 734 47
rect 788 21 818 47
rect 976 21 1006 47
rect 1060 21 1090 47
rect 1132 21 1162 47
rect 1320 21 1350 47
rect 1392 21 1422 47
rect 1487 21 1517 47
rect 1663 21 1693 47
rect 1783 21 1813 47
rect 1855 21 1885 47
rect 1955 21 1985 47
rect 2052 21 2082 47
rect 2268 21 2298 47
rect 2352 21 2382 47
rect 2553 21 2583 47
rect 2648 21 2678 47
rect 2732 21 2762 47
<< polycont >>
rect 34 215 68 249
rect 130 233 164 267
rect 1059 331 1093 365
rect 1195 331 1229 365
rect 233 169 267 203
rect 396 215 430 249
rect 497 215 531 249
rect 669 234 703 268
rect 765 234 799 268
rect 864 234 898 268
rect 1363 319 1397 353
rect 1695 331 1729 365
rect 1261 229 1295 263
rect 1142 169 1176 203
rect 1474 215 1508 249
rect 1577 215 1611 249
rect 1937 311 1971 345
rect 2043 321 2077 355
rect 1769 203 1803 237
rect 1869 187 1903 221
rect 2062 169 2096 203
rect 2635 215 2669 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2852 561
rect 17 431 69 493
rect 103 489 169 527
rect 103 455 119 489
rect 153 455 169 489
rect 203 485 421 493
rect 17 397 35 431
rect 203 451 371 485
rect 405 451 421 485
rect 203 415 237 451
rect 455 417 507 493
rect 541 485 620 527
rect 541 451 557 485
rect 591 451 620 485
rect 729 489 795 527
rect 541 428 620 451
rect 654 449 695 465
rect 729 455 745 489
rect 779 455 795 489
rect 829 477 888 493
rect 69 397 237 415
rect 17 369 237 397
rect 271 411 339 417
rect 271 377 287 411
rect 321 377 339 411
rect 271 369 339 377
rect 17 249 68 335
rect 17 215 34 249
rect 17 153 68 215
rect 108 267 164 335
rect 108 255 130 267
rect 108 221 121 255
rect 155 221 164 233
rect 108 153 164 221
rect 210 203 267 335
rect 210 169 233 203
rect 210 153 267 169
rect 301 323 339 369
rect 301 289 305 323
rect 301 144 339 289
rect 300 141 339 144
rect 396 415 507 417
rect 396 381 473 415
rect 654 415 661 449
rect 863 443 888 477
rect 829 427 888 443
rect 654 400 695 415
rect 396 352 507 381
rect 396 249 447 352
rect 581 323 620 394
rect 654 391 799 400
rect 654 366 765 391
rect 747 357 765 366
rect 430 215 447 249
rect 481 255 547 318
rect 481 221 489 255
rect 523 249 547 255
rect 481 215 497 221
rect 531 215 547 249
rect 581 268 713 323
rect 581 234 669 268
rect 703 234 713 268
rect 396 181 447 215
rect 581 211 713 234
rect 747 268 799 357
rect 747 234 765 268
rect 396 143 506 181
rect 581 145 620 211
rect 747 177 799 234
rect 299 129 339 141
rect 299 119 334 129
rect 17 103 140 119
rect 17 69 35 103
rect 69 69 140 103
rect 17 17 140 69
rect 174 98 334 119
rect 174 64 191 98
rect 225 64 334 98
rect 174 51 334 64
rect 368 93 418 109
rect 402 59 418 93
rect 368 17 418 59
rect 452 105 506 143
rect 654 143 799 177
rect 833 284 888 427
rect 933 477 978 493
rect 967 443 978 477
rect 933 323 978 443
rect 1012 477 1161 493
rect 1012 443 1028 477
rect 1062 443 1161 477
rect 1200 489 1266 527
rect 1200 455 1216 489
rect 1250 455 1266 489
rect 1321 474 1364 490
rect 1012 427 1161 443
rect 1041 357 1052 391
rect 1086 365 1093 391
rect 1041 331 1059 357
rect 933 318 960 323
rect 943 289 960 318
rect 1041 315 1093 331
rect 833 268 898 284
rect 833 255 864 268
rect 833 221 857 255
rect 891 221 898 234
rect 833 218 898 221
rect 452 71 472 105
rect 452 51 506 71
rect 540 93 620 111
rect 540 59 556 93
rect 590 59 620 93
rect 540 17 620 59
rect 654 105 694 143
rect 833 117 867 218
rect 943 184 977 289
rect 1127 279 1161 427
rect 1321 440 1326 474
rect 1360 440 1364 474
rect 1321 421 1364 440
rect 1412 489 1603 527
rect 1412 455 1428 489
rect 1462 455 1603 489
rect 1412 425 1603 455
rect 1637 475 1798 492
rect 1671 441 1798 475
rect 1832 489 1898 527
rect 1832 455 1848 489
rect 1882 455 1898 489
rect 1832 447 1898 455
rect 1932 474 1986 490
rect 1637 425 1798 441
rect 1195 387 1364 421
rect 1764 413 1798 425
rect 1966 440 1986 474
rect 2020 485 2086 527
rect 2020 451 2036 485
rect 2070 451 2086 485
rect 2020 447 2086 451
rect 2120 474 2169 493
rect 1932 413 1986 440
rect 2154 440 2169 474
rect 1195 365 1229 387
rect 1477 357 1512 391
rect 1546 357 1611 391
rect 1195 315 1229 331
rect 1328 323 1363 353
rect 1362 319 1363 323
rect 1397 319 1413 353
rect 1477 341 1611 357
rect 1362 289 1413 319
rect 1028 263 1295 279
rect 1028 255 1261 263
rect 654 71 660 105
rect 654 51 694 71
rect 728 89 788 109
rect 728 55 744 89
rect 778 55 788 89
rect 728 17 788 55
rect 822 101 867 117
rect 822 67 828 101
rect 862 67 867 101
rect 822 51 867 67
rect 901 101 977 184
rect 901 67 932 101
rect 966 67 977 101
rect 901 51 977 67
rect 1011 245 1261 255
rect 1011 101 1090 245
rect 1471 255 1541 265
rect 1295 249 1541 255
rect 1295 229 1474 249
rect 1261 215 1474 229
rect 1508 215 1541 249
rect 1124 169 1142 203
rect 1176 169 1203 203
rect 1261 195 1541 215
rect 1577 249 1611 341
rect 1684 365 1730 381
rect 1764 379 2086 413
rect 1684 331 1695 365
rect 1729 331 1730 365
rect 2021 355 2086 379
rect 1684 255 1730 331
rect 1776 323 1937 345
rect 1776 289 1788 323
rect 1822 311 1937 323
rect 1971 311 1987 345
rect 1822 305 1987 311
rect 2021 321 2043 355
rect 2077 321 2086 355
rect 2021 305 2086 321
rect 1822 289 1823 305
rect 1776 287 1823 289
rect 2120 271 2169 440
rect 2216 485 2258 527
rect 2216 451 2224 485
rect 2216 417 2258 451
rect 2216 383 2224 417
rect 2216 349 2258 383
rect 2216 315 2224 349
rect 2216 297 2258 315
rect 2292 484 2371 493
rect 2292 450 2308 484
rect 2342 450 2371 484
rect 2292 416 2371 450
rect 2292 382 2308 416
rect 2342 382 2371 416
rect 2292 348 2371 382
rect 2292 314 2308 348
rect 2342 314 2371 348
rect 1684 221 1696 255
rect 1684 215 1730 221
rect 1766 237 1817 253
rect 1124 161 1203 169
rect 1577 179 1611 215
rect 1766 203 1769 237
rect 1803 203 1817 237
rect 1766 179 1817 203
rect 1124 127 1310 161
rect 1011 67 1016 101
rect 1050 67 1090 101
rect 1267 119 1310 127
rect 1011 51 1090 67
rect 1133 59 1172 93
rect 1206 59 1233 93
rect 1133 17 1233 59
rect 1267 85 1276 119
rect 1267 51 1310 85
rect 1344 89 1541 161
rect 1577 139 1817 179
rect 1857 237 2182 271
rect 1857 221 1903 237
rect 1857 187 1869 221
rect 1857 171 1903 187
rect 1937 169 2062 203
rect 2096 169 2112 203
rect 1937 103 1971 169
rect 2146 117 2182 237
rect 1344 55 1432 89
rect 1466 55 1541 89
rect 1693 89 1971 103
rect 1693 55 1709 89
rect 1743 55 1971 89
rect 2007 89 2057 109
rect 2041 55 2057 89
rect 1344 17 1541 55
rect 2007 17 2057 55
rect 2093 101 2182 117
rect 2127 67 2182 101
rect 2093 51 2182 67
rect 2224 161 2258 177
rect 2224 93 2258 127
rect 2224 17 2258 59
rect 2292 161 2371 314
rect 2405 485 2463 527
rect 2439 451 2463 485
rect 2405 417 2463 451
rect 2439 383 2463 417
rect 2405 349 2463 383
rect 2439 315 2463 349
rect 2405 297 2463 315
rect 2506 472 2543 493
rect 2506 438 2509 472
rect 2506 404 2543 438
rect 2506 370 2509 404
rect 2506 265 2543 370
rect 2577 472 2648 527
rect 2577 438 2603 472
rect 2637 438 2648 472
rect 2577 404 2648 438
rect 2577 370 2603 404
rect 2637 370 2648 404
rect 2577 327 2648 370
rect 2682 474 2748 490
rect 2682 440 2688 474
rect 2722 440 2748 474
rect 2682 406 2748 440
rect 2682 372 2688 406
rect 2722 372 2748 406
rect 2682 299 2748 372
rect 2506 249 2669 265
rect 2506 215 2635 249
rect 2506 199 2669 215
rect 2292 127 2308 161
rect 2342 127 2371 161
rect 2292 93 2371 127
rect 2292 59 2308 93
rect 2342 59 2371 93
rect 2292 51 2371 59
rect 2405 161 2463 177
rect 2439 127 2463 161
rect 2405 93 2463 127
rect 2439 59 2463 93
rect 2405 17 2463 59
rect 2506 105 2543 199
rect 2703 165 2748 299
rect 2782 485 2835 527
rect 2816 451 2835 485
rect 2782 417 2835 451
rect 2816 383 2835 417
rect 2782 349 2835 383
rect 2816 315 2835 349
rect 2782 297 2835 315
rect 2506 71 2509 105
rect 2506 51 2543 71
rect 2577 89 2648 165
rect 2577 55 2598 89
rect 2632 55 2648 89
rect 2682 105 2748 165
rect 2682 71 2688 105
rect 2722 71 2748 105
rect 2682 55 2748 71
rect 2782 161 2835 177
rect 2816 127 2835 161
rect 2782 93 2835 127
rect 2816 59 2835 93
rect 2577 17 2648 55
rect 2782 17 2835 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2852 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 2605 527 2639 561
rect 2697 527 2731 561
rect 2789 527 2823 561
rect 121 233 130 255
rect 130 233 155 255
rect 121 221 155 233
rect 305 289 339 323
rect 765 357 799 391
rect 489 249 523 255
rect 489 221 497 249
rect 497 221 523 249
rect 1052 365 1086 391
rect 1052 357 1059 365
rect 1059 357 1086 365
rect 960 289 994 323
rect 857 234 864 255
rect 864 234 891 255
rect 857 221 891 234
rect 1512 357 1546 391
rect 1328 289 1362 323
rect 1788 289 1822 323
rect 1696 221 1730 255
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
rect 2697 -17 2731 17
rect 2789 -17 2823 17
<< metal1 >>
rect 0 561 2852 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2852 561
rect 0 496 2852 527
rect 753 391 811 397
rect 753 357 765 391
rect 799 388 811 391
rect 1040 391 1098 397
rect 1040 388 1052 391
rect 799 360 1052 388
rect 799 357 811 360
rect 753 351 811 357
rect 1040 357 1052 360
rect 1086 388 1098 391
rect 1500 391 1558 397
rect 1500 388 1512 391
rect 1086 360 1512 388
rect 1086 357 1098 360
rect 1040 351 1098 357
rect 1500 357 1512 360
rect 1546 357 1558 391
rect 1500 351 1558 357
rect 293 323 351 329
rect 293 289 305 323
rect 339 320 351 323
rect 948 323 1006 329
rect 948 320 960 323
rect 339 292 960 320
rect 339 289 351 292
rect 293 283 351 289
rect 948 289 960 292
rect 994 289 1006 323
rect 948 283 1006 289
rect 1316 323 1374 329
rect 1316 289 1328 323
rect 1362 320 1374 323
rect 1776 323 1834 329
rect 1776 320 1788 323
rect 1362 292 1788 320
rect 1362 289 1374 292
rect 1316 283 1374 289
rect 1776 289 1788 292
rect 1822 289 1834 323
rect 1776 283 1834 289
rect 109 255 167 261
rect 109 221 121 255
rect 155 252 167 255
rect 477 255 535 261
rect 477 252 489 255
rect 155 224 489 252
rect 155 221 167 224
rect 109 215 167 221
rect 477 221 489 224
rect 523 221 535 255
rect 477 215 535 221
rect 845 255 903 261
rect 845 221 857 255
rect 891 252 903 255
rect 1684 255 1742 261
rect 1684 252 1696 255
rect 891 224 1696 252
rect 891 221 903 224
rect 845 215 903 221
rect 1684 221 1696 224
rect 1730 221 1742 255
rect 1684 215 1742 221
rect 0 17 2852 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2852 17
rect 0 -48 2852 -17
<< labels >>
flabel locali s 29 153 63 187 0 FreeSans 200 0 0 0 SCD
port 3 nsew signal input
flabel locali s 581 357 615 391 0 FreeSans 200 0 0 0 CLK
port 1 nsew clock input
flabel locali s 2337 357 2371 391 0 FreeSans 200 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 213 289 247 323 0 FreeSans 200 0 0 0 D
port 2 nsew signal input
flabel locali s 2337 425 2371 459 0 FreeSans 200 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 29 289 63 323 0 FreeSans 200 0 0 0 SCD
port 3 nsew signal input
flabel locali s 2337 289 2371 323 0 FreeSans 200 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 2337 221 2371 255 0 FreeSans 200 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 2337 153 2371 187 0 FreeSans 200 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 2337 85 2371 119 0 FreeSans 200 0 0 0 Q_N
port 11 nsew signal output
flabel locali s 1328 289 1362 323 0 FreeSans 200 0 0 0 SET_B
port 5 nsew signal input
flabel locali s 121 221 155 255 0 FreeSans 200 0 0 0 SCE
port 4 nsew signal input
flabel locali s 213 153 247 187 0 FreeSans 200 0 0 0 D
port 2 nsew signal input
flabel locali s 581 221 615 255 0 FreeSans 200 0 0 0 CLK
port 1 nsew clock input
flabel locali s 581 153 615 187 0 FreeSans 200 0 0 0 CLK
port 1 nsew clock input
flabel locali s 673 221 707 255 0 FreeSans 200 0 0 0 CLK
port 1 nsew clock input
flabel locali s 2709 357 2743 391 0 FreeSans 200 0 0 0 Q
port 10 nsew signal output
flabel locali s 2709 425 2743 459 0 FreeSans 200 0 0 0 Q
port 10 nsew signal output
flabel locali s 2709 221 2743 255 0 FreeSans 200 0 0 0 Q
port 10 nsew signal output
flabel locali s 2709 153 2743 187 0 FreeSans 200 0 0 0 Q
port 10 nsew signal output
flabel locali s 2709 85 2743 119 0 FreeSans 200 0 0 0 Q
port 10 nsew signal output
flabel locali s 2709 289 2743 323 0 FreeSans 200 0 0 0 Q
port 10 nsew signal output
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 sdfsbp_2
flabel comment s 2095 229 2095 229 0 FreeSans 200 0 0 0 no_jumper_check
flabel comment s 1170 290 1170 290 0 FreeSans 200 0 0 0 no_jumper_check
rlabel locali s 481 215 547 318 1 SCE
port 4 nsew signal input
rlabel metal1 s 477 252 535 261 1 SCE
port 4 nsew signal input
rlabel metal1 s 477 215 535 224 1 SCE
port 4 nsew signal input
rlabel metal1 s 109 252 167 261 1 SCE
port 4 nsew signal input
rlabel metal1 s 109 224 535 252 1 SCE
port 4 nsew signal input
rlabel metal1 s 109 215 167 224 1 SCE
port 4 nsew signal input
rlabel locali s 1776 305 1987 345 1 SET_B
port 5 nsew signal input
rlabel locali s 1776 287 1823 305 1 SET_B
port 5 nsew signal input
rlabel metal1 s 1776 320 1834 329 1 SET_B
port 5 nsew signal input
rlabel metal1 s 1776 283 1834 292 1 SET_B
port 5 nsew signal input
rlabel metal1 s 1316 320 1374 329 1 SET_B
port 5 nsew signal input
rlabel metal1 s 1316 292 1834 320 1 SET_B
port 5 nsew signal input
rlabel metal1 s 1316 283 1374 292 1 SET_B
port 5 nsew signal input
rlabel metal1 s 0 -48 2852 48 1 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 2852 592 1 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2852 544
string GDS_END 264324
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 241692
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 2.720 14.260 2.720 
<< end >>
