magic
tech sky130A
magscale 1 2
timestamp 1666199351
<< nwell >>
rect 304 0 636 490
<< pwell >>
rect 147 328 249 462
<< psubdiff >>
rect 173 412 223 436
rect 173 378 181 412
rect 215 378 223 412
rect 173 354 223 378
<< nsubdiff >>
rect 445 412 495 436
rect 445 378 453 412
rect 487 378 495 412
rect 445 354 495 378
<< psubdiffcont >>
rect 181 378 215 412
<< nsubdiffcont >>
rect 453 378 487 412
<< poly >>
rect 44 214 110 230
rect 44 180 60 214
rect 94 212 110 214
rect 94 182 136 212
rect 260 182 332 212
rect 94 180 110 182
rect 44 164 110 180
<< polycont >>
rect 60 180 94 214
<< locali >>
rect 181 412 215 428
rect 181 362 215 378
rect 453 412 487 428
rect 453 362 487 378
rect 181 264 215 280
rect 60 214 94 230
rect 181 214 215 230
rect 453 264 487 280
rect 453 214 487 230
rect 60 164 94 180
rect 165 130 618 164
<< viali >>
rect 181 378 215 412
rect 453 378 487 412
rect 181 230 215 264
rect 453 230 487 264
<< metal1 >>
rect 169 412 227 418
rect 169 378 181 412
rect 215 378 227 412
rect 169 372 227 378
rect 441 412 499 418
rect 441 378 453 412
rect 487 378 499 412
rect 441 372 499 378
rect 184 270 212 372
rect 456 270 484 372
rect 169 264 227 270
rect 169 230 181 264
rect 215 230 227 264
rect 169 224 227 230
rect 441 264 499 270
rect 441 230 453 264
rect 487 230 499 264
rect 441 224 499 230
rect 184 0 212 224
rect 456 0 484 224
use contact_7  contact_7_0
timestamp 1666199351
transform 1 0 441 0 1 214
box 0 0 1 1
use contact_7  contact_7_1
timestamp 1666199351
transform 1 0 169 0 1 214
box 0 0 1 1
use contact_7  contact_7_2
timestamp 1666199351
transform 1 0 169 0 1 362
box 0 0 1 1
use contact_7  contact_7_3
timestamp 1666199351
transform 1 0 441 0 1 362
box 0 0 1 1
use contact_12  contact_12_0
timestamp 1666199351
transform 1 0 44 0 1 164
box 0 0 1 1
use contact_13  contact_13_0
timestamp 1666199351
transform 1 0 445 0 1 354
box 0 0 1 1
use contact_18  contact_18_0
timestamp 1666199351
transform 1 0 173 0 1 354
box 0 0 1 1
use nmos_m1_w0_360_sli_dli_da_p  nmos_m1_w0_360_sli_dli_da_p_0
timestamp 1666199351
transform 0 1 162 -1 0 272
box -26 -26 176 98
use pmos_m1_w1_120_sli_dli_da_p  pmos_m1_w1_120_sli_dli_da_p_0
timestamp 1666199351
transform 0 1 358 -1 0 272
box -59 -54 209 278
<< labels >>
rlabel locali s 391 147 391 147 4 Z
port 2 nsew
rlabel locali s 77 197 77 197 4 A
port 1 nsew
rlabel metal1 s 470 197 470 197 4 vdd
port 3 nsew
rlabel metal1 s 198 197 198 197 4 gnd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 618 395
string GDS_END 13946
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 12504
<< end >>
