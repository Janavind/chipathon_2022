magic
tech sky130B
magscale 1 2
timestamp 1666199351
<< nwell >>
rect -38 261 2062 582
<< pwell >>
rect 1 21 1951 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 331 47 361 177
rect 415 47 445 177
rect 499 47 529 177
rect 583 47 613 177
rect 667 47 697 177
rect 751 47 781 177
rect 835 47 865 177
rect 919 47 949 177
rect 1003 47 1033 177
rect 1087 47 1117 177
rect 1171 47 1201 177
rect 1255 47 1285 177
rect 1339 47 1369 177
rect 1423 47 1453 177
rect 1507 47 1537 177
rect 1591 47 1621 177
rect 1675 47 1705 177
rect 1759 47 1789 177
rect 1843 47 1873 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 331 297 361 497
rect 415 297 445 497
rect 499 297 529 497
rect 583 297 613 497
rect 667 297 697 497
rect 751 297 781 497
rect 835 297 865 497
rect 919 297 949 497
rect 1003 297 1033 497
rect 1087 297 1117 497
rect 1171 297 1201 497
rect 1255 297 1285 497
rect 1339 297 1369 497
rect 1423 297 1453 497
rect 1507 297 1537 497
rect 1591 297 1621 497
rect 1675 297 1705 497
rect 1759 297 1789 497
rect 1843 297 1873 497
<< ndiff >>
rect 27 165 79 177
rect 27 131 35 165
rect 69 131 79 165
rect 27 97 79 131
rect 27 63 35 97
rect 69 63 79 97
rect 27 47 79 63
rect 109 165 163 177
rect 109 131 119 165
rect 153 131 163 165
rect 109 97 163 131
rect 109 63 119 97
rect 153 63 163 97
rect 109 47 163 63
rect 193 97 247 177
rect 193 63 203 97
rect 237 63 247 97
rect 193 47 247 63
rect 277 165 331 177
rect 277 131 287 165
rect 321 131 331 165
rect 277 97 331 131
rect 277 63 287 97
rect 321 63 331 97
rect 277 47 331 63
rect 361 97 415 177
rect 361 63 371 97
rect 405 63 415 97
rect 361 47 415 63
rect 445 165 499 177
rect 445 131 455 165
rect 489 131 499 165
rect 445 97 499 131
rect 445 63 455 97
rect 489 63 499 97
rect 445 47 499 63
rect 529 97 583 177
rect 529 63 539 97
rect 573 63 583 97
rect 529 47 583 63
rect 613 165 667 177
rect 613 131 623 165
rect 657 131 667 165
rect 613 97 667 131
rect 613 63 623 97
rect 657 63 667 97
rect 613 47 667 63
rect 697 97 751 177
rect 697 63 707 97
rect 741 63 751 97
rect 697 47 751 63
rect 781 165 835 177
rect 781 131 791 165
rect 825 131 835 165
rect 781 97 835 131
rect 781 63 791 97
rect 825 63 835 97
rect 781 47 835 63
rect 865 97 919 177
rect 865 63 875 97
rect 909 63 919 97
rect 865 47 919 63
rect 949 165 1003 177
rect 949 131 959 165
rect 993 131 1003 165
rect 949 97 1003 131
rect 949 63 959 97
rect 993 63 1003 97
rect 949 47 1003 63
rect 1033 97 1087 177
rect 1033 63 1043 97
rect 1077 63 1087 97
rect 1033 47 1087 63
rect 1117 165 1171 177
rect 1117 131 1127 165
rect 1161 131 1171 165
rect 1117 97 1171 131
rect 1117 63 1127 97
rect 1161 63 1171 97
rect 1117 47 1171 63
rect 1201 97 1255 177
rect 1201 63 1211 97
rect 1245 63 1255 97
rect 1201 47 1255 63
rect 1285 165 1339 177
rect 1285 131 1295 165
rect 1329 131 1339 165
rect 1285 97 1339 131
rect 1285 63 1295 97
rect 1329 63 1339 97
rect 1285 47 1339 63
rect 1369 97 1423 177
rect 1369 63 1379 97
rect 1413 63 1423 97
rect 1369 47 1423 63
rect 1453 165 1507 177
rect 1453 131 1463 165
rect 1497 131 1507 165
rect 1453 97 1507 131
rect 1453 63 1463 97
rect 1497 63 1507 97
rect 1453 47 1507 63
rect 1537 97 1591 177
rect 1537 63 1547 97
rect 1581 63 1591 97
rect 1537 47 1591 63
rect 1621 165 1675 177
rect 1621 131 1631 165
rect 1665 131 1675 165
rect 1621 97 1675 131
rect 1621 63 1631 97
rect 1665 63 1675 97
rect 1621 47 1675 63
rect 1705 97 1759 177
rect 1705 63 1715 97
rect 1749 63 1759 97
rect 1705 47 1759 63
rect 1789 165 1843 177
rect 1789 131 1799 165
rect 1833 131 1843 165
rect 1789 97 1843 131
rect 1789 63 1799 97
rect 1833 63 1843 97
rect 1789 47 1843 63
rect 1873 97 1925 177
rect 1873 63 1883 97
rect 1917 63 1925 97
rect 1873 47 1925 63
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 349 79 383
rect 27 315 35 349
rect 69 315 79 349
rect 27 297 79 315
rect 109 479 163 497
rect 109 445 119 479
rect 153 445 163 479
rect 109 411 163 445
rect 109 377 119 411
rect 153 377 163 411
rect 109 343 163 377
rect 109 309 119 343
rect 153 309 163 343
rect 109 297 163 309
rect 193 485 247 497
rect 193 451 203 485
rect 237 451 247 485
rect 193 417 247 451
rect 193 383 203 417
rect 237 383 247 417
rect 193 297 247 383
rect 277 479 331 497
rect 277 445 287 479
rect 321 445 331 479
rect 277 411 331 445
rect 277 377 287 411
rect 321 377 331 411
rect 277 343 331 377
rect 277 309 287 343
rect 321 309 331 343
rect 277 297 331 309
rect 361 485 415 497
rect 361 451 371 485
rect 405 451 415 485
rect 361 417 415 451
rect 361 383 371 417
rect 405 383 415 417
rect 361 297 415 383
rect 445 479 499 497
rect 445 445 455 479
rect 489 445 499 479
rect 445 411 499 445
rect 445 377 455 411
rect 489 377 499 411
rect 445 343 499 377
rect 445 309 455 343
rect 489 309 499 343
rect 445 297 499 309
rect 529 485 583 497
rect 529 451 539 485
rect 573 451 583 485
rect 529 417 583 451
rect 529 383 539 417
rect 573 383 583 417
rect 529 297 583 383
rect 613 479 667 497
rect 613 445 623 479
rect 657 445 667 479
rect 613 411 667 445
rect 613 377 623 411
rect 657 377 667 411
rect 613 343 667 377
rect 613 309 623 343
rect 657 309 667 343
rect 613 297 667 309
rect 697 485 751 497
rect 697 451 707 485
rect 741 451 751 485
rect 697 417 751 451
rect 697 383 707 417
rect 741 383 751 417
rect 697 297 751 383
rect 781 479 835 497
rect 781 445 791 479
rect 825 445 835 479
rect 781 411 835 445
rect 781 377 791 411
rect 825 377 835 411
rect 781 343 835 377
rect 781 309 791 343
rect 825 309 835 343
rect 781 297 835 309
rect 865 485 919 497
rect 865 451 875 485
rect 909 451 919 485
rect 865 417 919 451
rect 865 383 875 417
rect 909 383 919 417
rect 865 297 919 383
rect 949 479 1003 497
rect 949 445 959 479
rect 993 445 1003 479
rect 949 411 1003 445
rect 949 377 959 411
rect 993 377 1003 411
rect 949 343 1003 377
rect 949 309 959 343
rect 993 309 1003 343
rect 949 297 1003 309
rect 1033 485 1087 497
rect 1033 451 1043 485
rect 1077 451 1087 485
rect 1033 417 1087 451
rect 1033 383 1043 417
rect 1077 383 1087 417
rect 1033 297 1087 383
rect 1117 479 1171 497
rect 1117 445 1127 479
rect 1161 445 1171 479
rect 1117 411 1171 445
rect 1117 377 1127 411
rect 1161 377 1171 411
rect 1117 343 1171 377
rect 1117 309 1127 343
rect 1161 309 1171 343
rect 1117 297 1171 309
rect 1201 485 1255 497
rect 1201 451 1211 485
rect 1245 451 1255 485
rect 1201 417 1255 451
rect 1201 383 1211 417
rect 1245 383 1255 417
rect 1201 297 1255 383
rect 1285 479 1339 497
rect 1285 445 1295 479
rect 1329 445 1339 479
rect 1285 411 1339 445
rect 1285 377 1295 411
rect 1329 377 1339 411
rect 1285 343 1339 377
rect 1285 309 1295 343
rect 1329 309 1339 343
rect 1285 297 1339 309
rect 1369 485 1423 497
rect 1369 451 1379 485
rect 1413 451 1423 485
rect 1369 417 1423 451
rect 1369 383 1379 417
rect 1413 383 1423 417
rect 1369 297 1423 383
rect 1453 479 1507 497
rect 1453 445 1463 479
rect 1497 445 1507 479
rect 1453 411 1507 445
rect 1453 377 1463 411
rect 1497 377 1507 411
rect 1453 343 1507 377
rect 1453 309 1463 343
rect 1497 309 1507 343
rect 1453 297 1507 309
rect 1537 485 1591 497
rect 1537 451 1547 485
rect 1581 451 1591 485
rect 1537 417 1591 451
rect 1537 383 1547 417
rect 1581 383 1591 417
rect 1537 297 1591 383
rect 1621 479 1675 497
rect 1621 445 1631 479
rect 1665 445 1675 479
rect 1621 411 1675 445
rect 1621 377 1631 411
rect 1665 377 1675 411
rect 1621 343 1675 377
rect 1621 309 1631 343
rect 1665 309 1675 343
rect 1621 297 1675 309
rect 1705 485 1759 497
rect 1705 451 1715 485
rect 1749 451 1759 485
rect 1705 417 1759 451
rect 1705 383 1715 417
rect 1749 383 1759 417
rect 1705 297 1759 383
rect 1789 479 1843 497
rect 1789 445 1799 479
rect 1833 445 1843 479
rect 1789 411 1843 445
rect 1789 377 1799 411
rect 1833 377 1843 411
rect 1789 343 1843 377
rect 1789 309 1799 343
rect 1833 309 1843 343
rect 1789 297 1843 309
rect 1873 485 1925 497
rect 1873 451 1883 485
rect 1917 451 1925 485
rect 1873 417 1925 451
rect 1873 383 1883 417
rect 1917 383 1925 417
rect 1873 297 1925 383
<< ndiffc >>
rect 35 131 69 165
rect 35 63 69 97
rect 119 131 153 165
rect 119 63 153 97
rect 203 63 237 97
rect 287 131 321 165
rect 287 63 321 97
rect 371 63 405 97
rect 455 131 489 165
rect 455 63 489 97
rect 539 63 573 97
rect 623 131 657 165
rect 623 63 657 97
rect 707 63 741 97
rect 791 131 825 165
rect 791 63 825 97
rect 875 63 909 97
rect 959 131 993 165
rect 959 63 993 97
rect 1043 63 1077 97
rect 1127 131 1161 165
rect 1127 63 1161 97
rect 1211 63 1245 97
rect 1295 131 1329 165
rect 1295 63 1329 97
rect 1379 63 1413 97
rect 1463 131 1497 165
rect 1463 63 1497 97
rect 1547 63 1581 97
rect 1631 131 1665 165
rect 1631 63 1665 97
rect 1715 63 1749 97
rect 1799 131 1833 165
rect 1799 63 1833 97
rect 1883 63 1917 97
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 119 445 153 479
rect 119 377 153 411
rect 119 309 153 343
rect 203 451 237 485
rect 203 383 237 417
rect 287 445 321 479
rect 287 377 321 411
rect 287 309 321 343
rect 371 451 405 485
rect 371 383 405 417
rect 455 445 489 479
rect 455 377 489 411
rect 455 309 489 343
rect 539 451 573 485
rect 539 383 573 417
rect 623 445 657 479
rect 623 377 657 411
rect 623 309 657 343
rect 707 451 741 485
rect 707 383 741 417
rect 791 445 825 479
rect 791 377 825 411
rect 791 309 825 343
rect 875 451 909 485
rect 875 383 909 417
rect 959 445 993 479
rect 959 377 993 411
rect 959 309 993 343
rect 1043 451 1077 485
rect 1043 383 1077 417
rect 1127 445 1161 479
rect 1127 377 1161 411
rect 1127 309 1161 343
rect 1211 451 1245 485
rect 1211 383 1245 417
rect 1295 445 1329 479
rect 1295 377 1329 411
rect 1295 309 1329 343
rect 1379 451 1413 485
rect 1379 383 1413 417
rect 1463 445 1497 479
rect 1463 377 1497 411
rect 1463 309 1497 343
rect 1547 451 1581 485
rect 1547 383 1581 417
rect 1631 445 1665 479
rect 1631 377 1665 411
rect 1631 309 1665 343
rect 1715 451 1749 485
rect 1715 383 1749 417
rect 1799 445 1833 479
rect 1799 377 1833 411
rect 1799 309 1833 343
rect 1883 451 1917 485
rect 1883 383 1917 417
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 331 497 361 523
rect 415 497 445 523
rect 499 497 529 523
rect 583 497 613 523
rect 667 497 697 523
rect 751 497 781 523
rect 835 497 865 523
rect 919 497 949 523
rect 1003 497 1033 523
rect 1087 497 1117 523
rect 1171 497 1201 523
rect 1255 497 1285 523
rect 1339 497 1369 523
rect 1423 497 1453 523
rect 1507 497 1537 523
rect 1591 497 1621 523
rect 1675 497 1705 523
rect 1759 497 1789 523
rect 1843 497 1873 523
rect 79 259 109 297
rect 163 259 193 297
rect 247 259 277 297
rect 331 259 361 297
rect 415 259 445 297
rect 499 259 529 297
rect 79 249 529 259
rect 79 215 103 249
rect 137 215 171 249
rect 205 215 239 249
rect 273 215 307 249
rect 341 215 375 249
rect 409 215 443 249
rect 477 215 529 249
rect 79 205 529 215
rect 79 177 109 205
rect 163 177 193 205
rect 247 177 277 205
rect 331 177 361 205
rect 415 177 445 205
rect 499 177 529 205
rect 583 259 613 297
rect 667 259 697 297
rect 751 259 781 297
rect 835 259 865 297
rect 919 259 949 297
rect 1003 259 1033 297
rect 1087 259 1117 297
rect 1171 259 1201 297
rect 1255 259 1285 297
rect 1339 259 1369 297
rect 1423 259 1453 297
rect 1507 259 1537 297
rect 1591 259 1621 297
rect 1675 259 1705 297
rect 1759 259 1789 297
rect 1843 259 1873 297
rect 583 249 1877 259
rect 583 215 603 249
rect 637 215 671 249
rect 705 215 739 249
rect 773 215 807 249
rect 841 215 875 249
rect 909 215 943 249
rect 977 215 1011 249
rect 1045 215 1079 249
rect 1113 215 1147 249
rect 1181 215 1215 249
rect 1249 215 1283 249
rect 1317 215 1351 249
rect 1385 215 1419 249
rect 1453 215 1487 249
rect 1521 215 1555 249
rect 1589 215 1623 249
rect 1657 215 1691 249
rect 1725 215 1759 249
rect 1793 215 1827 249
rect 1861 215 1877 249
rect 583 205 1877 215
rect 583 177 613 205
rect 667 177 697 205
rect 751 177 781 205
rect 835 177 865 205
rect 919 177 949 205
rect 1003 177 1033 205
rect 1087 177 1117 205
rect 1171 177 1201 205
rect 1255 177 1285 205
rect 1339 177 1369 205
rect 1423 177 1453 205
rect 1507 177 1537 205
rect 1591 177 1621 205
rect 1675 177 1705 205
rect 1759 177 1789 205
rect 1843 177 1873 205
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 331 21 361 47
rect 415 21 445 47
rect 499 21 529 47
rect 583 21 613 47
rect 667 21 697 47
rect 751 21 781 47
rect 835 21 865 47
rect 919 21 949 47
rect 1003 21 1033 47
rect 1087 21 1117 47
rect 1171 21 1201 47
rect 1255 21 1285 47
rect 1339 21 1369 47
rect 1423 21 1453 47
rect 1507 21 1537 47
rect 1591 21 1621 47
rect 1675 21 1705 47
rect 1759 21 1789 47
rect 1843 21 1873 47
<< polycont >>
rect 103 215 137 249
rect 171 215 205 249
rect 239 215 273 249
rect 307 215 341 249
rect 375 215 409 249
rect 443 215 477 249
rect 603 215 637 249
rect 671 215 705 249
rect 739 215 773 249
rect 807 215 841 249
rect 875 215 909 249
rect 943 215 977 249
rect 1011 215 1045 249
rect 1079 215 1113 249
rect 1147 215 1181 249
rect 1215 215 1249 249
rect 1283 215 1317 249
rect 1351 215 1385 249
rect 1419 215 1453 249
rect 1487 215 1521 249
rect 1555 215 1589 249
rect 1623 215 1657 249
rect 1691 215 1725 249
rect 1759 215 1793 249
rect 1827 215 1861 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 35 485 69 527
rect 35 417 69 451
rect 35 349 69 383
rect 35 289 69 315
rect 103 479 169 493
rect 103 445 119 479
rect 153 445 169 479
rect 103 411 169 445
rect 103 377 119 411
rect 153 377 169 411
rect 103 343 169 377
rect 203 485 237 527
rect 203 417 237 451
rect 203 367 237 383
rect 271 479 337 493
rect 271 445 287 479
rect 321 445 337 479
rect 271 411 337 445
rect 271 377 287 411
rect 321 377 337 411
rect 103 309 119 343
rect 153 323 169 343
rect 271 343 337 377
rect 371 485 405 527
rect 371 417 405 451
rect 371 367 405 383
rect 439 479 505 493
rect 439 445 455 479
rect 489 445 505 479
rect 439 411 505 445
rect 439 377 455 411
rect 489 377 505 411
rect 271 323 287 343
rect 153 309 287 323
rect 321 323 337 343
rect 439 343 505 377
rect 539 485 573 527
rect 539 417 573 451
rect 539 367 573 383
rect 607 479 673 493
rect 607 445 623 479
rect 657 445 673 479
rect 607 411 673 445
rect 607 377 623 411
rect 657 377 673 411
rect 439 323 455 343
rect 321 309 455 323
rect 489 323 505 343
rect 607 343 673 377
rect 707 485 741 527
rect 707 417 741 451
rect 707 367 741 383
rect 775 479 841 493
rect 775 445 791 479
rect 825 445 841 479
rect 775 411 841 445
rect 775 377 791 411
rect 825 377 841 411
rect 489 309 573 323
rect 103 289 573 309
rect 607 309 623 343
rect 657 323 673 343
rect 775 343 841 377
rect 875 485 909 527
rect 875 417 909 451
rect 875 367 909 383
rect 943 479 1009 493
rect 943 445 959 479
rect 993 445 1009 479
rect 943 411 1009 445
rect 943 377 959 411
rect 993 377 1009 411
rect 775 323 791 343
rect 657 309 791 323
rect 825 323 841 343
rect 943 343 1009 377
rect 1043 485 1077 527
rect 1043 417 1077 451
rect 1043 367 1077 383
rect 1111 479 1177 493
rect 1111 445 1127 479
rect 1161 445 1177 479
rect 1111 411 1177 445
rect 1111 377 1127 411
rect 1161 377 1177 411
rect 943 323 959 343
rect 825 309 959 323
rect 993 323 1009 343
rect 1111 343 1177 377
rect 1211 485 1245 527
rect 1211 417 1245 451
rect 1211 367 1245 383
rect 1279 479 1345 493
rect 1279 445 1295 479
rect 1329 445 1345 479
rect 1279 411 1345 445
rect 1279 377 1295 411
rect 1329 377 1345 411
rect 1111 323 1127 343
rect 993 309 1127 323
rect 1161 323 1177 343
rect 1279 343 1345 377
rect 1379 485 1413 527
rect 1379 417 1413 451
rect 1379 367 1413 383
rect 1447 479 1513 493
rect 1447 445 1463 479
rect 1497 445 1513 479
rect 1447 411 1513 445
rect 1447 377 1463 411
rect 1497 377 1513 411
rect 1279 323 1295 343
rect 1161 309 1295 323
rect 1329 323 1345 343
rect 1447 343 1513 377
rect 1547 485 1581 527
rect 1547 417 1581 451
rect 1547 367 1581 383
rect 1615 479 1681 493
rect 1615 445 1631 479
rect 1665 445 1681 479
rect 1615 411 1681 445
rect 1615 377 1631 411
rect 1665 377 1681 411
rect 1447 323 1463 343
rect 1329 309 1463 323
rect 1497 323 1513 343
rect 1615 343 1681 377
rect 1715 485 1749 527
rect 1715 417 1749 451
rect 1715 367 1749 383
rect 1783 479 1849 493
rect 1783 445 1799 479
rect 1833 445 1849 479
rect 1783 411 1849 445
rect 1783 377 1799 411
rect 1833 377 1849 411
rect 1615 323 1631 343
rect 1497 309 1631 323
rect 1665 323 1681 343
rect 1783 343 1849 377
rect 1883 485 1917 527
rect 1883 417 1917 451
rect 1883 367 1917 383
rect 1783 323 1799 343
rect 1665 309 1799 323
rect 1833 323 1849 343
rect 1952 323 2007 472
rect 1833 309 2007 323
rect 607 289 2007 309
rect 538 255 573 289
rect 17 249 497 255
rect 17 215 103 249
rect 137 215 171 249
rect 205 215 239 249
rect 273 215 307 249
rect 341 215 375 249
rect 409 215 443 249
rect 477 215 497 249
rect 538 249 1882 255
rect 538 215 603 249
rect 637 215 671 249
rect 705 215 739 249
rect 773 215 807 249
rect 841 215 875 249
rect 909 215 943 249
rect 977 215 1011 249
rect 1045 215 1079 249
rect 1113 215 1147 249
rect 1181 215 1215 249
rect 1249 215 1283 249
rect 1317 215 1351 249
rect 1385 215 1419 249
rect 1453 215 1487 249
rect 1521 215 1555 249
rect 1589 215 1623 249
rect 1657 215 1691 249
rect 1725 215 1759 249
rect 1793 215 1827 249
rect 1861 215 1882 249
rect 538 181 573 215
rect 1931 181 2007 289
rect 35 165 69 181
rect 35 97 69 131
rect 35 17 69 63
rect 103 165 573 181
rect 103 131 119 165
rect 153 147 287 165
rect 153 131 169 147
rect 103 97 169 131
rect 271 131 287 147
rect 321 147 455 165
rect 321 131 337 147
rect 103 63 119 97
rect 153 63 169 97
rect 103 52 169 63
rect 203 97 237 113
rect 203 17 237 63
rect 271 97 337 131
rect 439 131 455 147
rect 489 147 573 165
rect 607 165 2007 181
rect 489 131 505 147
rect 271 63 287 97
rect 321 63 337 97
rect 271 52 337 63
rect 371 97 405 113
rect 371 17 405 63
rect 439 97 505 131
rect 607 131 623 165
rect 657 147 791 165
rect 657 131 673 147
rect 439 63 455 97
rect 489 63 505 97
rect 439 52 505 63
rect 539 97 573 113
rect 539 17 573 63
rect 607 97 673 131
rect 775 131 791 147
rect 825 147 959 165
rect 825 131 841 147
rect 607 63 623 97
rect 657 63 673 97
rect 607 52 673 63
rect 707 97 741 113
rect 607 51 657 52
rect 707 17 741 63
rect 775 97 841 131
rect 943 131 959 147
rect 993 147 1127 165
rect 993 131 1009 147
rect 775 63 791 97
rect 825 63 841 97
rect 775 52 841 63
rect 875 97 909 113
rect 791 51 825 52
rect 875 17 909 63
rect 943 97 1009 131
rect 1111 131 1127 147
rect 1161 147 1295 165
rect 1161 131 1177 147
rect 943 63 959 97
rect 993 63 1009 97
rect 943 52 1009 63
rect 1043 97 1077 113
rect 959 51 993 52
rect 1043 17 1077 63
rect 1111 97 1177 131
rect 1279 131 1295 147
rect 1329 147 1463 165
rect 1329 131 1345 147
rect 1111 63 1127 97
rect 1161 63 1177 97
rect 1111 52 1177 63
rect 1211 97 1245 113
rect 1211 17 1245 63
rect 1279 97 1345 131
rect 1447 131 1463 147
rect 1497 147 1631 165
rect 1497 131 1513 147
rect 1279 63 1295 97
rect 1329 63 1345 97
rect 1279 52 1345 63
rect 1379 97 1413 113
rect 1379 17 1413 63
rect 1447 97 1513 131
rect 1615 131 1631 147
rect 1665 147 1799 165
rect 1665 131 1681 147
rect 1447 63 1463 97
rect 1497 63 1513 97
rect 1447 52 1513 63
rect 1547 97 1581 113
rect 1547 17 1581 63
rect 1615 97 1681 131
rect 1783 131 1799 147
rect 1833 147 2007 165
rect 1833 131 1849 147
rect 1615 63 1631 97
rect 1665 63 1681 97
rect 1615 52 1681 63
rect 1715 97 1749 113
rect 1715 17 1749 63
rect 1783 97 1849 131
rect 1783 63 1799 97
rect 1833 63 1849 97
rect 1783 52 1849 63
rect 1883 97 1917 113
rect 1952 73 2007 147
rect 1883 17 1917 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
<< metal1 >>
rect 0 561 2024 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 0 496 2024 527
rect 0 17 2024 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
rect 0 -48 2024 -17
<< labels >>
flabel locali s 398 221 432 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 306 221 340 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 1961 221 1995 255 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 1961 289 1995 323 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 buf_16
rlabel metal1 s 0 -48 2024 48 1 VGND
port 2 nsew ground bidirectional abutment
rlabel metal1 s 0 496 2024 592 1 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2024 544
string GDS_END 3162694
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3147186
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 13.600 50.600 13.600 
<< end >>
