magic
tech sky130B
magscale 1 2
timestamp 1666464484
<< nwell >>
rect -38 261 1786 582
<< pwell >>
rect 1 201 1433 203
rect 1 23 1744 201
rect 1 21 289 23
rect 747 21 937 23
rect 1348 21 1744 23
rect 30 -17 64 21
<< locali >>
rect 109 288 165 493
rect 109 185 158 288
rect 109 70 161 185
rect 415 215 528 265
rect 1337 289 1453 323
rect 1337 199 1371 289
rect 1501 215 1583 265
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 17 298 75 527
rect 199 443 266 527
rect 302 447 596 481
rect 737 447 803 527
rect 870 455 1489 489
rect 1571 455 1638 527
rect 302 409 336 447
rect 870 413 904 455
rect 199 375 336 409
rect 404 379 904 413
rect 199 265 233 375
rect 279 307 596 341
rect 192 199 233 265
rect 17 17 75 147
rect 198 173 233 199
rect 198 139 313 173
rect 195 17 245 105
rect 279 85 313 139
rect 347 119 381 307
rect 562 265 596 307
rect 630 305 707 339
rect 651 275 707 305
rect 562 199 617 265
rect 441 159 517 181
rect 651 159 685 275
rect 741 241 775 379
rect 821 289 905 343
rect 441 125 685 159
rect 719 207 775 241
rect 719 91 753 207
rect 506 85 593 91
rect 279 51 593 85
rect 627 57 753 91
rect 787 17 821 173
rect 857 83 905 289
rect 941 119 975 421
rect 1009 178 1043 455
rect 1672 421 1731 493
rect 1079 323 1162 409
rect 1269 387 1731 421
rect 1079 289 1235 323
rect 1082 199 1167 254
rect 1009 165 1051 178
rect 1009 144 1091 165
rect 1017 131 1091 144
rect 941 97 983 119
rect 941 53 1023 97
rect 1057 64 1091 131
rect 1125 126 1167 199
rect 1201 85 1235 289
rect 1269 119 1303 387
rect 1634 375 1731 387
rect 1487 299 1651 341
rect 1617 265 1651 299
rect 1405 189 1467 255
rect 1617 199 1663 265
rect 1405 146 1446 189
rect 1617 181 1651 199
rect 1503 150 1651 181
rect 1495 147 1651 150
rect 1337 85 1430 93
rect 1201 51 1430 85
rect 1495 59 1553 147
rect 1697 117 1731 375
rect 1587 17 1621 113
rect 1671 51 1731 117
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
<< metal1 >>
rect 0 561 1748 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 0 496 1748 527
rect 0 17 1748 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
rect 0 -48 1748 -17
<< obsm1 >>
rect 661 320 719 329
rect 1121 320 1179 329
rect 661 292 1179 320
rect 661 283 719 292
rect 1121 283 1179 292
rect 845 184 903 193
rect 1121 184 1179 193
rect 1397 184 1455 193
rect 845 156 1455 184
rect 845 147 903 156
rect 1121 147 1179 156
rect 1397 147 1455 156
rect 937 116 995 125
rect 1489 116 1547 125
rect 937 88 1547 116
rect 937 79 995 88
rect 1489 79 1547 88
<< labels >>
rlabel locali s 1501 215 1583 265 6 A
port 1 nsew signal input
rlabel locali s 1337 199 1371 289 6 B
port 2 nsew signal input
rlabel locali s 1337 289 1453 323 6 B
port 2 nsew signal input
rlabel locali s 415 215 528 265 6 C
port 3 nsew signal input
rlabel metal1 s 0 -48 1748 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1348 21 1744 23 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 747 21 937 23 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 21 289 23 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 23 1744 201 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 201 1433 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 1786 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 1748 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 109 70 161 185 6 X
port 8 nsew signal output
rlabel locali s 109 185 158 288 6 X
port 8 nsew signal output
rlabel locali s 109 288 165 493 6 X
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1748 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 584754
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 572576
<< end >>
