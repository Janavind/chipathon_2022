magic
tech sky130B
magscale 1 2
timestamp 1666464484
<< nwell >>
rect -38 261 1418 582
<< pwell >>
rect 826 157 1379 203
rect 1 21 1379 157
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 351 47 381 131
rect 435 47 465 131
rect 530 47 560 119
rect 621 47 651 119
rect 716 47 746 131
rect 904 47 934 177
rect 988 47 1018 177
rect 1176 47 1206 131
rect 1271 47 1301 177
<< scpmoshvt >>
rect 79 363 109 491
rect 163 363 193 491
rect 353 369 383 497
rect 437 369 467 497
rect 532 413 562 497
rect 618 413 648 497
rect 716 413 746 497
rect 904 297 934 497
rect 988 297 1018 497
rect 1176 369 1206 497
rect 1271 297 1301 497
<< ndiff >>
rect 27 119 79 131
rect 27 85 35 119
rect 69 85 79 119
rect 27 47 79 85
rect 109 93 163 131
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 119 245 131
rect 193 85 203 119
rect 237 85 245 119
rect 193 47 245 85
rect 299 119 351 131
rect 299 85 307 119
rect 341 85 351 119
rect 299 47 351 85
rect 381 89 435 131
rect 381 55 391 89
rect 425 55 435 89
rect 381 47 435 55
rect 465 119 515 131
rect 852 133 904 177
rect 666 119 716 131
rect 465 47 530 119
rect 560 107 621 119
rect 560 73 577 107
rect 611 73 621 107
rect 560 47 621 73
rect 651 47 716 119
rect 746 106 798 131
rect 746 72 756 106
rect 790 72 798 106
rect 746 47 798 72
rect 852 99 860 133
rect 894 99 904 133
rect 852 47 904 99
rect 934 127 988 177
rect 934 93 944 127
rect 978 93 988 127
rect 934 47 988 93
rect 1018 101 1070 177
rect 1221 131 1271 177
rect 1018 67 1028 101
rect 1062 67 1070 101
rect 1018 47 1070 67
rect 1124 119 1176 131
rect 1124 85 1132 119
rect 1166 85 1176 119
rect 1124 47 1176 85
rect 1206 93 1271 131
rect 1206 59 1227 93
rect 1261 59 1271 93
rect 1206 47 1271 59
rect 1301 129 1353 177
rect 1301 95 1311 129
rect 1345 95 1353 129
rect 1301 47 1353 95
<< pdiff >>
rect 27 477 79 491
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 363 79 375
rect 109 461 163 491
rect 109 427 119 461
rect 153 427 163 461
rect 109 363 163 427
rect 193 477 245 491
rect 193 443 203 477
rect 237 443 245 477
rect 193 409 245 443
rect 193 375 203 409
rect 237 375 245 409
rect 193 363 245 375
rect 301 483 353 497
rect 301 449 309 483
rect 343 449 353 483
rect 301 415 353 449
rect 301 381 309 415
rect 343 381 353 415
rect 301 369 353 381
rect 383 485 437 497
rect 383 451 393 485
rect 427 451 437 485
rect 383 417 437 451
rect 383 383 393 417
rect 427 383 437 417
rect 383 369 437 383
rect 467 413 532 497
rect 562 485 618 497
rect 562 451 573 485
rect 607 451 618 485
rect 562 413 618 451
rect 648 413 716 497
rect 746 485 798 497
rect 746 451 756 485
rect 790 451 798 485
rect 746 413 798 451
rect 852 471 904 497
rect 852 437 860 471
rect 894 437 904 471
rect 467 369 517 413
rect 852 368 904 437
rect 852 334 860 368
rect 894 334 904 368
rect 852 297 904 334
rect 934 484 988 497
rect 934 450 944 484
rect 978 450 988 484
rect 934 364 988 450
rect 934 330 944 364
rect 978 330 988 364
rect 934 297 988 330
rect 1018 475 1070 497
rect 1018 441 1028 475
rect 1062 441 1070 475
rect 1018 384 1070 441
rect 1018 350 1028 384
rect 1062 350 1070 384
rect 1124 450 1176 497
rect 1124 416 1132 450
rect 1166 416 1176 450
rect 1124 369 1176 416
rect 1206 485 1271 497
rect 1206 451 1227 485
rect 1261 451 1271 485
rect 1206 417 1271 451
rect 1206 383 1227 417
rect 1261 383 1271 417
rect 1206 369 1271 383
rect 1018 297 1070 350
rect 1221 297 1271 369
rect 1301 449 1353 497
rect 1301 415 1311 449
rect 1345 415 1353 449
rect 1301 381 1353 415
rect 1301 347 1311 381
rect 1345 347 1353 381
rect 1301 297 1353 347
<< ndiffc >>
rect 35 85 69 119
rect 119 59 153 93
rect 203 85 237 119
rect 307 85 341 119
rect 391 55 425 89
rect 577 73 611 107
rect 756 72 790 106
rect 860 99 894 133
rect 944 93 978 127
rect 1028 67 1062 101
rect 1132 85 1166 119
rect 1227 59 1261 93
rect 1311 95 1345 129
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 119 427 153 461
rect 203 443 237 477
rect 203 375 237 409
rect 309 449 343 483
rect 309 381 343 415
rect 393 451 427 485
rect 393 383 427 417
rect 573 451 607 485
rect 756 451 790 485
rect 860 437 894 471
rect 860 334 894 368
rect 944 450 978 484
rect 944 330 978 364
rect 1028 441 1062 475
rect 1028 350 1062 384
rect 1132 416 1166 450
rect 1227 451 1261 485
rect 1227 383 1261 417
rect 1311 415 1345 449
rect 1311 347 1345 381
<< poly >>
rect 79 491 109 517
rect 163 491 193 517
rect 353 497 383 523
rect 437 497 467 523
rect 532 497 562 523
rect 618 497 648 523
rect 716 497 746 523
rect 904 497 934 523
rect 988 497 1018 523
rect 1176 497 1206 523
rect 1271 497 1301 523
rect 79 348 109 363
rect 46 318 109 348
rect 46 280 76 318
rect 21 264 76 280
rect 163 274 193 363
rect 353 338 383 369
rect 21 230 32 264
rect 66 230 76 264
rect 21 214 76 230
rect 118 264 193 274
rect 118 230 134 264
rect 168 230 193 264
rect 301 308 383 338
rect 301 241 331 308
rect 437 247 467 369
rect 532 337 562 413
rect 618 376 648 413
rect 608 366 674 376
rect 509 321 563 337
rect 608 332 624 366
rect 658 332 674 366
rect 608 326 674 332
rect 609 324 674 326
rect 610 322 674 324
rect 716 373 746 413
rect 716 357 808 373
rect 716 323 764 357
rect 798 323 808 357
rect 509 287 519 321
rect 553 299 563 321
rect 716 307 808 323
rect 553 295 570 299
rect 553 288 577 295
rect 553 287 585 288
rect 509 284 585 287
rect 509 283 592 284
rect 509 282 594 283
rect 509 281 597 282
rect 509 280 600 281
rect 509 271 658 280
rect 526 251 658 271
rect 591 250 658 251
rect 594 249 658 250
rect 597 248 658 249
rect 599 247 658 248
rect 118 220 193 230
rect 46 176 76 214
rect 46 146 109 176
rect 79 131 109 146
rect 163 131 193 220
rect 277 225 331 241
rect 277 191 287 225
rect 321 191 331 225
rect 277 176 331 191
rect 417 231 471 247
rect 601 246 658 247
rect 606 243 658 246
rect 611 239 658 243
rect 614 235 658 239
rect 417 197 427 231
rect 461 197 471 231
rect 417 181 471 197
rect 513 207 581 209
rect 513 205 582 207
rect 513 199 583 205
rect 277 175 368 176
rect 299 171 368 175
rect 299 167 373 171
rect 299 161 377 167
rect 299 157 379 161
rect 299 146 381 157
rect 351 131 381 146
rect 435 131 465 181
rect 513 165 533 199
rect 567 165 583 199
rect 513 164 583 165
rect 513 161 582 164
rect 513 158 581 161
rect 513 153 579 158
rect 628 157 658 235
rect 627 156 658 157
rect 625 153 658 156
rect 513 146 560 153
rect 624 151 658 153
rect 623 148 658 151
rect 530 119 560 146
rect 622 145 658 148
rect 621 144 658 145
rect 621 143 657 144
rect 621 142 655 143
rect 621 140 654 142
rect 621 139 653 140
rect 621 137 652 139
rect 621 119 651 137
rect 716 131 746 307
rect 1176 354 1206 369
rect 1170 324 1206 354
rect 904 265 934 297
rect 988 265 1018 297
rect 1170 265 1200 324
rect 1271 265 1301 297
rect 791 249 934 265
rect 791 215 801 249
rect 835 215 934 249
rect 791 199 934 215
rect 986 249 1200 265
rect 986 215 996 249
rect 1030 215 1200 249
rect 986 199 1200 215
rect 1242 249 1301 265
rect 1242 215 1252 249
rect 1286 215 1301 249
rect 1242 199 1301 215
rect 904 177 934 199
rect 988 177 1018 199
rect 1170 176 1200 199
rect 1271 177 1301 199
rect 1170 146 1206 176
rect 1176 131 1206 146
rect 79 21 109 47
rect 163 21 193 47
rect 351 21 381 47
rect 435 21 465 47
rect 530 21 560 47
rect 621 21 651 47
rect 716 21 746 47
rect 904 21 934 47
rect 988 21 1018 47
rect 1176 21 1206 47
rect 1271 21 1301 47
<< polycont >>
rect 32 230 66 264
rect 134 230 168 264
rect 624 332 658 366
rect 764 323 798 357
rect 519 287 553 321
rect 287 191 321 225
rect 427 197 461 231
rect 533 165 567 199
rect 801 215 835 249
rect 996 215 1030 249
rect 1252 215 1286 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 35 477 69 493
rect 35 409 69 443
rect 103 461 169 527
rect 103 427 119 461
rect 153 427 169 461
rect 203 477 248 493
rect 393 485 449 527
rect 756 485 796 527
rect 237 443 248 477
rect 203 409 248 443
rect 69 375 156 393
rect 35 359 156 375
rect 17 264 66 325
rect 17 230 32 264
rect 17 197 66 230
rect 122 323 156 359
rect 122 280 156 289
rect 237 391 248 409
rect 203 357 214 375
rect 203 337 248 357
rect 286 449 309 483
rect 343 449 359 483
rect 286 415 359 449
rect 286 381 309 415
rect 343 381 359 415
rect 122 264 168 280
rect 122 230 134 264
rect 122 214 168 230
rect 122 161 156 214
rect 35 127 156 161
rect 35 119 69 127
rect 203 119 237 337
rect 286 333 359 381
rect 427 451 449 485
rect 550 451 573 485
rect 607 451 722 485
rect 393 417 449 451
rect 427 383 449 417
rect 685 418 722 451
rect 790 451 796 485
rect 756 435 796 451
rect 857 471 903 487
rect 857 437 860 471
rect 894 437 903 471
rect 685 413 726 418
rect 685 407 730 413
rect 686 404 730 407
rect 687 402 730 404
rect 688 399 730 402
rect 393 367 449 383
rect 593 391 639 399
rect 627 382 639 391
rect 627 366 658 382
rect 286 299 423 333
rect 271 225 337 265
rect 271 191 287 225
rect 321 191 337 225
rect 371 247 423 299
rect 493 323 559 337
rect 493 289 511 323
rect 545 321 559 323
rect 493 287 519 289
rect 553 287 559 321
rect 493 271 559 287
rect 593 332 624 357
rect 593 315 658 332
rect 371 231 467 247
rect 371 197 427 231
rect 461 197 467 231
rect 593 213 627 315
rect 692 265 730 399
rect 857 373 903 437
rect 764 368 903 373
rect 764 357 860 368
rect 798 334 860 357
rect 894 334 903 368
rect 798 323 903 334
rect 764 307 903 323
rect 937 484 994 527
rect 937 450 944 484
rect 978 450 994 484
rect 937 364 994 450
rect 937 330 944 364
rect 978 330 994 364
rect 1028 475 1098 491
rect 1062 441 1098 475
rect 1028 384 1098 441
rect 1062 350 1098 384
rect 1028 334 1098 350
rect 937 314 994 330
rect 869 265 903 307
rect 692 249 835 265
rect 692 233 801 249
rect 371 175 467 197
rect 516 199 627 213
rect 371 157 427 175
rect 35 69 69 85
rect 103 59 119 93
rect 153 59 169 93
rect 203 69 237 85
rect 302 123 427 157
rect 516 165 533 199
rect 567 165 627 199
rect 516 141 627 165
rect 661 215 801 233
rect 661 199 835 215
rect 869 249 1030 265
rect 869 215 996 249
rect 869 199 1030 215
rect 302 119 341 123
rect 302 85 307 119
rect 661 107 695 199
rect 869 149 910 199
rect 1064 164 1098 334
rect 302 69 341 85
rect 103 17 169 59
rect 375 55 391 89
rect 425 55 441 89
rect 560 73 577 107
rect 611 73 695 107
rect 857 133 910 149
rect 375 17 441 55
rect 740 72 756 106
rect 790 72 809 106
rect 857 99 860 133
rect 894 99 910 133
rect 857 83 910 99
rect 944 127 994 143
rect 978 93 994 127
rect 740 17 809 72
rect 944 17 994 93
rect 1028 101 1098 164
rect 1062 67 1098 101
rect 1028 51 1098 67
rect 1132 450 1182 493
rect 1166 416 1182 450
rect 1132 265 1182 416
rect 1218 485 1277 527
rect 1218 451 1227 485
rect 1261 451 1277 485
rect 1218 417 1277 451
rect 1218 383 1227 417
rect 1261 383 1277 417
rect 1218 367 1277 383
rect 1311 449 1363 493
rect 1345 415 1363 449
rect 1311 381 1363 415
rect 1345 347 1363 381
rect 1311 289 1363 347
rect 1132 249 1286 265
rect 1132 215 1252 249
rect 1132 199 1286 215
rect 1132 119 1182 199
rect 1320 165 1363 289
rect 1166 85 1182 119
rect 1311 129 1363 165
rect 1132 51 1182 85
rect 1218 93 1277 109
rect 1218 59 1227 93
rect 1261 59 1277 93
rect 1218 17 1277 59
rect 1345 95 1363 129
rect 1311 51 1363 95
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 122 289 156 323
rect 214 375 237 391
rect 237 375 248 391
rect 214 357 248 375
rect 593 366 627 391
rect 593 357 624 366
rect 624 357 627 366
rect 511 321 545 323
rect 511 289 519 321
rect 519 289 545 321
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
<< metal1 >>
rect 0 561 1380 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 0 496 1380 527
rect 202 391 260 397
rect 202 357 214 391
rect 248 388 260 391
rect 581 391 639 397
rect 581 388 593 391
rect 248 360 593 388
rect 248 357 260 360
rect 202 351 260 357
rect 581 357 593 360
rect 627 357 639 391
rect 581 351 639 357
rect 110 323 168 329
rect 110 289 122 323
rect 156 320 168 323
rect 499 323 557 329
rect 499 320 511 323
rect 156 292 511 320
rect 156 289 168 292
rect 110 283 168 289
rect 499 289 511 292
rect 545 289 557 323
rect 499 283 557 289
rect 0 17 1380 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
rect 0 -48 1380 -17
<< labels >>
flabel locali s 289 221 323 255 0 FreeSans 200 0 0 0 D
port 1 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 GATE
port 2 nsew clock input
flabel locali s 1039 357 1073 391 0 FreeSans 200 0 0 0 Q
port 7 nsew signal output
flabel locali s 30 289 64 323 0 FreeSans 200 0 0 0 GATE
port 2 nsew clock input
flabel locali s 1039 425 1073 459 0 FreeSans 200 0 0 0 Q
port 7 nsew signal output
flabel locali s 1039 85 1073 119 0 FreeSans 200 0 0 0 Q
port 7 nsew signal output
flabel locali s 1319 425 1353 459 0 FreeSans 200 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 1319 357 1353 391 0 FreeSans 200 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 1319 85 1353 119 0 FreeSans 200 0 0 0 Q_N
port 8 nsew signal output
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel nwell s 47 544 47 544 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel pwell s 47 0 47 0 0 FreeSans 200 0 0 0 VNB
port 4 nsew
rlabel comment s 0 0 0 0 4 dlxbp_1
rlabel metal1 s 0 -48 1380 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1380 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1380 544
string GDS_END 2849306
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2836820
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 34.500 0.000 
<< end >>
