magic
tech sky130B
magscale 1 2
timestamp 1666464484
<< pwell >>
rect -26 -26 326 3026
<< pdiff >>
rect 0 2945 300 3000
rect 0 55 31 2945
rect 269 55 300 2945
rect 0 0 300 55
<< psubdiffcont >>
rect 31 55 269 2945
use sky130_fd_io__gnd2gnd_strap  sky130_fd_io__gnd2gnd_strap_0
timestamp 1666464484
transform 1 0 0 0 1 0
box 0 0 300 3000
<< properties >>
string GDS_END 8041808
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 8041624
<< end >>
