magic
tech sky130B
timestamp 1666199351
<< properties >>
string GDS_END 29892360
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 29891972
<< end >>
