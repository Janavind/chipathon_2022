magic
tech sky130B
magscale 1 2
timestamp 1668728499
<< viali >>
rect 4721 47209 4755 47243
rect 5365 47209 5399 47243
rect 6009 47209 6043 47243
rect 7113 47209 7147 47243
rect 7757 47209 7791 47243
rect 8401 47209 8435 47243
rect 9137 47209 9171 47243
rect 10241 47209 10275 47243
rect 11161 47209 11195 47243
rect 12449 47209 12483 47243
rect 13553 47209 13587 47243
rect 14657 47209 14691 47243
rect 15669 47209 15703 47243
rect 16313 47209 16347 47243
rect 18889 47209 18923 47243
rect 27169 47209 27203 47243
rect 38485 47209 38519 47243
rect 42625 47209 42659 47243
rect 43269 47209 43303 47243
rect 43913 47209 43947 47243
rect 45201 47209 45235 47243
rect 45845 47209 45879 47243
rect 46489 47209 46523 47243
rect 18245 47141 18279 47175
rect 19533 47141 19567 47175
rect 25973 47141 26007 47175
rect 28917 47141 28951 47175
rect 30205 47141 30239 47175
rect 36369 47141 36403 47175
rect 41337 47141 41371 47175
rect 17601 47073 17635 47107
rect 21465 47073 21499 47107
rect 23581 47073 23615 47107
rect 23857 47073 23891 47107
rect 27905 47073 27939 47107
rect 36001 47073 36035 47107
rect 37933 47073 37967 47107
rect 41981 47073 42015 47107
rect 19441 47005 19475 47039
rect 19963 47005 19997 47039
rect 21189 47005 21223 47039
rect 21373 47005 21407 47039
rect 22293 47005 22327 47039
rect 22477 47005 22511 47039
rect 23673 47005 23707 47039
rect 23765 47005 23799 47039
rect 24041 47005 24075 47039
rect 24869 47005 24903 47039
rect 25053 47005 25087 47039
rect 25789 47005 25823 47039
rect 26065 47005 26099 47039
rect 28089 47005 28123 47039
rect 28457 47005 28491 47039
rect 30021 47005 30055 47039
rect 30297 47005 30331 47039
rect 30941 47005 30975 47039
rect 31769 47005 31803 47039
rect 33888 47005 33922 47039
rect 35173 47005 35207 47039
rect 36185 47005 36219 47039
rect 36461 47005 36495 47039
rect 37749 47005 37783 47039
rect 38025 47005 38059 47039
rect 39129 47005 39163 47039
rect 40049 47005 40083 47039
rect 40693 47005 40727 47039
rect 23397 46937 23431 46971
rect 24685 46937 24719 46971
rect 25605 46937 25639 46971
rect 28365 46937 28399 46971
rect 30757 46937 30791 46971
rect 31125 46937 31159 46971
rect 32321 46937 32355 46971
rect 32505 46937 32539 46971
rect 32873 46937 32907 46971
rect 33517 46937 33551 46971
rect 34989 46937 35023 46971
rect 35449 46937 35483 46971
rect 37565 46937 37599 46971
rect 44557 46937 44591 46971
rect 16957 46869 16991 46903
rect 19901 46869 19935 46903
rect 20085 46869 20119 46903
rect 22109 46869 22143 46903
rect 26617 46869 26651 46903
rect 29837 46869 29871 46903
rect 31677 46869 31711 46903
rect 32597 46869 32631 46903
rect 32689 46869 32723 46903
rect 33425 46869 33459 46903
rect 33609 46869 33643 46903
rect 33701 46869 33735 46903
rect 35357 46869 35391 46903
rect 17877 46665 17911 46699
rect 21189 46665 21223 46699
rect 25973 46665 26007 46699
rect 26157 46665 26191 46699
rect 29285 46665 29319 46699
rect 30205 46665 30239 46699
rect 32505 46665 32539 46699
rect 34437 46665 34471 46699
rect 34621 46665 34655 46699
rect 23857 46597 23891 46631
rect 27261 46597 27295 46631
rect 28181 46597 28215 46631
rect 31585 46597 31619 46631
rect 38577 46597 38611 46631
rect 6929 46529 6963 46563
rect 17417 46529 17451 46563
rect 18061 46529 18095 46563
rect 18521 46529 18555 46563
rect 20085 46529 20119 46563
rect 21251 46529 21285 46563
rect 22477 46529 22511 46563
rect 22569 46529 22603 46563
rect 24041 46529 24075 46563
rect 24410 46529 24444 46563
rect 24593 46529 24627 46563
rect 25237 46529 25271 46563
rect 25421 46529 25455 46563
rect 26155 46529 26189 46563
rect 27721 46529 27755 46563
rect 28365 46529 28399 46563
rect 29009 46529 29043 46563
rect 29285 46529 29319 46563
rect 29515 46529 29549 46563
rect 30665 46529 30699 46563
rect 31769 46529 31803 46563
rect 32505 46529 32539 46563
rect 34439 46529 34473 46563
rect 35817 46529 35851 46563
rect 36369 46529 36403 46563
rect 36553 46529 36587 46563
rect 38025 46529 38059 46563
rect 38761 46529 38795 46563
rect 39037 46529 39071 46563
rect 41429 46529 41463 46563
rect 42625 46529 42659 46563
rect 43729 46529 43763 46563
rect 44465 46529 44499 46563
rect 19349 46461 19383 46495
rect 20269 46461 20303 46495
rect 20729 46461 20763 46495
rect 22845 46461 22879 46495
rect 24225 46461 24259 46495
rect 24317 46461 24351 46495
rect 26617 46461 26651 46495
rect 27445 46461 27479 46495
rect 30113 46461 30147 46495
rect 30297 46461 30331 46495
rect 30941 46461 30975 46495
rect 31401 46461 31435 46495
rect 32321 46461 32355 46495
rect 32873 46461 32907 46495
rect 33977 46461 34011 46495
rect 35173 46461 35207 46495
rect 36001 46461 36035 46495
rect 37749 46461 37783 46495
rect 38945 46461 38979 46495
rect 40785 46461 40819 46495
rect 18705 46393 18739 46427
rect 20821 46393 20855 46427
rect 22293 46393 22327 46427
rect 22753 46393 22787 46427
rect 25053 46393 25087 46427
rect 27629 46393 27663 46427
rect 35909 46393 35943 46427
rect 37933 46393 37967 46427
rect 40141 46393 40175 46427
rect 19901 46325 19935 46359
rect 21373 46325 21407 46359
rect 23397 46325 23431 46359
rect 26525 46325 26559 46359
rect 28457 46325 28491 46359
rect 33333 46325 33367 46359
rect 34069 46325 34103 46359
rect 37565 46325 37599 46359
rect 39497 46325 39531 46359
rect 17509 46121 17543 46155
rect 19717 46121 19751 46155
rect 20637 46121 20671 46155
rect 24777 46121 24811 46155
rect 27353 46121 27387 46155
rect 29837 46121 29871 46155
rect 30849 46121 30883 46155
rect 35541 46121 35575 46155
rect 40693 46121 40727 46155
rect 41337 46121 41371 46155
rect 41981 46121 42015 46155
rect 43821 46121 43855 46155
rect 18245 46053 18279 46087
rect 21465 46053 21499 46087
rect 28921 46053 28955 46087
rect 29009 46053 29043 46087
rect 32965 46053 32999 46087
rect 40049 46053 40083 46087
rect 42625 46053 42659 46087
rect 43177 46053 43211 46087
rect 23397 45985 23431 46019
rect 25513 45985 25547 46019
rect 36553 45985 36587 46019
rect 37933 45985 37967 46019
rect 38669 45985 38703 46019
rect 18889 45917 18923 45951
rect 19901 45917 19935 45951
rect 20085 45917 20119 45951
rect 20729 45917 20763 45951
rect 21645 45917 21679 45951
rect 21833 45917 21867 45951
rect 22293 45917 22327 45951
rect 22477 45917 22511 45951
rect 22661 45917 22695 45951
rect 22937 45917 22971 45951
rect 23581 45917 23615 45951
rect 25697 45917 25731 45951
rect 25789 45917 25823 45951
rect 26525 45917 26559 45951
rect 26801 45917 26835 45951
rect 27537 45917 27571 45951
rect 27629 45917 27663 45951
rect 27813 45917 27847 45951
rect 27905 45917 27939 45951
rect 28549 45917 28583 45951
rect 28825 45917 28859 45951
rect 29101 45917 29135 45951
rect 30021 45917 30055 45951
rect 31033 45917 31067 45951
rect 32045 45917 32079 45951
rect 32321 45917 32355 45951
rect 33793 45917 33827 45951
rect 33977 45917 34011 45951
rect 34345 45917 34379 45951
rect 34989 45917 35023 45951
rect 35716 45905 35750 45939
rect 35817 45917 35851 45951
rect 36001 45917 36035 45951
rect 36093 45917 36127 45951
rect 37749 45917 37783 45951
rect 38761 45917 38795 45951
rect 39037 45917 39071 45951
rect 39221 45917 39255 45951
rect 20913 45849 20947 45883
rect 23949 45849 23983 45883
rect 26341 45849 26375 45883
rect 30297 45849 30331 45883
rect 31309 45849 31343 45883
rect 31861 45849 31895 45883
rect 33333 45849 33367 45883
rect 18705 45781 18739 45815
rect 23673 45781 23707 45815
rect 23765 45781 23799 45815
rect 25329 45781 25363 45815
rect 26709 45781 26743 45815
rect 30205 45781 30239 45815
rect 31217 45781 31251 45815
rect 32229 45781 32263 45815
rect 32873 45781 32907 45815
rect 33977 45781 34011 45815
rect 37105 45781 37139 45815
rect 20637 45577 20671 45611
rect 20821 45577 20855 45611
rect 23213 45577 23247 45611
rect 24685 45577 24719 45611
rect 24869 45577 24903 45611
rect 24961 45577 24995 45611
rect 26157 45577 26191 45611
rect 26249 45577 26283 45611
rect 32873 45577 32907 45611
rect 38025 45577 38059 45611
rect 19993 45509 20027 45543
rect 24133 45509 24167 45543
rect 24777 45509 24811 45543
rect 25145 45509 25179 45543
rect 27353 45509 27387 45543
rect 30205 45509 30239 45543
rect 33609 45509 33643 45543
rect 34069 45509 34103 45543
rect 38853 45509 38887 45543
rect 19257 45441 19291 45475
rect 19901 45441 19935 45475
rect 20819 45441 20853 45475
rect 22293 45441 22327 45475
rect 23213 45441 23247 45475
rect 23581 45441 23615 45475
rect 25789 45441 25823 45475
rect 27169 45441 27203 45475
rect 28457 45441 28491 45475
rect 28733 45441 28767 45475
rect 29745 45441 29779 45475
rect 31033 45441 31067 45475
rect 32321 45441 32355 45475
rect 32413 45441 32447 45475
rect 32597 45441 32631 45475
rect 32689 45441 32723 45475
rect 33953 45441 33987 45475
rect 35173 45441 35207 45475
rect 36151 45441 36185 45475
rect 36553 45441 36587 45475
rect 37565 45441 37599 45475
rect 37657 45441 37691 45475
rect 37841 45441 37875 45475
rect 39037 45441 39071 45475
rect 39589 45441 39623 45475
rect 21281 45373 21315 45407
rect 22477 45373 22511 45407
rect 23029 45373 23063 45407
rect 25605 45373 25639 45407
rect 26048 45373 26082 45407
rect 26341 45373 26375 45407
rect 28089 45373 28123 45407
rect 31125 45373 31159 45407
rect 33865 45373 33899 45407
rect 34161 45373 34195 45407
rect 36461 45373 36495 45407
rect 37745 45373 37779 45407
rect 38761 45373 38795 45407
rect 19441 45305 19475 45339
rect 21189 45305 21223 45339
rect 27537 45305 27571 45339
rect 40233 45305 40267 45339
rect 40785 45305 40819 45339
rect 41337 45305 41371 45339
rect 18705 45237 18739 45271
rect 22109 45237 22143 45271
rect 33425 45237 33459 45271
rect 34713 45237 34747 45271
rect 34897 45237 34931 45271
rect 36001 45237 36035 45271
rect 41981 45237 42015 45271
rect 42625 45237 42659 45271
rect 18797 45033 18831 45067
rect 21833 45033 21867 45067
rect 25973 45033 26007 45067
rect 27169 45033 27203 45067
rect 29009 45033 29043 45067
rect 30757 45033 30791 45067
rect 31769 45033 31803 45067
rect 34161 45033 34195 45067
rect 34989 45033 35023 45067
rect 38393 45033 38427 45067
rect 40601 45033 40635 45067
rect 41153 45033 41187 45067
rect 41797 45033 41831 45067
rect 23581 44965 23615 44999
rect 25145 44965 25179 44999
rect 29837 44965 29871 44999
rect 39129 44965 39163 44999
rect 33701 44897 33735 44931
rect 36369 44897 36403 44931
rect 36829 44897 36863 44931
rect 37565 44897 37599 44931
rect 19809 44829 19843 44863
rect 20545 44829 20579 44863
rect 20729 44829 20763 44863
rect 22017 44829 22051 44863
rect 22661 44829 22695 44863
rect 22845 44829 22879 44863
rect 24593 44829 24627 44863
rect 24685 44829 24719 44863
rect 24869 44829 24903 44863
rect 24961 44829 24995 44863
rect 25881 44829 25915 44863
rect 27629 44829 27663 44863
rect 27721 44829 27755 44863
rect 28088 44829 28122 44863
rect 28733 44829 28767 44863
rect 29929 44829 29963 44863
rect 30205 44829 30239 44863
rect 31953 44829 31987 44863
rect 32137 44829 32171 44863
rect 32689 44829 32723 44863
rect 35081 44829 35115 44863
rect 35725 44829 35759 44863
rect 35909 44829 35943 44863
rect 36185 44829 36219 44863
rect 37473 44829 37507 44863
rect 23857 44761 23891 44795
rect 28273 44761 28307 44795
rect 29009 44761 29043 44795
rect 29193 44761 29227 44795
rect 40049 44761 40083 44795
rect 19993 44693 20027 44727
rect 20913 44693 20947 44727
rect 22753 44693 22787 44727
rect 23397 44693 23431 44727
rect 26341 44693 26375 44727
rect 19717 44489 19751 44523
rect 20269 44489 20303 44523
rect 21005 44489 21039 44523
rect 23213 44489 23247 44523
rect 25421 44489 25455 44523
rect 28641 44489 28675 44523
rect 32689 44489 32723 44523
rect 36185 44489 36219 44523
rect 37565 44489 37599 44523
rect 38577 44489 38611 44523
rect 40785 44489 40819 44523
rect 22109 44421 22143 44455
rect 26525 44421 26559 44455
rect 28181 44421 28215 44455
rect 30757 44421 30791 44455
rect 33609 44421 33643 44455
rect 33977 44421 34011 44455
rect 36093 44421 36127 44455
rect 39129 44421 39163 44455
rect 39681 44421 39715 44455
rect 40233 44421 40267 44455
rect 20821 44353 20855 44387
rect 23581 44353 23615 44387
rect 23949 44353 23983 44387
rect 25053 44353 25087 44387
rect 25421 44353 25455 44387
rect 26341 44353 26375 44387
rect 26617 44353 26651 44387
rect 27537 44353 27571 44387
rect 27721 44353 27755 44387
rect 27997 44353 28031 44387
rect 29285 44353 29319 44387
rect 29653 44353 29687 44387
rect 32505 44353 32539 44387
rect 33793 44353 33827 44387
rect 34069 44353 34103 44387
rect 34621 44353 34655 44387
rect 34805 44353 34839 44387
rect 35633 44353 35667 44387
rect 36369 44353 36403 44387
rect 37749 44353 37783 44387
rect 38025 44353 38059 44387
rect 25605 44285 25639 44319
rect 30205 44285 30239 44319
rect 30849 44285 30883 44319
rect 31401 44285 31435 44319
rect 32321 44285 32355 44319
rect 37933 44285 37967 44319
rect 22753 44217 22787 44251
rect 26157 44217 26191 44251
rect 36553 44149 36587 44183
rect 22385 43945 22419 43979
rect 23029 43945 23063 43979
rect 28089 43945 28123 43979
rect 29193 43945 29227 43979
rect 29837 43945 29871 43979
rect 30757 43945 30791 43979
rect 31401 43945 31435 43979
rect 32321 43945 32355 43979
rect 33701 43945 33735 43979
rect 34989 43945 35023 43979
rect 35357 43945 35391 43979
rect 36001 43945 36035 43979
rect 36185 43945 36219 43979
rect 36921 43945 36955 43979
rect 38485 43945 38519 43979
rect 39037 43945 39071 43979
rect 40049 43945 40083 43979
rect 40601 43945 40635 43979
rect 23949 43877 23983 43911
rect 37381 43877 37415 43911
rect 38025 43877 38059 43911
rect 24041 43809 24075 43843
rect 25053 43809 25087 43843
rect 25881 43809 25915 43843
rect 26617 43809 26651 43843
rect 27537 43809 27571 43843
rect 30021 43809 30055 43843
rect 34345 43809 34379 43843
rect 23489 43741 23523 43775
rect 23673 43741 23707 43775
rect 26893 43741 26927 43775
rect 28273 43741 28307 43775
rect 28549 43741 28583 43775
rect 30205 43741 30239 43775
rect 30297 43741 30331 43775
rect 32597 43741 32631 43775
rect 33425 43741 33459 43775
rect 33609 43741 33643 43775
rect 35449 43741 35483 43775
rect 20729 43673 20763 43707
rect 28457 43673 28491 43707
rect 32413 43673 32447 43707
rect 36185 43673 36219 43707
rect 36369 43673 36403 43707
rect 21189 43605 21223 43639
rect 21833 43605 21867 43639
rect 22845 43401 22879 43435
rect 24593 43401 24627 43435
rect 26157 43401 26191 43435
rect 27261 43401 27295 43435
rect 28825 43401 28859 43435
rect 29377 43401 29411 43435
rect 29929 43401 29963 43435
rect 32321 43401 32355 43435
rect 32873 43401 32907 43435
rect 35449 43401 35483 43435
rect 36553 43401 36587 43435
rect 37565 43401 37599 43435
rect 38577 43401 38611 43435
rect 39129 43401 39163 43435
rect 34529 43333 34563 43367
rect 34713 43333 34747 43367
rect 35909 43333 35943 43367
rect 38117 43333 38151 43367
rect 24777 43265 24811 43299
rect 25421 43265 25455 43299
rect 27721 43265 27755 43299
rect 30481 43265 30515 43299
rect 31585 43265 31619 43299
rect 33793 43265 33827 43299
rect 34897 43265 34931 43299
rect 23489 43197 23523 43231
rect 24961 43197 24995 43231
rect 28181 43197 28215 43231
rect 24041 43061 24075 43095
rect 27445 43061 27479 43095
rect 39681 43061 39715 43095
rect 24685 42857 24719 42891
rect 25973 42857 26007 42891
rect 26617 42857 26651 42891
rect 27905 42857 27939 42891
rect 29745 42857 29779 42891
rect 30389 42857 30423 42891
rect 31953 42857 31987 42891
rect 32597 42857 32631 42891
rect 33885 42857 33919 42891
rect 36645 42857 36679 42891
rect 29101 42789 29135 42823
rect 23029 42721 23063 42755
rect 24041 42721 24075 42755
rect 25513 42721 25547 42755
rect 27077 42721 27111 42755
rect 30849 42721 30883 42755
rect 31401 42721 31435 42755
rect 33057 42721 33091 42755
rect 34897 42721 34931 42755
rect 35449 42721 35483 42755
rect 37197 42721 37231 42755
rect 24777 42653 24811 42687
rect 24961 42653 24995 42687
rect 28549 42653 28583 42687
rect 36093 42585 36127 42619
rect 24133 42313 24167 42347
rect 25145 42313 25179 42347
rect 25605 42313 25639 42347
rect 26249 42313 26283 42347
rect 28641 42313 28675 42347
rect 29193 42313 29227 42347
rect 29745 42313 29779 42347
rect 30941 42313 30975 42347
rect 32413 42313 32447 42347
rect 33609 42313 33643 42347
rect 34529 42313 34563 42347
rect 35725 42313 35759 42347
rect 36369 42313 36403 42347
rect 27261 42245 27295 42279
rect 30481 42245 30515 42279
rect 31493 42245 31527 42279
rect 33057 42245 33091 42279
rect 34989 42245 35023 42279
rect 27721 41973 27755 42007
rect 25329 41769 25363 41803
rect 26249 41769 26283 41803
rect 27997 41769 28031 41803
rect 29745 41769 29779 41803
rect 30849 41769 30883 41803
rect 26985 41701 27019 41735
rect 28641 41701 28675 41735
rect 30297 41701 30331 41735
rect 28641 41225 28675 41259
rect 22937 6749 22971 6783
rect 25329 6749 25363 6783
rect 25789 6681 25823 6715
rect 23029 6613 23063 6647
rect 25145 6613 25179 6647
rect 20545 6409 20579 6443
rect 27169 6409 27203 6443
rect 23765 6341 23799 6375
rect 24501 6341 24535 6375
rect 25973 6341 26007 6375
rect 22293 6273 22327 6307
rect 22937 6273 22971 6307
rect 23673 6273 23707 6307
rect 24409 6205 24443 6239
rect 25881 6205 25915 6239
rect 26525 6205 26559 6239
rect 24961 6137 24995 6171
rect 22385 6069 22419 6103
rect 23029 6069 23063 6103
rect 19533 5865 19567 5899
rect 24041 5865 24075 5899
rect 25053 5865 25087 5899
rect 21925 5729 21959 5763
rect 22477 5729 22511 5763
rect 22937 5729 22971 5763
rect 25973 5729 26007 5763
rect 20177 5661 20211 5695
rect 21097 5661 21131 5695
rect 24961 5661 24995 5695
rect 26801 5661 26835 5695
rect 27629 5661 27663 5695
rect 28089 5661 28123 5695
rect 28917 5661 28951 5695
rect 22569 5593 22603 5627
rect 26157 5593 26191 5627
rect 26249 5593 26283 5627
rect 21189 5525 21223 5559
rect 26893 5525 26927 5559
rect 27537 5525 27571 5559
rect 28181 5525 28215 5559
rect 20821 5321 20855 5355
rect 23121 5253 23155 5287
rect 24593 5253 24627 5287
rect 27353 5253 27387 5287
rect 28549 5253 28583 5287
rect 19993 5185 20027 5219
rect 20637 5185 20671 5219
rect 25789 5185 25823 5219
rect 26433 5185 26467 5219
rect 29745 5185 29779 5219
rect 21465 5117 21499 5151
rect 23029 5117 23063 5151
rect 24501 5117 24535 5151
rect 25145 5117 25179 5151
rect 27261 5117 27295 5151
rect 28457 5117 28491 5151
rect 29101 5117 29135 5151
rect 22477 5049 22511 5083
rect 23581 5049 23615 5083
rect 27813 5049 27847 5083
rect 19441 4981 19475 5015
rect 20085 4981 20119 5015
rect 29653 4981 29687 5015
rect 27353 4777 27387 4811
rect 19717 4709 19751 4743
rect 22201 4709 22235 4743
rect 20269 4641 20303 4675
rect 21649 4641 21683 4675
rect 23581 4641 23615 4675
rect 25053 4641 25087 4675
rect 25605 4641 25639 4675
rect 26065 4641 26099 4675
rect 28825 4641 28859 4675
rect 29101 4641 29135 4675
rect 16957 4573 16991 4607
rect 18889 4573 18923 4607
rect 26893 4573 26927 4607
rect 20361 4505 20395 4539
rect 20913 4505 20947 4539
rect 21741 4505 21775 4539
rect 23121 4505 23155 4539
rect 23213 4505 23247 4539
rect 25697 4505 25731 4539
rect 29009 4505 29043 4539
rect 26709 4437 26743 4471
rect 23581 4233 23615 4267
rect 25605 4233 25639 4267
rect 22293 4165 22327 4199
rect 24317 4165 24351 4199
rect 27721 4165 27755 4199
rect 29009 4165 29043 4199
rect 29745 4165 29779 4199
rect 19993 4097 20027 4131
rect 20085 4097 20119 4131
rect 23489 4097 23523 4131
rect 25513 4097 25547 4131
rect 29837 4097 29871 4131
rect 19533 4029 19567 4063
rect 22201 4029 22235 4063
rect 22477 4029 22511 4063
rect 24225 4029 24259 4063
rect 24685 4029 24719 4063
rect 27445 4029 27479 4063
rect 27813 4029 27847 4063
rect 29101 4029 29135 4063
rect 18245 3961 18279 3995
rect 21465 3961 21499 3995
rect 26617 3961 26651 3995
rect 28549 3961 28583 3995
rect 15025 3893 15059 3927
rect 16129 3893 16163 3927
rect 17601 3893 17635 3927
rect 18889 3893 18923 3927
rect 20821 3893 20855 3927
rect 30297 3893 30331 3927
rect 18245 3689 18279 3723
rect 23305 3689 23339 3723
rect 26893 3689 26927 3723
rect 28917 3689 28951 3723
rect 29745 3689 29779 3723
rect 16313 3621 16347 3655
rect 17601 3621 17635 3655
rect 20637 3621 20671 3655
rect 33609 3621 33643 3655
rect 37473 3621 37507 3655
rect 15025 3553 15059 3587
rect 16957 3553 16991 3587
rect 21189 3553 21223 3587
rect 21465 3553 21499 3587
rect 22753 3553 22787 3587
rect 25237 3553 25271 3587
rect 25513 3553 25547 3587
rect 28089 3553 28123 3587
rect 31033 3553 31067 3587
rect 35541 3553 35575 3587
rect 4261 3485 4295 3519
rect 5181 3485 5215 3519
rect 6009 3485 6043 3519
rect 6837 3485 6871 3519
rect 7665 3485 7699 3519
rect 8493 3485 8527 3519
rect 9321 3485 9355 3519
rect 10149 3485 10183 3519
rect 10977 3485 11011 3519
rect 11713 3485 11747 3519
rect 12357 3485 12391 3519
rect 13001 3485 13035 3519
rect 13645 3485 13679 3519
rect 15669 3485 15703 3519
rect 18705 3485 18739 3519
rect 19809 3485 19843 3519
rect 23213 3485 23247 3519
rect 24041 3485 24075 3519
rect 26801 3485 26835 3519
rect 30573 3485 30607 3519
rect 31677 3485 31711 3519
rect 32321 3485 32355 3519
rect 32965 3485 32999 3519
rect 34897 3485 34931 3519
rect 36185 3485 36219 3519
rect 36829 3485 36863 3519
rect 38117 3485 38151 3519
rect 38761 3485 38795 3519
rect 40049 3485 40083 3519
rect 40693 3485 40727 3519
rect 41337 3485 41371 3519
rect 41981 3485 42015 3519
rect 42901 3485 42935 3519
rect 43361 3485 43395 3519
rect 45201 3485 45235 3519
rect 45845 3485 45879 3519
rect 46489 3485 46523 3519
rect 47133 3485 47167 3519
rect 47777 3485 47811 3519
rect 18797 3417 18831 3451
rect 21281 3417 21315 3451
rect 25338 3417 25372 3451
rect 28273 3417 28307 3451
rect 28365 3417 28399 3451
rect 19901 3349 19935 3383
rect 23949 3349 23983 3383
rect 30481 3349 30515 3383
rect 20177 3145 20211 3179
rect 18245 3077 18279 3111
rect 20913 3077 20947 3111
rect 23029 3077 23063 3111
rect 24133 3077 24167 3111
rect 24225 3077 24259 3111
rect 25973 3077 26007 3111
rect 27353 3077 27387 3111
rect 28917 3077 28951 3111
rect 29009 3077 29043 3111
rect 30113 3077 30147 3111
rect 31493 3077 31527 3111
rect 15025 3009 15059 3043
rect 17049 3009 17083 3043
rect 18337 3009 18371 3043
rect 19441 3009 19475 3043
rect 20085 3009 20119 3043
rect 22201 3009 22235 3043
rect 31401 3009 31435 3043
rect 34253 3009 34287 3043
rect 4721 2941 4755 2975
rect 7297 2941 7331 2975
rect 9229 2941 9263 2975
rect 16313 2941 16347 2975
rect 17693 2941 17727 2975
rect 20821 2941 20855 2975
rect 21465 2941 21499 2975
rect 22937 2941 22971 2975
rect 23581 2941 23615 2975
rect 24409 2941 24443 2975
rect 25789 2941 25823 2975
rect 26065 2941 26099 2975
rect 27261 2941 27295 2975
rect 27537 2941 27571 2975
rect 28549 2941 28583 2975
rect 29561 2941 29595 2975
rect 30205 2941 30239 2975
rect 33609 2941 33643 2975
rect 35541 2941 35575 2975
rect 38117 2941 38151 2975
rect 39405 2941 39439 2975
rect 41337 2941 41371 2975
rect 43269 2941 43303 2975
rect 45201 2941 45235 2975
rect 4077 2873 4111 2907
rect 5365 2873 5399 2907
rect 10517 2873 10551 2907
rect 12449 2873 12483 2907
rect 13737 2873 13771 2907
rect 15669 2873 15703 2907
rect 19533 2873 19567 2907
rect 22293 2873 22327 2907
rect 30757 2873 30791 2907
rect 32965 2873 32999 2907
rect 34897 2873 34931 2907
rect 36185 2873 36219 2907
rect 2789 2805 2823 2839
rect 3433 2805 3467 2839
rect 6009 2805 6043 2839
rect 7941 2805 7975 2839
rect 8585 2805 8619 2839
rect 9873 2805 9907 2839
rect 11161 2805 11195 2839
rect 13093 2805 13127 2839
rect 14381 2805 14415 2839
rect 18981 2805 19015 2839
rect 32321 2805 32355 2839
rect 37473 2805 37507 2839
rect 38761 2805 38795 2839
rect 40049 2805 40083 2839
rect 40693 2805 40727 2839
rect 42625 2805 42659 2839
rect 43913 2805 43947 2839
rect 44557 2805 44591 2839
rect 45845 2805 45879 2839
rect 46489 2805 46523 2839
rect 47777 2805 47811 2839
rect 15025 2601 15059 2635
rect 19625 2601 19659 2635
rect 23949 2601 23983 2635
rect 26341 2601 26375 2635
rect 29745 2601 29779 2635
rect 30481 2601 30515 2635
rect 31033 2601 31067 2635
rect 32321 2601 32355 2635
rect 5365 2533 5399 2567
rect 7941 2533 7975 2567
rect 9873 2533 9907 2567
rect 12449 2533 12483 2567
rect 15669 2533 15703 2567
rect 20177 2533 20211 2567
rect 34897 2533 34931 2567
rect 37473 2533 37507 2567
rect 40049 2533 40083 2567
rect 43913 2533 43947 2567
rect 46489 2533 46523 2567
rect 2789 2465 2823 2499
rect 7297 2465 7331 2499
rect 8585 2465 8619 2499
rect 11161 2465 11195 2499
rect 13093 2465 13127 2499
rect 17601 2465 17635 2499
rect 20821 2465 20855 2499
rect 22477 2465 22511 2499
rect 22753 2465 22787 2499
rect 24961 2465 24995 2499
rect 27813 2465 27847 2499
rect 28365 2465 28399 2499
rect 33609 2465 33643 2499
rect 36185 2465 36219 2499
rect 38761 2465 38795 2499
rect 40693 2465 40727 2499
rect 42625 2465 42659 2499
rect 45201 2465 45235 2499
rect 2145 2397 2179 2431
rect 3433 2397 3467 2431
rect 4721 2397 4755 2431
rect 6009 2397 6043 2431
rect 10517 2397 10551 2431
rect 13737 2397 13771 2431
rect 16313 2397 16347 2431
rect 18245 2397 18279 2431
rect 18889 2397 18923 2431
rect 20085 2397 20119 2431
rect 23857 2397 23891 2431
rect 29193 2397 29227 2431
rect 30573 2397 30607 2431
rect 32965 2397 32999 2431
rect 35541 2397 35575 2431
rect 38117 2397 38151 2431
rect 41337 2397 41371 2431
rect 43269 2397 43303 2431
rect 45845 2397 45879 2431
rect 47777 2397 47811 2431
rect 18153 2329 18187 2363
rect 20913 2329 20947 2363
rect 21465 2329 21499 2363
rect 22569 2329 22603 2363
rect 24685 2329 24719 2363
rect 24777 2329 24811 2363
rect 27169 2329 27203 2363
rect 27721 2329 27755 2363
rect 29101 2329 29135 2363
<< metal1 >>
rect 28994 47608 29000 47660
rect 29052 47648 29058 47660
rect 32950 47648 32956 47660
rect 29052 47620 32956 47648
rect 29052 47608 29058 47620
rect 32950 47608 32956 47620
rect 33008 47608 33014 47660
rect 19426 47540 19432 47592
rect 19484 47580 19490 47592
rect 20254 47580 20260 47592
rect 19484 47552 20260 47580
rect 19484 47540 19490 47552
rect 20254 47540 20260 47552
rect 20312 47540 20318 47592
rect 21910 47540 21916 47592
rect 21968 47580 21974 47592
rect 22094 47580 22100 47592
rect 21968 47552 22100 47580
rect 21968 47540 21974 47552
rect 22094 47540 22100 47552
rect 22152 47540 22158 47592
rect 26786 47540 26792 47592
rect 26844 47580 26850 47592
rect 28810 47580 28816 47592
rect 26844 47552 28816 47580
rect 26844 47540 26850 47552
rect 28810 47540 28816 47552
rect 28868 47540 28874 47592
rect 33318 47580 33324 47592
rect 31726 47552 33324 47580
rect 19886 47472 19892 47524
rect 19944 47512 19950 47524
rect 31726 47512 31754 47552
rect 33318 47540 33324 47552
rect 33376 47540 33382 47592
rect 19944 47484 31754 47512
rect 19944 47472 19950 47484
rect 34146 47472 34152 47524
rect 34204 47512 34210 47524
rect 37734 47512 37740 47524
rect 34204 47484 37740 47512
rect 34204 47472 34210 47484
rect 37734 47472 37740 47484
rect 37792 47512 37798 47524
rect 38746 47512 38752 47524
rect 37792 47484 38752 47512
rect 37792 47472 37798 47484
rect 38746 47472 38752 47484
rect 38804 47472 38810 47524
rect 38838 47472 38844 47524
rect 38896 47512 38902 47524
rect 40770 47512 40776 47524
rect 38896 47484 40776 47512
rect 38896 47472 38902 47484
rect 40770 47472 40776 47484
rect 40828 47472 40834 47524
rect 18874 47404 18880 47456
rect 18932 47444 18938 47456
rect 23474 47444 23480 47456
rect 18932 47416 23480 47444
rect 18932 47404 18938 47416
rect 23474 47404 23480 47416
rect 23532 47404 23538 47456
rect 24118 47404 24124 47456
rect 24176 47444 24182 47456
rect 30190 47444 30196 47456
rect 24176 47416 30196 47444
rect 24176 47404 24182 47416
rect 30190 47404 30196 47416
rect 30248 47404 30254 47456
rect 35342 47404 35348 47456
rect 35400 47444 35406 47456
rect 39758 47444 39764 47456
rect 35400 47416 39764 47444
rect 35400 47404 35406 47416
rect 39758 47404 39764 47416
rect 39816 47404 39822 47456
rect 1104 47354 48852 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 48852 47354
rect 1104 47280 48852 47302
rect 4706 47240 4712 47252
rect 4667 47212 4712 47240
rect 4706 47200 4712 47212
rect 4764 47200 4770 47252
rect 5353 47243 5411 47249
rect 5353 47209 5365 47243
rect 5399 47240 5411 47243
rect 5810 47240 5816 47252
rect 5399 47212 5816 47240
rect 5399 47209 5411 47212
rect 5353 47203 5411 47209
rect 5810 47200 5816 47212
rect 5868 47200 5874 47252
rect 5994 47240 6000 47252
rect 5955 47212 6000 47240
rect 5994 47200 6000 47212
rect 6052 47200 6058 47252
rect 7098 47240 7104 47252
rect 7059 47212 7104 47240
rect 7098 47200 7104 47212
rect 7156 47200 7162 47252
rect 7742 47240 7748 47252
rect 7703 47212 7748 47240
rect 7742 47200 7748 47212
rect 7800 47200 7806 47252
rect 8386 47240 8392 47252
rect 8347 47212 8392 47240
rect 8386 47200 8392 47212
rect 8444 47200 8450 47252
rect 9122 47240 9128 47252
rect 9083 47212 9128 47240
rect 9122 47200 9128 47212
rect 9180 47200 9186 47252
rect 10226 47240 10232 47252
rect 10187 47212 10232 47240
rect 10226 47200 10232 47212
rect 10284 47200 10290 47252
rect 11146 47240 11152 47252
rect 11107 47212 11152 47240
rect 11146 47200 11152 47212
rect 11204 47200 11210 47252
rect 12434 47200 12440 47252
rect 12492 47240 12498 47252
rect 13538 47240 13544 47252
rect 12492 47212 12537 47240
rect 13499 47212 13544 47240
rect 12492 47200 12498 47212
rect 13538 47200 13544 47212
rect 13596 47200 13602 47252
rect 14642 47240 14648 47252
rect 14603 47212 14648 47240
rect 14642 47200 14648 47212
rect 14700 47200 14706 47252
rect 15654 47240 15660 47252
rect 15615 47212 15660 47240
rect 15654 47200 15660 47212
rect 15712 47200 15718 47252
rect 16301 47243 16359 47249
rect 16301 47209 16313 47243
rect 16347 47240 16359 47243
rect 16850 47240 16856 47252
rect 16347 47212 16856 47240
rect 16347 47209 16359 47212
rect 16301 47203 16359 47209
rect 16850 47200 16856 47212
rect 16908 47200 16914 47252
rect 18874 47240 18880 47252
rect 18835 47212 18880 47240
rect 18874 47200 18880 47212
rect 18932 47200 18938 47252
rect 21266 47240 21272 47252
rect 19352 47212 21272 47240
rect 18233 47175 18291 47181
rect 18233 47141 18245 47175
rect 18279 47172 18291 47175
rect 19352 47172 19380 47212
rect 21266 47200 21272 47212
rect 21324 47200 21330 47252
rect 23952 47212 26188 47240
rect 18279 47144 19380 47172
rect 18279 47141 18291 47144
rect 18233 47135 18291 47141
rect 19426 47132 19432 47184
rect 19484 47172 19490 47184
rect 19521 47175 19579 47181
rect 19521 47172 19533 47175
rect 19484 47144 19533 47172
rect 19484 47132 19490 47144
rect 19521 47141 19533 47144
rect 19567 47172 19579 47175
rect 20530 47172 20536 47184
rect 19567 47144 20536 47172
rect 19567 47141 19579 47144
rect 19521 47135 19579 47141
rect 20530 47132 20536 47144
rect 20588 47132 20594 47184
rect 23106 47172 23112 47184
rect 21284 47144 23112 47172
rect 17589 47107 17647 47113
rect 17589 47073 17601 47107
rect 17635 47104 17647 47107
rect 20162 47104 20168 47116
rect 17635 47076 20168 47104
rect 17635 47073 17647 47076
rect 17589 47067 17647 47073
rect 20162 47064 20168 47076
rect 20220 47064 20226 47116
rect 17862 46996 17868 47048
rect 17920 47036 17926 47048
rect 19429 47039 19487 47045
rect 19429 47036 19441 47039
rect 17920 47008 19441 47036
rect 17920 46996 17926 47008
rect 19429 47005 19441 47008
rect 19475 47005 19487 47039
rect 19429 46999 19487 47005
rect 19951 47039 20009 47045
rect 19951 47005 19963 47039
rect 19997 47036 20009 47039
rect 20346 47036 20352 47048
rect 19997 47008 20352 47036
rect 19997 47005 20009 47008
rect 19951 46999 20009 47005
rect 20346 46996 20352 47008
rect 20404 46996 20410 47048
rect 21177 47039 21235 47045
rect 21177 47005 21189 47039
rect 21223 47036 21235 47039
rect 21284 47036 21312 47144
rect 23106 47132 23112 47144
rect 23164 47132 23170 47184
rect 21453 47107 21511 47113
rect 21453 47073 21465 47107
rect 21499 47104 21511 47107
rect 23569 47107 23627 47113
rect 23569 47104 23581 47107
rect 21499 47076 23581 47104
rect 21499 47073 21511 47076
rect 21453 47067 21511 47073
rect 23569 47073 23581 47076
rect 23615 47073 23627 47107
rect 23842 47104 23848 47116
rect 23803 47076 23848 47104
rect 23569 47067 23627 47073
rect 23842 47064 23848 47076
rect 23900 47064 23906 47116
rect 21223 47008 21312 47036
rect 21361 47039 21419 47045
rect 21223 47005 21235 47008
rect 21177 46999 21235 47005
rect 21361 47005 21373 47039
rect 21407 47036 21419 47039
rect 21407 47008 22094 47036
rect 21407 47005 21419 47008
rect 21361 46999 21419 47005
rect 19334 46928 19340 46980
rect 19392 46968 19398 46980
rect 20162 46968 20168 46980
rect 19392 46940 20168 46968
rect 19392 46928 19398 46940
rect 20162 46928 20168 46940
rect 20220 46928 20226 46980
rect 22066 46968 22094 47008
rect 22186 46996 22192 47048
rect 22244 47036 22250 47048
rect 22281 47039 22339 47045
rect 22281 47036 22293 47039
rect 22244 47008 22293 47036
rect 22244 46996 22250 47008
rect 22281 47005 22293 47008
rect 22327 47005 22339 47039
rect 22462 47036 22468 47048
rect 22423 47008 22468 47036
rect 22281 46999 22339 47005
rect 22462 46996 22468 47008
rect 22520 46996 22526 47048
rect 22738 46996 22744 47048
rect 22796 47036 22802 47048
rect 23661 47039 23719 47045
rect 23661 47036 23673 47039
rect 22796 47008 23673 47036
rect 22796 46996 22802 47008
rect 23661 47005 23673 47008
rect 23707 47005 23719 47039
rect 23661 46999 23719 47005
rect 23753 47039 23811 47045
rect 23753 47005 23765 47039
rect 23799 47036 23811 47039
rect 23952 47036 23980 47212
rect 24026 47132 24032 47184
rect 24084 47172 24090 47184
rect 25958 47172 25964 47184
rect 24084 47144 25636 47172
rect 25919 47144 25964 47172
rect 24084 47132 24090 47144
rect 25498 47104 25504 47116
rect 24872 47076 25504 47104
rect 23799 47008 23980 47036
rect 24029 47039 24087 47045
rect 23799 47005 23811 47008
rect 23753 46999 23811 47005
rect 24029 47005 24041 47039
rect 24075 47036 24087 47039
rect 24118 47036 24124 47048
rect 24075 47008 24124 47036
rect 24075 47005 24087 47008
rect 24029 46999 24087 47005
rect 23198 46968 23204 46980
rect 22066 46940 23204 46968
rect 23198 46928 23204 46940
rect 23256 46928 23262 46980
rect 23382 46968 23388 46980
rect 23343 46940 23388 46968
rect 23382 46928 23388 46940
rect 23440 46928 23446 46980
rect 16942 46900 16948 46912
rect 16903 46872 16948 46900
rect 16942 46860 16948 46872
rect 17000 46860 17006 46912
rect 19886 46900 19892 46912
rect 19847 46872 19892 46900
rect 19886 46860 19892 46872
rect 19944 46860 19950 46912
rect 19978 46860 19984 46912
rect 20036 46900 20042 46912
rect 20073 46903 20131 46909
rect 20073 46900 20085 46903
rect 20036 46872 20085 46900
rect 20036 46860 20042 46872
rect 20073 46869 20085 46872
rect 20119 46869 20131 46903
rect 20073 46863 20131 46869
rect 20438 46860 20444 46912
rect 20496 46900 20502 46912
rect 22097 46903 22155 46909
rect 22097 46900 22109 46903
rect 20496 46872 22109 46900
rect 20496 46860 20502 46872
rect 22097 46869 22109 46872
rect 22143 46869 22155 46903
rect 22097 46863 22155 46869
rect 22278 46860 22284 46912
rect 22336 46900 22342 46912
rect 24044 46900 24072 46999
rect 24118 46996 24124 47008
rect 24176 46996 24182 47048
rect 24872 47045 24900 47076
rect 25498 47064 25504 47076
rect 25556 47064 25562 47116
rect 24857 47039 24915 47045
rect 24857 47005 24869 47039
rect 24903 47005 24915 47039
rect 24857 46999 24915 47005
rect 25041 47039 25099 47045
rect 25041 47005 25053 47039
rect 25087 47036 25099 47039
rect 25222 47036 25228 47048
rect 25087 47008 25228 47036
rect 25087 47005 25099 47008
rect 25041 46999 25099 47005
rect 25222 46996 25228 47008
rect 25280 46996 25286 47048
rect 25608 47036 25636 47144
rect 25958 47132 25964 47144
rect 26016 47132 26022 47184
rect 26160 47172 26188 47212
rect 26234 47200 26240 47252
rect 26292 47240 26298 47252
rect 27157 47243 27215 47249
rect 27157 47240 27169 47243
rect 26292 47212 27169 47240
rect 26292 47200 26298 47212
rect 27157 47209 27169 47212
rect 27203 47209 27215 47243
rect 30834 47240 30840 47252
rect 27157 47203 27215 47209
rect 27632 47212 30840 47240
rect 27632 47172 27660 47212
rect 30834 47200 30840 47212
rect 30892 47200 30898 47252
rect 32674 47200 32680 47252
rect 32732 47240 32738 47252
rect 38473 47243 38531 47249
rect 38473 47240 38485 47243
rect 32732 47212 38485 47240
rect 32732 47200 32738 47212
rect 38473 47209 38485 47212
rect 38519 47209 38531 47243
rect 38473 47203 38531 47209
rect 40678 47200 40684 47252
rect 40736 47240 40742 47252
rect 42613 47243 42671 47249
rect 42613 47240 42625 47243
rect 40736 47212 42625 47240
rect 40736 47200 40742 47212
rect 42613 47209 42625 47212
rect 42659 47209 42671 47243
rect 42613 47203 42671 47209
rect 42794 47200 42800 47252
rect 42852 47240 42858 47252
rect 43257 47243 43315 47249
rect 43257 47240 43269 47243
rect 42852 47212 43269 47240
rect 42852 47200 42858 47212
rect 43257 47209 43269 47212
rect 43303 47209 43315 47243
rect 43257 47203 43315 47209
rect 43346 47200 43352 47252
rect 43404 47240 43410 47252
rect 43901 47243 43959 47249
rect 43901 47240 43913 47243
rect 43404 47212 43913 47240
rect 43404 47200 43410 47212
rect 43901 47209 43913 47212
rect 43947 47209 43959 47243
rect 43901 47203 43959 47209
rect 44818 47200 44824 47252
rect 44876 47240 44882 47252
rect 45189 47243 45247 47249
rect 45189 47240 45201 47243
rect 44876 47212 45201 47240
rect 44876 47200 44882 47212
rect 45189 47209 45201 47212
rect 45235 47209 45247 47243
rect 45830 47240 45836 47252
rect 45791 47212 45836 47240
rect 45189 47203 45247 47209
rect 45830 47200 45836 47212
rect 45888 47200 45894 47252
rect 45922 47200 45928 47252
rect 45980 47240 45986 47252
rect 46477 47243 46535 47249
rect 46477 47240 46489 47243
rect 45980 47212 46489 47240
rect 45980 47200 45986 47212
rect 46477 47209 46489 47212
rect 46523 47209 46535 47243
rect 46477 47203 46535 47209
rect 28350 47172 28356 47184
rect 26160 47144 27660 47172
rect 27724 47144 28356 47172
rect 26142 47104 26148 47116
rect 26055 47076 26148 47104
rect 25777 47039 25835 47045
rect 25608 47008 25728 47036
rect 24670 46968 24676 46980
rect 24631 46940 24676 46968
rect 24670 46928 24676 46940
rect 24728 46928 24734 46980
rect 25590 46968 25596 46980
rect 25551 46940 25596 46968
rect 25590 46928 25596 46940
rect 25648 46928 25654 46980
rect 25700 46968 25728 47008
rect 25777 47005 25789 47039
rect 25823 47036 25835 47039
rect 25866 47036 25872 47048
rect 25823 47008 25872 47036
rect 25823 47005 25835 47008
rect 25777 46999 25835 47005
rect 25866 46996 25872 47008
rect 25924 46996 25930 47048
rect 26068 47045 26096 47076
rect 26142 47064 26148 47076
rect 26200 47104 26206 47116
rect 27724 47104 27752 47144
rect 28350 47132 28356 47144
rect 28408 47172 28414 47184
rect 28718 47172 28724 47184
rect 28408 47144 28724 47172
rect 28408 47132 28414 47144
rect 28718 47132 28724 47144
rect 28776 47132 28782 47184
rect 28810 47132 28816 47184
rect 28868 47172 28874 47184
rect 28905 47175 28963 47181
rect 28905 47172 28917 47175
rect 28868 47144 28917 47172
rect 28868 47132 28874 47144
rect 28905 47141 28917 47144
rect 28951 47141 28963 47175
rect 28905 47135 28963 47141
rect 29914 47132 29920 47184
rect 29972 47172 29978 47184
rect 30193 47175 30251 47181
rect 30193 47172 30205 47175
rect 29972 47144 30205 47172
rect 29972 47132 29978 47144
rect 30193 47141 30205 47144
rect 30239 47141 30251 47175
rect 34606 47172 34612 47184
rect 30193 47135 30251 47141
rect 31726 47144 34612 47172
rect 26200 47076 27752 47104
rect 27893 47107 27951 47113
rect 26200 47064 26206 47076
rect 27893 47073 27905 47107
rect 27939 47104 27951 47107
rect 29086 47104 29092 47116
rect 27939 47076 29092 47104
rect 27939 47073 27951 47076
rect 27893 47067 27951 47073
rect 29086 47064 29092 47076
rect 29144 47064 29150 47116
rect 29730 47064 29736 47116
rect 29788 47104 29794 47116
rect 31726 47104 31754 47144
rect 34606 47132 34612 47144
rect 34664 47132 34670 47184
rect 34698 47132 34704 47184
rect 34756 47172 34762 47184
rect 36357 47175 36415 47181
rect 36357 47172 36369 47175
rect 34756 47144 36369 47172
rect 34756 47132 34762 47144
rect 36357 47141 36369 47144
rect 36403 47141 36415 47175
rect 36357 47135 36415 47141
rect 37090 47132 37096 47184
rect 37148 47172 37154 47184
rect 41325 47175 41383 47181
rect 41325 47172 41337 47175
rect 37148 47144 41337 47172
rect 37148 47132 37154 47144
rect 41325 47141 41337 47144
rect 41371 47141 41383 47175
rect 41325 47135 41383 47141
rect 35989 47107 36047 47113
rect 35989 47104 36001 47107
rect 29788 47076 30328 47104
rect 29788 47064 29794 47076
rect 26053 47039 26111 47045
rect 26053 47005 26065 47039
rect 26099 47005 26111 47039
rect 26053 46999 26111 47005
rect 26418 46996 26424 47048
rect 26476 47036 26482 47048
rect 28077 47039 28135 47045
rect 28077 47036 28089 47039
rect 26476 47008 28089 47036
rect 26476 46996 26482 47008
rect 28077 47005 28089 47008
rect 28123 47036 28135 47039
rect 28166 47036 28172 47048
rect 28123 47008 28172 47036
rect 28123 47005 28135 47008
rect 28077 46999 28135 47005
rect 28166 46996 28172 47008
rect 28224 46996 28230 47048
rect 28442 47036 28448 47048
rect 28403 47008 28448 47036
rect 28442 46996 28448 47008
rect 28500 46996 28506 47048
rect 29362 46996 29368 47048
rect 29420 47036 29426 47048
rect 30300 47045 30328 47076
rect 30392 47076 31800 47104
rect 30009 47039 30067 47045
rect 30009 47036 30021 47039
rect 29420 47008 30021 47036
rect 29420 46996 29426 47008
rect 30009 47005 30021 47008
rect 30055 47005 30067 47039
rect 30009 46999 30067 47005
rect 30285 47039 30343 47045
rect 30285 47005 30297 47039
rect 30331 47005 30343 47039
rect 30285 46999 30343 47005
rect 28353 46971 28411 46977
rect 28353 46968 28365 46971
rect 25700 46940 28365 46968
rect 28353 46937 28365 46940
rect 28399 46937 28411 46971
rect 30392 46968 30420 47076
rect 30558 46996 30564 47048
rect 30616 47036 30622 47048
rect 30929 47039 30987 47045
rect 30616 47008 30880 47036
rect 30616 46996 30622 47008
rect 30742 46968 30748 46980
rect 28353 46931 28411 46937
rect 28460 46940 30420 46968
rect 30703 46940 30748 46968
rect 22336 46872 24072 46900
rect 22336 46860 22342 46872
rect 24210 46860 24216 46912
rect 24268 46900 24274 46912
rect 25958 46900 25964 46912
rect 24268 46872 25964 46900
rect 24268 46860 24274 46872
rect 25958 46860 25964 46872
rect 26016 46860 26022 46912
rect 26234 46860 26240 46912
rect 26292 46900 26298 46912
rect 26605 46903 26663 46909
rect 26605 46900 26617 46903
rect 26292 46872 26617 46900
rect 26292 46860 26298 46872
rect 26605 46869 26617 46872
rect 26651 46900 26663 46903
rect 27706 46900 27712 46912
rect 26651 46872 27712 46900
rect 26651 46869 26663 46872
rect 26605 46863 26663 46869
rect 27706 46860 27712 46872
rect 27764 46900 27770 46912
rect 28460 46900 28488 46940
rect 30300 46912 30328 46940
rect 30742 46928 30748 46940
rect 30800 46928 30806 46980
rect 30852 46968 30880 47008
rect 30929 47005 30941 47039
rect 30975 47036 30987 47039
rect 31018 47036 31024 47048
rect 30975 47008 31024 47036
rect 30975 47005 30987 47008
rect 30929 46999 30987 47005
rect 31018 46996 31024 47008
rect 31076 46996 31082 47048
rect 31772 47045 31800 47076
rect 33980 47076 36001 47104
rect 31757 47039 31815 47045
rect 31757 47005 31769 47039
rect 31803 47005 31815 47039
rect 33594 47036 33600 47048
rect 31757 46999 31815 47005
rect 32968 47008 33600 47036
rect 31113 46971 31171 46977
rect 31113 46968 31125 46971
rect 30852 46940 31125 46968
rect 31113 46937 31125 46940
rect 31159 46968 31171 46971
rect 32309 46971 32367 46977
rect 32309 46968 32321 46971
rect 31159 46940 32321 46968
rect 31159 46937 31171 46940
rect 31113 46931 31171 46937
rect 32309 46937 32321 46940
rect 32355 46937 32367 46971
rect 32309 46931 32367 46937
rect 32398 46928 32404 46980
rect 32456 46968 32462 46980
rect 32493 46971 32551 46977
rect 32493 46968 32505 46971
rect 32456 46940 32505 46968
rect 32456 46928 32462 46940
rect 32493 46937 32505 46940
rect 32539 46937 32551 46971
rect 32493 46931 32551 46937
rect 32861 46971 32919 46977
rect 32861 46937 32873 46971
rect 32907 46968 32919 46971
rect 32968 46968 32996 47008
rect 33594 46996 33600 47008
rect 33652 46996 33658 47048
rect 33876 47039 33934 47045
rect 33876 47005 33888 47039
rect 33922 47038 33934 47039
rect 33980 47038 34008 47076
rect 35989 47073 36001 47076
rect 36035 47073 36047 47107
rect 35989 47067 36047 47073
rect 36538 47064 36544 47116
rect 36596 47104 36602 47116
rect 37921 47107 37979 47113
rect 37921 47104 37933 47107
rect 36596 47076 37933 47104
rect 36596 47064 36602 47076
rect 37921 47073 37933 47076
rect 37967 47104 37979 47107
rect 37967 47076 38700 47104
rect 37967 47073 37979 47076
rect 37921 47067 37979 47073
rect 33922 47010 34008 47038
rect 35158 47036 35164 47048
rect 33922 47005 33934 47010
rect 35119 47008 35164 47036
rect 33876 46999 33934 47005
rect 35158 46996 35164 47008
rect 35216 46996 35222 47048
rect 35250 46996 35256 47048
rect 35308 47036 35314 47048
rect 36173 47039 36231 47045
rect 36173 47036 36185 47039
rect 35308 47008 36185 47036
rect 35308 46996 35314 47008
rect 36173 47005 36185 47008
rect 36219 47005 36231 47039
rect 36173 46999 36231 47005
rect 36449 47039 36507 47045
rect 36449 47005 36461 47039
rect 36495 47036 36507 47039
rect 37274 47036 37280 47048
rect 36495 47008 37280 47036
rect 36495 47005 36507 47008
rect 36449 46999 36507 47005
rect 37274 46996 37280 47008
rect 37332 46996 37338 47048
rect 37734 47036 37740 47048
rect 37695 47008 37740 47036
rect 37734 46996 37740 47008
rect 37792 46996 37798 47048
rect 38013 47039 38071 47045
rect 38013 47005 38025 47039
rect 38059 47036 38071 47039
rect 38562 47036 38568 47048
rect 38059 47008 38568 47036
rect 38059 47005 38071 47008
rect 38013 46999 38071 47005
rect 32907 46940 32996 46968
rect 32907 46937 32919 46940
rect 32861 46931 32919 46937
rect 33226 46928 33232 46980
rect 33284 46968 33290 46980
rect 33505 46971 33563 46977
rect 33505 46968 33517 46971
rect 33284 46940 33517 46968
rect 33284 46928 33290 46940
rect 33505 46937 33517 46940
rect 33551 46968 33563 46971
rect 33551 46940 34008 46968
rect 33551 46937 33563 46940
rect 33505 46931 33563 46937
rect 27764 46872 28488 46900
rect 27764 46860 27770 46872
rect 28534 46860 28540 46912
rect 28592 46900 28598 46912
rect 29825 46903 29883 46909
rect 29825 46900 29837 46903
rect 28592 46872 29837 46900
rect 28592 46860 28598 46872
rect 29825 46869 29837 46872
rect 29871 46869 29883 46903
rect 29825 46863 29883 46869
rect 30282 46860 30288 46912
rect 30340 46860 30346 46912
rect 30374 46860 30380 46912
rect 30432 46900 30438 46912
rect 31665 46903 31723 46909
rect 31665 46900 31677 46903
rect 30432 46872 31677 46900
rect 30432 46860 30438 46872
rect 31665 46869 31677 46872
rect 31711 46869 31723 46903
rect 32582 46900 32588 46912
rect 32543 46872 32588 46900
rect 31665 46863 31723 46869
rect 32582 46860 32588 46872
rect 32640 46860 32646 46912
rect 32677 46903 32735 46909
rect 32677 46869 32689 46903
rect 32723 46900 32735 46903
rect 32766 46900 32772 46912
rect 32723 46872 32772 46900
rect 32723 46869 32735 46872
rect 32677 46863 32735 46869
rect 32766 46860 32772 46872
rect 32824 46860 32830 46912
rect 33318 46860 33324 46912
rect 33376 46900 33382 46912
rect 33413 46903 33471 46909
rect 33413 46900 33425 46903
rect 33376 46872 33425 46900
rect 33376 46860 33382 46872
rect 33413 46869 33425 46872
rect 33459 46869 33471 46903
rect 33594 46900 33600 46912
rect 33555 46872 33600 46900
rect 33413 46863 33471 46869
rect 33594 46860 33600 46872
rect 33652 46860 33658 46912
rect 33689 46903 33747 46909
rect 33689 46869 33701 46903
rect 33735 46900 33747 46903
rect 33870 46900 33876 46912
rect 33735 46872 33876 46900
rect 33735 46869 33747 46872
rect 33689 46863 33747 46869
rect 33870 46860 33876 46872
rect 33928 46860 33934 46912
rect 33980 46900 34008 46940
rect 34054 46928 34060 46980
rect 34112 46968 34118 46980
rect 34977 46971 35035 46977
rect 34977 46968 34989 46971
rect 34112 46940 34989 46968
rect 34112 46928 34118 46940
rect 34977 46937 34989 46940
rect 35023 46937 35035 46971
rect 35434 46968 35440 46980
rect 35395 46940 35440 46968
rect 34977 46931 35035 46937
rect 35434 46928 35440 46940
rect 35492 46928 35498 46980
rect 36078 46928 36084 46980
rect 36136 46968 36142 46980
rect 37553 46971 37611 46977
rect 37553 46968 37565 46971
rect 36136 46940 37565 46968
rect 36136 46928 36142 46940
rect 37553 46937 37565 46940
rect 37599 46937 37611 46971
rect 37553 46931 37611 46937
rect 37642 46928 37648 46980
rect 37700 46968 37706 46980
rect 38028 46968 38056 46999
rect 38562 46996 38568 47008
rect 38620 46996 38626 47048
rect 37700 46940 38056 46968
rect 37700 46928 37706 46940
rect 34422 46900 34428 46912
rect 33980 46872 34428 46900
rect 34422 46860 34428 46872
rect 34480 46900 34486 46912
rect 34698 46900 34704 46912
rect 34480 46872 34704 46900
rect 34480 46860 34486 46872
rect 34698 46860 34704 46872
rect 34756 46860 34762 46912
rect 35345 46903 35403 46909
rect 35345 46869 35357 46903
rect 35391 46900 35403 46903
rect 35526 46900 35532 46912
rect 35391 46872 35532 46900
rect 35391 46869 35403 46872
rect 35345 46863 35403 46869
rect 35526 46860 35532 46872
rect 35584 46900 35590 46912
rect 36538 46900 36544 46912
rect 35584 46872 36544 46900
rect 35584 46860 35590 46872
rect 36538 46860 36544 46872
rect 36596 46860 36602 46912
rect 36630 46860 36636 46912
rect 36688 46900 36694 46912
rect 38562 46900 38568 46912
rect 36688 46872 38568 46900
rect 36688 46860 36694 46872
rect 38562 46860 38568 46872
rect 38620 46860 38626 46912
rect 38672 46900 38700 47076
rect 40218 47064 40224 47116
rect 40276 47104 40282 47116
rect 41969 47107 42027 47113
rect 41969 47104 41981 47107
rect 40276 47076 41981 47104
rect 40276 47064 40282 47076
rect 41969 47073 41981 47076
rect 42015 47073 42027 47107
rect 41969 47067 42027 47073
rect 39114 47036 39120 47048
rect 39075 47008 39120 47036
rect 39114 46996 39120 47008
rect 39172 46996 39178 47048
rect 40037 47039 40095 47045
rect 40037 47005 40049 47039
rect 40083 47036 40095 47039
rect 40126 47036 40132 47048
rect 40083 47008 40132 47036
rect 40083 47005 40095 47008
rect 40037 46999 40095 47005
rect 40126 46996 40132 47008
rect 40184 46996 40190 47048
rect 40678 47036 40684 47048
rect 40639 47008 40684 47036
rect 40678 46996 40684 47008
rect 40736 46996 40742 47048
rect 38746 46928 38752 46980
rect 38804 46968 38810 46980
rect 44545 46971 44603 46977
rect 44545 46968 44557 46971
rect 38804 46940 44557 46968
rect 38804 46928 38810 46940
rect 44545 46937 44557 46940
rect 44591 46937 44603 46971
rect 44545 46931 44603 46937
rect 38930 46900 38936 46912
rect 38672 46872 38936 46900
rect 38930 46860 38936 46872
rect 38988 46860 38994 46912
rect 1104 46810 48852 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 48852 46810
rect 1104 46736 48852 46758
rect 16114 46656 16120 46708
rect 16172 46696 16178 46708
rect 17862 46696 17868 46708
rect 16172 46668 17868 46696
rect 16172 46656 16178 46668
rect 17862 46656 17868 46668
rect 17920 46656 17926 46708
rect 20346 46696 20352 46708
rect 20088 46668 20352 46696
rect 12802 46588 12808 46640
rect 12860 46628 12866 46640
rect 19334 46628 19340 46640
rect 12860 46600 19340 46628
rect 12860 46588 12866 46600
rect 19334 46588 19340 46600
rect 19392 46588 19398 46640
rect 6914 46520 6920 46572
rect 6972 46560 6978 46572
rect 17405 46563 17463 46569
rect 6972 46532 7017 46560
rect 6972 46520 6978 46532
rect 17405 46529 17417 46563
rect 17451 46560 17463 46563
rect 17954 46560 17960 46572
rect 17451 46532 17960 46560
rect 17451 46529 17463 46532
rect 17405 46523 17463 46529
rect 17954 46520 17960 46532
rect 18012 46520 18018 46572
rect 18046 46520 18052 46572
rect 18104 46560 18110 46572
rect 18509 46563 18567 46569
rect 18104 46532 18149 46560
rect 18104 46520 18110 46532
rect 18509 46529 18521 46563
rect 18555 46560 18567 46563
rect 19886 46560 19892 46572
rect 18555 46532 19892 46560
rect 18555 46529 18567 46532
rect 18509 46523 18567 46529
rect 19886 46520 19892 46532
rect 19944 46520 19950 46572
rect 20088 46569 20116 46668
rect 20346 46656 20352 46668
rect 20404 46656 20410 46708
rect 21177 46699 21235 46705
rect 21177 46665 21189 46699
rect 21223 46696 21235 46699
rect 22186 46696 22192 46708
rect 21223 46668 22192 46696
rect 21223 46665 21235 46668
rect 21177 46659 21235 46665
rect 22186 46656 22192 46668
rect 22244 46656 22250 46708
rect 22388 46668 23980 46696
rect 20254 46588 20260 46640
rect 20312 46628 20318 46640
rect 22278 46628 22284 46640
rect 20312 46600 22284 46628
rect 20312 46588 20318 46600
rect 22278 46588 22284 46600
rect 22336 46588 22342 46640
rect 20073 46563 20131 46569
rect 20073 46529 20085 46563
rect 20119 46529 20131 46563
rect 21239 46563 21297 46569
rect 20073 46523 20131 46529
rect 20180 46532 20852 46560
rect 19337 46495 19395 46501
rect 19337 46461 19349 46495
rect 19383 46492 19395 46495
rect 20180 46492 20208 46532
rect 19383 46464 20208 46492
rect 19383 46461 19395 46464
rect 19337 46455 19395 46461
rect 20254 46452 20260 46504
rect 20312 46492 20318 46504
rect 20714 46492 20720 46504
rect 20312 46464 20357 46492
rect 20675 46464 20720 46492
rect 20312 46452 20318 46464
rect 20714 46452 20720 46464
rect 20772 46452 20778 46504
rect 20824 46492 20852 46532
rect 21239 46529 21251 46563
rect 21285 46560 21297 46563
rect 21450 46560 21456 46572
rect 21285 46532 21456 46560
rect 21285 46529 21297 46532
rect 21239 46523 21297 46529
rect 21450 46520 21456 46532
rect 21508 46560 21514 46572
rect 22388 46560 22416 46668
rect 22646 46628 22652 46640
rect 22480 46600 22652 46628
rect 22480 46569 22508 46600
rect 22646 46588 22652 46600
rect 22704 46588 22710 46640
rect 23842 46628 23848 46640
rect 23803 46600 23848 46628
rect 23842 46588 23848 46600
rect 23900 46588 23906 46640
rect 23952 46628 23980 46668
rect 25866 46656 25872 46708
rect 25924 46696 25930 46708
rect 25961 46699 26019 46705
rect 25961 46696 25973 46699
rect 25924 46668 25973 46696
rect 25924 46656 25930 46668
rect 25961 46665 25973 46668
rect 26007 46665 26019 46699
rect 25961 46659 26019 46665
rect 26050 46656 26056 46708
rect 26108 46696 26114 46708
rect 26145 46699 26203 46705
rect 26145 46696 26157 46699
rect 26108 46668 26157 46696
rect 26108 46656 26114 46668
rect 26145 46665 26157 46668
rect 26191 46665 26203 46699
rect 26145 46659 26203 46665
rect 26694 46656 26700 46708
rect 26752 46696 26758 46708
rect 26752 46668 28212 46696
rect 26752 46656 26758 46668
rect 28184 46637 28212 46668
rect 28350 46656 28356 46708
rect 28408 46696 28414 46708
rect 28534 46696 28540 46708
rect 28408 46668 28540 46696
rect 28408 46656 28414 46668
rect 28534 46656 28540 46668
rect 28592 46656 28598 46708
rect 29270 46696 29276 46708
rect 29231 46668 29276 46696
rect 29270 46656 29276 46668
rect 29328 46656 29334 46708
rect 30190 46696 30196 46708
rect 30151 46668 30196 46696
rect 30190 46656 30196 46668
rect 30248 46656 30254 46708
rect 31018 46656 31024 46708
rect 31076 46696 31082 46708
rect 32493 46699 32551 46705
rect 32493 46696 32505 46699
rect 31076 46668 32505 46696
rect 31076 46656 31082 46668
rect 32493 46665 32505 46668
rect 32539 46665 32551 46699
rect 32493 46659 32551 46665
rect 33962 46656 33968 46708
rect 34020 46696 34026 46708
rect 34020 46668 34376 46696
rect 34020 46656 34026 46668
rect 27249 46631 27307 46637
rect 27249 46628 27261 46631
rect 23952 46600 27261 46628
rect 27249 46597 27261 46600
rect 27295 46597 27307 46631
rect 27249 46591 27307 46597
rect 28169 46631 28227 46637
rect 28169 46597 28181 46631
rect 28215 46597 28227 46631
rect 28169 46591 28227 46597
rect 31573 46631 31631 46637
rect 31573 46597 31585 46631
rect 31619 46628 31631 46631
rect 32214 46628 32220 46640
rect 31619 46600 32220 46628
rect 31619 46597 31631 46600
rect 31573 46591 31631 46597
rect 32214 46588 32220 46600
rect 32272 46588 32278 46640
rect 32306 46588 32312 46640
rect 32364 46628 32370 46640
rect 34146 46628 34152 46640
rect 32364 46600 34152 46628
rect 32364 46588 32370 46600
rect 34146 46588 34152 46600
rect 34204 46588 34210 46640
rect 34348 46628 34376 46668
rect 34422 46656 34428 46708
rect 34480 46696 34486 46708
rect 34609 46699 34667 46705
rect 34480 46668 34525 46696
rect 34480 46656 34486 46668
rect 34609 46665 34621 46699
rect 34655 46696 34667 46699
rect 35250 46696 35256 46708
rect 34655 46668 35256 46696
rect 34655 46665 34667 46668
rect 34609 46659 34667 46665
rect 35250 46656 35256 46668
rect 35308 46656 35314 46708
rect 35986 46656 35992 46708
rect 36044 46696 36050 46708
rect 36044 46668 39160 46696
rect 36044 46656 36050 46668
rect 38565 46631 38623 46637
rect 38565 46628 38577 46631
rect 34348 46600 34652 46628
rect 21508 46532 22416 46560
rect 22465 46563 22523 46569
rect 21508 46520 21514 46532
rect 22465 46529 22477 46563
rect 22511 46529 22523 46563
rect 22465 46523 22523 46529
rect 22557 46563 22615 46569
rect 22557 46529 22569 46563
rect 22603 46529 22615 46563
rect 22557 46523 22615 46529
rect 21910 46492 21916 46504
rect 20824 46464 21916 46492
rect 21910 46452 21916 46464
rect 21968 46452 21974 46504
rect 22370 46452 22376 46504
rect 22428 46492 22434 46504
rect 22572 46492 22600 46523
rect 23106 46520 23112 46572
rect 23164 46560 23170 46572
rect 24029 46563 24087 46569
rect 24029 46560 24041 46563
rect 23164 46532 24041 46560
rect 23164 46520 23170 46532
rect 24029 46529 24041 46532
rect 24075 46560 24087 46563
rect 24118 46560 24124 46572
rect 24075 46532 24124 46560
rect 24075 46529 24087 46532
rect 24029 46523 24087 46529
rect 24118 46520 24124 46532
rect 24176 46520 24182 46572
rect 24394 46520 24400 46572
rect 24452 46560 24458 46572
rect 24581 46563 24639 46569
rect 24452 46532 24497 46560
rect 24452 46520 24458 46532
rect 24581 46529 24593 46563
rect 24627 46560 24639 46563
rect 24762 46560 24768 46572
rect 24627 46532 24768 46560
rect 24627 46529 24639 46532
rect 24581 46523 24639 46529
rect 24762 46520 24768 46532
rect 24820 46520 24826 46572
rect 25222 46560 25228 46572
rect 25183 46532 25228 46560
rect 25222 46520 25228 46532
rect 25280 46520 25286 46572
rect 25409 46563 25467 46569
rect 25409 46529 25421 46563
rect 25455 46560 25467 46563
rect 25498 46560 25504 46572
rect 25455 46532 25504 46560
rect 25455 46529 25467 46532
rect 25409 46523 25467 46529
rect 25498 46520 25504 46532
rect 25556 46520 25562 46572
rect 25958 46520 25964 46572
rect 26016 46560 26022 46572
rect 26142 46560 26148 46572
rect 26016 46532 26148 46560
rect 26016 46520 26022 46532
rect 26142 46520 26148 46532
rect 26200 46520 26206 46572
rect 27706 46560 27712 46572
rect 27667 46532 27712 46560
rect 27706 46520 27712 46532
rect 27764 46520 27770 46572
rect 27798 46520 27804 46572
rect 27856 46560 27862 46572
rect 28353 46563 28411 46569
rect 28353 46560 28365 46563
rect 27856 46532 28365 46560
rect 27856 46520 27862 46532
rect 28353 46529 28365 46532
rect 28399 46560 28411 46563
rect 28994 46560 29000 46572
rect 28399 46532 28856 46560
rect 28955 46532 29000 46560
rect 28399 46529 28411 46532
rect 28353 46523 28411 46529
rect 22830 46492 22836 46504
rect 22428 46464 22600 46492
rect 22791 46464 22836 46492
rect 22428 46452 22434 46464
rect 22830 46452 22836 46464
rect 22888 46452 22894 46504
rect 23198 46452 23204 46504
rect 23256 46492 23262 46504
rect 24213 46495 24271 46501
rect 24213 46492 24225 46495
rect 23256 46464 24225 46492
rect 23256 46452 23262 46464
rect 24213 46461 24225 46464
rect 24259 46461 24271 46495
rect 24213 46455 24271 46461
rect 24302 46452 24308 46504
rect 24360 46492 24366 46504
rect 26602 46492 26608 46504
rect 24360 46464 24405 46492
rect 26563 46464 26608 46492
rect 24360 46452 24366 46464
rect 26602 46452 26608 46464
rect 26660 46452 26666 46504
rect 27338 46452 27344 46504
rect 27396 46492 27402 46504
rect 27433 46495 27491 46501
rect 27433 46492 27445 46495
rect 27396 46464 27445 46492
rect 27396 46452 27402 46464
rect 27433 46461 27445 46464
rect 27479 46461 27491 46495
rect 28828 46492 28856 46532
rect 28994 46520 29000 46532
rect 29052 46520 29058 46572
rect 29270 46560 29276 46572
rect 29231 46532 29276 46560
rect 29270 46520 29276 46532
rect 29328 46520 29334 46572
rect 29503 46563 29561 46569
rect 29503 46529 29515 46563
rect 29549 46560 29561 46563
rect 30558 46560 30564 46572
rect 29549 46532 30564 46560
rect 29549 46529 29561 46532
rect 29503 46523 29561 46529
rect 30558 46520 30564 46532
rect 30616 46520 30622 46572
rect 30653 46563 30711 46569
rect 30653 46529 30665 46563
rect 30699 46560 30711 46563
rect 31662 46560 31668 46572
rect 30699 46532 31668 46560
rect 30699 46529 30711 46532
rect 30653 46523 30711 46529
rect 31662 46520 31668 46532
rect 31720 46520 31726 46572
rect 31754 46520 31760 46572
rect 31812 46560 31818 46572
rect 32490 46560 32496 46572
rect 31812 46532 31857 46560
rect 32140 46532 32496 46560
rect 31812 46520 31818 46532
rect 29914 46492 29920 46504
rect 28828 46464 29920 46492
rect 27433 46455 27491 46461
rect 29914 46452 29920 46464
rect 29972 46452 29978 46504
rect 30006 46452 30012 46504
rect 30064 46492 30070 46504
rect 30101 46495 30159 46501
rect 30101 46492 30113 46495
rect 30064 46464 30113 46492
rect 30064 46452 30070 46464
rect 30101 46461 30113 46464
rect 30147 46461 30159 46495
rect 30101 46455 30159 46461
rect 30285 46495 30343 46501
rect 30285 46461 30297 46495
rect 30331 46492 30343 46495
rect 30742 46492 30748 46504
rect 30331 46464 30748 46492
rect 30331 46461 30343 46464
rect 30285 46455 30343 46461
rect 30742 46452 30748 46464
rect 30800 46452 30806 46504
rect 30929 46495 30987 46501
rect 30929 46461 30941 46495
rect 30975 46492 30987 46495
rect 31294 46492 31300 46504
rect 30975 46464 31300 46492
rect 30975 46461 30987 46464
rect 30929 46455 30987 46461
rect 31294 46452 31300 46464
rect 31352 46452 31358 46504
rect 31389 46495 31447 46501
rect 31389 46461 31401 46495
rect 31435 46492 31447 46495
rect 32140 46492 32168 46532
rect 32490 46520 32496 46532
rect 32548 46520 32554 46572
rect 32692 46532 34100 46560
rect 32306 46492 32312 46504
rect 31435 46464 32168 46492
rect 32267 46464 32312 46492
rect 31435 46461 31447 46464
rect 31389 46455 31447 46461
rect 32306 46452 32312 46464
rect 32364 46452 32370 46504
rect 18693 46427 18751 46433
rect 18693 46393 18705 46427
rect 18739 46424 18751 46427
rect 20809 46427 20867 46433
rect 20809 46424 20821 46427
rect 18739 46396 20821 46424
rect 18739 46393 18751 46396
rect 18693 46387 18751 46393
rect 20809 46393 20821 46396
rect 20855 46424 20867 46427
rect 21542 46424 21548 46436
rect 20855 46396 21548 46424
rect 20855 46393 20867 46396
rect 20809 46387 20867 46393
rect 21542 46384 21548 46396
rect 21600 46384 21606 46436
rect 22278 46424 22284 46436
rect 22239 46396 22284 46424
rect 22278 46384 22284 46396
rect 22336 46384 22342 46436
rect 22741 46427 22799 46433
rect 22741 46393 22753 46427
rect 22787 46424 22799 46427
rect 22922 46424 22928 46436
rect 22787 46396 22928 46424
rect 22787 46393 22799 46396
rect 22741 46387 22799 46393
rect 22922 46384 22928 46396
rect 22980 46384 22986 46436
rect 23658 46384 23664 46436
rect 23716 46424 23722 46436
rect 25041 46427 25099 46433
rect 25041 46424 25053 46427
rect 23716 46396 25053 46424
rect 23716 46384 23722 46396
rect 25041 46393 25053 46396
rect 25087 46393 25099 46427
rect 25041 46387 25099 46393
rect 25314 46384 25320 46436
rect 25372 46424 25378 46436
rect 25372 46396 27476 46424
rect 25372 46384 25378 46396
rect 18322 46316 18328 46368
rect 18380 46356 18386 46368
rect 19242 46356 19248 46368
rect 18380 46328 19248 46356
rect 18380 46316 18386 46328
rect 19242 46316 19248 46328
rect 19300 46316 19306 46368
rect 19426 46316 19432 46368
rect 19484 46356 19490 46368
rect 19889 46359 19947 46365
rect 19889 46356 19901 46359
rect 19484 46328 19901 46356
rect 19484 46316 19490 46328
rect 19889 46325 19901 46328
rect 19935 46325 19947 46359
rect 19889 46319 19947 46325
rect 20162 46316 20168 46368
rect 20220 46356 20226 46368
rect 21361 46359 21419 46365
rect 21361 46356 21373 46359
rect 20220 46328 21373 46356
rect 20220 46316 20226 46328
rect 21361 46325 21373 46328
rect 21407 46325 21419 46359
rect 21361 46319 21419 46325
rect 23385 46359 23443 46365
rect 23385 46325 23397 46359
rect 23431 46356 23443 46359
rect 25774 46356 25780 46368
rect 23431 46328 25780 46356
rect 23431 46325 23443 46328
rect 23385 46319 23443 46325
rect 25774 46316 25780 46328
rect 25832 46356 25838 46368
rect 26418 46356 26424 46368
rect 25832 46328 26424 46356
rect 25832 46316 25838 46328
rect 26418 46316 26424 46328
rect 26476 46316 26482 46368
rect 26513 46359 26571 46365
rect 26513 46325 26525 46359
rect 26559 46356 26571 46359
rect 26786 46356 26792 46368
rect 26559 46328 26792 46356
rect 26559 46325 26571 46328
rect 26513 46319 26571 46325
rect 26786 46316 26792 46328
rect 26844 46316 26850 46368
rect 27448 46356 27476 46396
rect 27522 46384 27528 46436
rect 27580 46424 27586 46436
rect 27617 46427 27675 46433
rect 27617 46424 27629 46427
rect 27580 46396 27629 46424
rect 27580 46384 27586 46396
rect 27617 46393 27629 46396
rect 27663 46393 27675 46427
rect 29362 46424 29368 46436
rect 27617 46387 27675 46393
rect 27724 46396 29368 46424
rect 27724 46356 27752 46396
rect 29362 46384 29368 46396
rect 29420 46384 29426 46436
rect 30650 46384 30656 46436
rect 30708 46424 30714 46436
rect 32692 46424 32720 46532
rect 32858 46492 32864 46504
rect 32819 46464 32864 46492
rect 32858 46452 32864 46464
rect 32916 46452 32922 46504
rect 33134 46452 33140 46504
rect 33192 46492 33198 46504
rect 33962 46492 33968 46504
rect 33192 46464 33968 46492
rect 33192 46452 33198 46464
rect 33962 46452 33968 46464
rect 34020 46452 34026 46504
rect 34072 46492 34100 46532
rect 34238 46520 34244 46572
rect 34296 46560 34302 46572
rect 34427 46563 34485 46569
rect 34427 46560 34439 46563
rect 34296 46532 34439 46560
rect 34296 46520 34302 46532
rect 34427 46529 34439 46532
rect 34473 46529 34485 46563
rect 34624 46560 34652 46600
rect 35820 46600 38577 46628
rect 35820 46569 35848 46600
rect 38565 46597 38577 46600
rect 38611 46597 38623 46631
rect 38565 46591 38623 46597
rect 35805 46563 35863 46569
rect 34624 46532 35296 46560
rect 34427 46523 34485 46529
rect 35161 46495 35219 46501
rect 35161 46492 35173 46495
rect 34072 46464 35173 46492
rect 35161 46461 35173 46464
rect 35207 46461 35219 46495
rect 35268 46492 35296 46532
rect 35805 46529 35817 46563
rect 35851 46529 35863 46563
rect 36354 46560 36360 46572
rect 36315 46532 36360 46560
rect 35805 46523 35863 46529
rect 36354 46520 36360 46532
rect 36412 46520 36418 46572
rect 36538 46560 36544 46572
rect 36499 46532 36544 46560
rect 36538 46520 36544 46532
rect 36596 46520 36602 46572
rect 38013 46563 38071 46569
rect 36648 46532 37872 46560
rect 35710 46492 35716 46504
rect 35268 46464 35716 46492
rect 35161 46455 35219 46461
rect 35710 46452 35716 46464
rect 35768 46492 35774 46504
rect 35989 46495 36047 46501
rect 35989 46492 36001 46495
rect 35768 46464 36001 46492
rect 35768 46452 35774 46464
rect 35989 46461 36001 46464
rect 36035 46461 36047 46495
rect 36648 46492 36676 46532
rect 35989 46455 36047 46461
rect 36096 46464 36676 46492
rect 30708 46396 32720 46424
rect 30708 46384 30714 46396
rect 32766 46384 32772 46436
rect 32824 46424 32830 46436
rect 35897 46427 35955 46433
rect 35897 46424 35909 46427
rect 32824 46396 35909 46424
rect 32824 46384 32830 46396
rect 35897 46393 35909 46396
rect 35943 46393 35955 46427
rect 35897 46387 35955 46393
rect 27448 46328 27752 46356
rect 27982 46316 27988 46368
rect 28040 46356 28046 46368
rect 28445 46359 28503 46365
rect 28445 46356 28457 46359
rect 28040 46328 28457 46356
rect 28040 46316 28046 46328
rect 28445 46325 28457 46328
rect 28491 46325 28503 46359
rect 28445 46319 28503 46325
rect 29270 46316 29276 46368
rect 29328 46356 29334 46368
rect 31018 46356 31024 46368
rect 29328 46328 31024 46356
rect 29328 46316 29334 46328
rect 31018 46316 31024 46328
rect 31076 46316 31082 46368
rect 32950 46316 32956 46368
rect 33008 46356 33014 46368
rect 33321 46359 33379 46365
rect 33321 46356 33333 46359
rect 33008 46328 33333 46356
rect 33008 46316 33014 46328
rect 33321 46325 33333 46328
rect 33367 46325 33379 46359
rect 33321 46319 33379 46325
rect 34057 46359 34115 46365
rect 34057 46325 34069 46359
rect 34103 46356 34115 46359
rect 34422 46356 34428 46368
rect 34103 46328 34428 46356
rect 34103 46325 34115 46328
rect 34057 46319 34115 46325
rect 34422 46316 34428 46328
rect 34480 46316 34486 46368
rect 34514 46316 34520 46368
rect 34572 46356 34578 46368
rect 36096 46356 36124 46464
rect 36722 46452 36728 46504
rect 36780 46492 36786 46504
rect 37737 46495 37795 46501
rect 37737 46492 37749 46495
rect 36780 46464 37749 46492
rect 36780 46452 36786 46464
rect 37737 46461 37749 46464
rect 37783 46461 37795 46495
rect 37844 46492 37872 46532
rect 38013 46529 38025 46563
rect 38059 46560 38071 46563
rect 38102 46560 38108 46572
rect 38059 46532 38108 46560
rect 38059 46529 38071 46532
rect 38013 46523 38071 46529
rect 38102 46520 38108 46532
rect 38160 46520 38166 46572
rect 38654 46520 38660 46572
rect 38712 46560 38718 46572
rect 38749 46563 38807 46569
rect 38749 46560 38761 46563
rect 38712 46532 38761 46560
rect 38712 46520 38718 46532
rect 38749 46529 38761 46532
rect 38795 46529 38807 46563
rect 38749 46523 38807 46529
rect 38838 46520 38844 46572
rect 38896 46560 38902 46572
rect 39025 46563 39083 46569
rect 39025 46560 39037 46563
rect 38896 46532 39037 46560
rect 38896 46520 38902 46532
rect 39025 46529 39037 46532
rect 39071 46529 39083 46563
rect 39025 46523 39083 46529
rect 38930 46492 38936 46504
rect 37844 46464 38056 46492
rect 38891 46464 38936 46492
rect 37737 46455 37795 46461
rect 36170 46384 36176 46436
rect 36228 46424 36234 46436
rect 37921 46427 37979 46433
rect 37921 46424 37933 46427
rect 36228 46396 37933 46424
rect 36228 46384 36234 46396
rect 37921 46393 37933 46396
rect 37967 46393 37979 46427
rect 37921 46387 37979 46393
rect 37550 46356 37556 46368
rect 34572 46328 36124 46356
rect 37511 46328 37556 46356
rect 34572 46316 34578 46328
rect 37550 46316 37556 46328
rect 37608 46316 37614 46368
rect 38028 46356 38056 46464
rect 38930 46452 38936 46464
rect 38988 46452 38994 46504
rect 39132 46424 39160 46668
rect 39390 46656 39396 46708
rect 39448 46696 39454 46708
rect 41874 46696 41880 46708
rect 39448 46668 41880 46696
rect 39448 46656 39454 46668
rect 41874 46656 41880 46668
rect 41932 46656 41938 46708
rect 40034 46520 40040 46572
rect 40092 46560 40098 46572
rect 41417 46563 41475 46569
rect 41417 46560 41429 46563
rect 40092 46532 41429 46560
rect 40092 46520 40098 46532
rect 41417 46529 41429 46532
rect 41463 46529 41475 46563
rect 41417 46523 41475 46529
rect 42242 46520 42248 46572
rect 42300 46560 42306 46572
rect 42613 46563 42671 46569
rect 42613 46560 42625 46563
rect 42300 46532 42625 46560
rect 42300 46520 42306 46532
rect 42613 46529 42625 46532
rect 42659 46529 42671 46563
rect 43714 46560 43720 46572
rect 43675 46532 43720 46560
rect 42613 46523 42671 46529
rect 43714 46520 43720 46532
rect 43772 46520 43778 46572
rect 44450 46560 44456 46572
rect 44411 46532 44456 46560
rect 44450 46520 44456 46532
rect 44508 46520 44514 46572
rect 39206 46452 39212 46504
rect 39264 46492 39270 46504
rect 40773 46495 40831 46501
rect 40773 46492 40785 46495
rect 39264 46464 40785 46492
rect 39264 46452 39270 46464
rect 40773 46461 40785 46464
rect 40819 46461 40831 46495
rect 40773 46455 40831 46461
rect 40129 46427 40187 46433
rect 40129 46424 40141 46427
rect 39132 46396 40141 46424
rect 40129 46393 40141 46396
rect 40175 46393 40187 46427
rect 40129 46387 40187 46393
rect 39485 46359 39543 46365
rect 39485 46356 39497 46359
rect 38028 46328 39497 46356
rect 39485 46325 39497 46328
rect 39531 46325 39543 46359
rect 39485 46319 39543 46325
rect 1104 46266 48852 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 48852 46266
rect 1104 46192 48852 46214
rect 16942 46112 16948 46164
rect 17000 46152 17006 46164
rect 17497 46155 17555 46161
rect 17497 46152 17509 46155
rect 17000 46124 17509 46152
rect 17000 46112 17006 46124
rect 17497 46121 17509 46124
rect 17543 46152 17555 46155
rect 17862 46152 17868 46164
rect 17543 46124 17868 46152
rect 17543 46121 17555 46124
rect 17497 46115 17555 46121
rect 17862 46112 17868 46124
rect 17920 46112 17926 46164
rect 18046 46112 18052 46164
rect 18104 46152 18110 46164
rect 19705 46155 19763 46161
rect 19705 46152 19717 46155
rect 18104 46124 19717 46152
rect 18104 46112 18110 46124
rect 19705 46121 19717 46124
rect 19751 46121 19763 46155
rect 20530 46152 20536 46164
rect 19705 46115 19763 46121
rect 19812 46124 20536 46152
rect 18233 46087 18291 46093
rect 18233 46053 18245 46087
rect 18279 46084 18291 46087
rect 19058 46084 19064 46096
rect 18279 46056 19064 46084
rect 18279 46053 18291 46056
rect 18233 46047 18291 46053
rect 19058 46044 19064 46056
rect 19116 46044 19122 46096
rect 19242 46044 19248 46096
rect 19300 46084 19306 46096
rect 19812 46084 19840 46124
rect 20530 46112 20536 46124
rect 20588 46112 20594 46164
rect 20625 46155 20683 46161
rect 20625 46121 20637 46155
rect 20671 46152 20683 46155
rect 22830 46152 22836 46164
rect 20671 46124 22836 46152
rect 20671 46121 20683 46124
rect 20625 46115 20683 46121
rect 22830 46112 22836 46124
rect 22888 46112 22894 46164
rect 24765 46155 24823 46161
rect 24765 46121 24777 46155
rect 24811 46152 24823 46155
rect 25682 46152 25688 46164
rect 24811 46124 25688 46152
rect 24811 46121 24823 46124
rect 24765 46115 24823 46121
rect 25682 46112 25688 46124
rect 25740 46112 25746 46164
rect 27338 46152 27344 46164
rect 27299 46124 27344 46152
rect 27338 46112 27344 46124
rect 27396 46112 27402 46164
rect 28810 46112 28816 46164
rect 28868 46152 28874 46164
rect 29825 46155 29883 46161
rect 29825 46152 29837 46155
rect 28868 46124 29837 46152
rect 28868 46112 28874 46124
rect 29825 46121 29837 46124
rect 29871 46121 29883 46155
rect 30834 46152 30840 46164
rect 30795 46124 30840 46152
rect 29825 46115 29883 46121
rect 30834 46112 30840 46124
rect 30892 46112 30898 46164
rect 32490 46112 32496 46164
rect 32548 46152 32554 46164
rect 32548 46124 32996 46152
rect 32548 46112 32554 46124
rect 19300 46056 19840 46084
rect 19300 46044 19306 46056
rect 19886 46044 19892 46096
rect 19944 46084 19950 46096
rect 21453 46087 21511 46093
rect 21453 46084 21465 46087
rect 19944 46056 21465 46084
rect 19944 46044 19950 46056
rect 21453 46053 21465 46056
rect 21499 46053 21511 46087
rect 22646 46084 22652 46096
rect 21453 46047 21511 46053
rect 22066 46056 22652 46084
rect 19978 46016 19984 46028
rect 12406 45988 19984 46016
rect 11698 45908 11704 45960
rect 11756 45948 11762 45960
rect 12406 45948 12434 45988
rect 19978 45976 19984 45988
rect 20036 45976 20042 46028
rect 22066 46016 22094 46056
rect 22646 46044 22652 46056
rect 22704 46044 22710 46096
rect 25222 46044 25228 46096
rect 25280 46084 25286 46096
rect 26142 46084 26148 46096
rect 25280 46056 26148 46084
rect 25280 46044 25286 46056
rect 25516 46025 25544 46056
rect 26142 46044 26148 46056
rect 26200 46084 26206 46096
rect 27430 46084 27436 46096
rect 26200 46056 27436 46084
rect 26200 46044 26206 46056
rect 27430 46044 27436 46056
rect 27488 46044 27494 46096
rect 27614 46044 27620 46096
rect 27672 46084 27678 46096
rect 27672 46056 27936 46084
rect 27672 46044 27678 46056
rect 23385 46019 23443 46025
rect 23385 46016 23397 46019
rect 20732 45988 22094 46016
rect 22480 45988 23397 46016
rect 11756 45920 12434 45948
rect 18877 45951 18935 45957
rect 11756 45908 11762 45920
rect 18877 45917 18889 45951
rect 18923 45917 18935 45951
rect 19886 45948 19892 45960
rect 19847 45920 19892 45948
rect 18877 45911 18935 45917
rect 17218 45840 17224 45892
rect 17276 45880 17282 45892
rect 18892 45880 18920 45911
rect 19886 45908 19892 45920
rect 19944 45908 19950 45960
rect 20073 45951 20131 45957
rect 20073 45917 20085 45951
rect 20119 45948 20131 45951
rect 20162 45948 20168 45960
rect 20119 45920 20168 45948
rect 20119 45917 20131 45920
rect 20073 45911 20131 45917
rect 20162 45908 20168 45920
rect 20220 45908 20226 45960
rect 20732 45957 20760 45988
rect 20717 45951 20775 45957
rect 20717 45917 20729 45951
rect 20763 45917 20775 45951
rect 20717 45911 20775 45917
rect 21450 45908 21456 45960
rect 21508 45948 21514 45960
rect 21633 45951 21691 45957
rect 21633 45948 21645 45951
rect 21508 45920 21645 45948
rect 21508 45908 21514 45920
rect 21633 45917 21645 45920
rect 21679 45917 21691 45951
rect 21633 45911 21691 45917
rect 21821 45951 21879 45957
rect 21821 45917 21833 45951
rect 21867 45948 21879 45951
rect 22002 45948 22008 45960
rect 21867 45920 22008 45948
rect 21867 45917 21879 45920
rect 21821 45911 21879 45917
rect 22002 45908 22008 45920
rect 22060 45908 22066 45960
rect 22278 45948 22284 45960
rect 22239 45920 22284 45948
rect 22278 45908 22284 45920
rect 22336 45908 22342 45960
rect 22480 45957 22508 45988
rect 23385 45985 23397 45988
rect 23431 45985 23443 46019
rect 23385 45979 23443 45985
rect 25501 46019 25559 46025
rect 25501 45985 25513 46019
rect 25547 45985 25559 46019
rect 25501 45979 25559 45985
rect 26602 45976 26608 46028
rect 26660 46016 26666 46028
rect 27706 46016 27712 46028
rect 26660 45988 27712 46016
rect 26660 45976 26666 45988
rect 27706 45976 27712 45988
rect 27764 46016 27770 46028
rect 27908 46016 27936 46056
rect 28718 46044 28724 46096
rect 28776 46084 28782 46096
rect 28909 46087 28967 46093
rect 28909 46084 28921 46087
rect 28776 46056 28921 46084
rect 28776 46044 28782 46056
rect 28909 46053 28921 46056
rect 28955 46053 28967 46087
rect 28909 46047 28967 46053
rect 28997 46087 29055 46093
rect 28997 46053 29009 46087
rect 29043 46084 29055 46087
rect 29043 46056 29224 46084
rect 29043 46053 29055 46056
rect 28997 46047 29055 46053
rect 28074 46016 28080 46028
rect 27764 45988 27844 46016
rect 27908 45988 28080 46016
rect 27764 45976 27770 45988
rect 22465 45951 22523 45957
rect 22465 45917 22477 45951
rect 22511 45917 22523 45951
rect 22646 45948 22652 45960
rect 22607 45920 22652 45948
rect 22465 45911 22523 45917
rect 20438 45880 20444 45892
rect 17276 45852 18736 45880
rect 18892 45852 20444 45880
rect 17276 45840 17282 45852
rect 18708 45821 18736 45852
rect 20438 45840 20444 45852
rect 20496 45840 20502 45892
rect 20901 45883 20959 45889
rect 20901 45849 20913 45883
rect 20947 45880 20959 45883
rect 21726 45880 21732 45892
rect 20947 45852 21732 45880
rect 20947 45849 20959 45852
rect 20901 45843 20959 45849
rect 21726 45840 21732 45852
rect 21784 45840 21790 45892
rect 21910 45840 21916 45892
rect 21968 45880 21974 45892
rect 22480 45880 22508 45911
rect 22646 45908 22652 45920
rect 22704 45908 22710 45960
rect 22922 45948 22928 45960
rect 22883 45920 22928 45948
rect 22922 45908 22928 45920
rect 22980 45908 22986 45960
rect 23569 45951 23627 45957
rect 23569 45917 23581 45951
rect 23615 45948 23627 45951
rect 23750 45948 23756 45960
rect 23615 45920 23756 45948
rect 23615 45917 23627 45920
rect 23569 45911 23627 45917
rect 23750 45908 23756 45920
rect 23808 45908 23814 45960
rect 25685 45951 25743 45957
rect 25685 45917 25697 45951
rect 25731 45917 25743 45951
rect 25685 45911 25743 45917
rect 21968 45852 22508 45880
rect 21968 45840 21974 45852
rect 18693 45815 18751 45821
rect 18693 45781 18705 45815
rect 18739 45812 18751 45815
rect 20714 45812 20720 45824
rect 18739 45784 20720 45812
rect 18739 45781 18751 45784
rect 18693 45775 18751 45781
rect 20714 45772 20720 45784
rect 20772 45772 20778 45824
rect 20990 45772 20996 45824
rect 21048 45812 21054 45824
rect 22940 45812 22968 45908
rect 23937 45883 23995 45889
rect 23937 45849 23949 45883
rect 23983 45880 23995 45883
rect 24118 45880 24124 45892
rect 23983 45852 24124 45880
rect 23983 45849 23995 45852
rect 23937 45843 23995 45849
rect 24118 45840 24124 45852
rect 24176 45880 24182 45892
rect 24854 45880 24860 45892
rect 24176 45852 24860 45880
rect 24176 45840 24182 45852
rect 24854 45840 24860 45852
rect 24912 45840 24918 45892
rect 23658 45812 23664 45824
rect 21048 45784 22968 45812
rect 23619 45784 23664 45812
rect 21048 45772 21054 45784
rect 23658 45772 23664 45784
rect 23716 45772 23722 45824
rect 23753 45815 23811 45821
rect 23753 45781 23765 45815
rect 23799 45812 23811 45815
rect 24026 45812 24032 45824
rect 23799 45784 24032 45812
rect 23799 45781 23811 45784
rect 23753 45775 23811 45781
rect 24026 45772 24032 45784
rect 24084 45772 24090 45824
rect 24394 45772 24400 45824
rect 24452 45812 24458 45824
rect 25317 45815 25375 45821
rect 25317 45812 25329 45815
rect 24452 45784 25329 45812
rect 24452 45772 24458 45784
rect 25317 45781 25329 45784
rect 25363 45781 25375 45815
rect 25700 45812 25728 45911
rect 25774 45908 25780 45960
rect 25832 45948 25838 45960
rect 26510 45948 26516 45960
rect 25832 45920 25877 45948
rect 26471 45920 26516 45948
rect 25832 45908 25838 45920
rect 26510 45908 26516 45920
rect 26568 45908 26574 45960
rect 26694 45908 26700 45960
rect 26752 45948 26758 45960
rect 26789 45951 26847 45957
rect 26789 45948 26801 45951
rect 26752 45920 26801 45948
rect 26752 45908 26758 45920
rect 26789 45917 26801 45920
rect 26835 45917 26847 45951
rect 26789 45911 26847 45917
rect 27525 45951 27583 45957
rect 27525 45917 27537 45951
rect 27571 45917 27583 45951
rect 27525 45911 27583 45917
rect 26326 45880 26332 45892
rect 26287 45852 26332 45880
rect 26326 45840 26332 45852
rect 26384 45840 26390 45892
rect 27540 45880 27568 45911
rect 27614 45908 27620 45960
rect 27672 45948 27678 45960
rect 27816 45957 27844 45988
rect 28074 45976 28080 45988
rect 28132 46016 28138 46028
rect 29012 46016 29040 46047
rect 28132 45988 29040 46016
rect 29196 46016 29224 46056
rect 31018 46044 31024 46096
rect 31076 46084 31082 46096
rect 31938 46084 31944 46096
rect 31076 46056 31944 46084
rect 31076 46044 31082 46056
rect 31938 46044 31944 46056
rect 31996 46044 32002 46096
rect 32766 46084 32772 46096
rect 32048 46056 32772 46084
rect 29730 46016 29736 46028
rect 28132 45976 28138 45988
rect 27801 45951 27859 45957
rect 27672 45920 27717 45948
rect 27672 45908 27678 45920
rect 27801 45917 27813 45951
rect 27847 45917 27859 45951
rect 27801 45911 27859 45917
rect 27893 45951 27951 45957
rect 27893 45917 27905 45951
rect 27939 45948 27951 45951
rect 27939 45920 28212 45948
rect 27939 45917 27951 45920
rect 27893 45911 27951 45917
rect 27706 45880 27712 45892
rect 27540 45852 27712 45880
rect 26697 45815 26755 45821
rect 26697 45812 26709 45815
rect 25700 45784 26709 45812
rect 25317 45775 25375 45781
rect 26697 45781 26709 45784
rect 26743 45812 26755 45815
rect 26786 45812 26792 45824
rect 26743 45784 26792 45812
rect 26743 45781 26755 45784
rect 26697 45775 26755 45781
rect 26786 45772 26792 45784
rect 26844 45812 26850 45824
rect 27540 45812 27568 45852
rect 27706 45840 27712 45852
rect 27764 45840 27770 45892
rect 28184 45880 28212 45920
rect 28442 45908 28448 45960
rect 28500 45948 28506 45960
rect 28537 45951 28595 45957
rect 28537 45948 28549 45951
rect 28500 45920 28549 45948
rect 28500 45908 28506 45920
rect 28537 45917 28549 45920
rect 28583 45917 28595 45951
rect 28537 45911 28595 45917
rect 28718 45908 28724 45960
rect 28776 45950 28782 45960
rect 28813 45951 28871 45957
rect 28813 45950 28825 45951
rect 28776 45922 28825 45950
rect 28776 45908 28782 45922
rect 28813 45917 28825 45922
rect 28859 45917 28871 45951
rect 29086 45942 29092 45994
rect 29144 45942 29150 45994
rect 29196 45988 29736 46016
rect 29730 45976 29736 45988
rect 29788 45976 29794 46028
rect 32048 46016 32076 46056
rect 32766 46044 32772 46056
rect 32824 46044 32830 46096
rect 32968 46093 32996 46124
rect 33594 46112 33600 46164
rect 33652 46152 33658 46164
rect 34330 46152 34336 46164
rect 33652 46124 34336 46152
rect 33652 46112 33658 46124
rect 34330 46112 34336 46124
rect 34388 46112 34394 46164
rect 35529 46155 35587 46161
rect 35529 46121 35541 46155
rect 35575 46152 35587 46155
rect 36722 46152 36728 46164
rect 35575 46124 36728 46152
rect 35575 46121 35587 46124
rect 35529 46115 35587 46121
rect 36722 46112 36728 46124
rect 36780 46112 36786 46164
rect 37918 46112 37924 46164
rect 37976 46152 37982 46164
rect 38286 46152 38292 46164
rect 37976 46124 38292 46152
rect 37976 46112 37982 46124
rect 38286 46112 38292 46124
rect 38344 46112 38350 46164
rect 39298 46112 39304 46164
rect 39356 46152 39362 46164
rect 40681 46155 40739 46161
rect 40681 46152 40693 46155
rect 39356 46124 40693 46152
rect 39356 46112 39362 46124
rect 40681 46121 40693 46124
rect 40727 46121 40739 46155
rect 41322 46152 41328 46164
rect 41283 46124 41328 46152
rect 40681 46115 40739 46121
rect 41322 46112 41328 46124
rect 41380 46112 41386 46164
rect 41506 46112 41512 46164
rect 41564 46152 41570 46164
rect 41969 46155 42027 46161
rect 41969 46152 41981 46155
rect 41564 46124 41981 46152
rect 41564 46112 41570 46124
rect 41969 46121 41981 46124
rect 42015 46121 42027 46155
rect 43806 46152 43812 46164
rect 43767 46124 43812 46152
rect 41969 46115 42027 46121
rect 43806 46112 43812 46124
rect 43864 46112 43870 46164
rect 32953 46087 33011 46093
rect 32953 46053 32965 46087
rect 32999 46053 33011 46087
rect 32953 46047 33011 46053
rect 36998 46044 37004 46096
rect 37056 46084 37062 46096
rect 40037 46087 40095 46093
rect 40037 46084 40049 46087
rect 37056 46056 40049 46084
rect 37056 46044 37062 46056
rect 40037 46053 40049 46056
rect 40083 46053 40095 46087
rect 40037 46047 40095 46053
rect 40770 46044 40776 46096
rect 40828 46084 40834 46096
rect 42613 46087 42671 46093
rect 42613 46084 42625 46087
rect 40828 46056 42625 46084
rect 40828 46044 40834 46056
rect 42613 46053 42625 46056
rect 42659 46084 42671 46087
rect 43165 46087 43223 46093
rect 43165 46084 43177 46087
rect 42659 46056 43177 46084
rect 42659 46053 42671 46056
rect 42613 46047 42671 46053
rect 43165 46053 43177 46056
rect 43211 46053 43223 46087
rect 43165 46047 43223 46053
rect 36541 46019 36599 46025
rect 36541 46016 36553 46019
rect 31726 45988 32076 46016
rect 32140 45988 36553 46016
rect 30009 45951 30067 45957
rect 30009 45948 30021 45951
rect 28813 45911 28871 45917
rect 29089 45917 29101 45942
rect 29135 45917 29147 45942
rect 29089 45911 29147 45917
rect 29196 45920 30021 45948
rect 28350 45880 28356 45892
rect 28184 45852 28356 45880
rect 28350 45840 28356 45852
rect 28408 45840 28414 45892
rect 28994 45840 29000 45892
rect 29052 45880 29058 45892
rect 29196 45880 29224 45920
rect 30009 45917 30021 45920
rect 30055 45948 30067 45951
rect 30374 45948 30380 45960
rect 30055 45920 30380 45948
rect 30055 45917 30067 45920
rect 30009 45911 30067 45917
rect 30374 45908 30380 45920
rect 30432 45908 30438 45960
rect 30742 45908 30748 45960
rect 30800 45948 30806 45960
rect 31021 45951 31079 45957
rect 31021 45948 31033 45951
rect 30800 45920 31033 45948
rect 30800 45908 30806 45920
rect 31021 45917 31033 45920
rect 31067 45948 31079 45951
rect 31726 45948 31754 45988
rect 32030 45948 32036 45960
rect 31067 45920 31754 45948
rect 31991 45920 32036 45948
rect 31067 45917 31079 45920
rect 31021 45911 31079 45917
rect 32030 45908 32036 45920
rect 32088 45908 32094 45960
rect 30282 45880 30288 45892
rect 29052 45852 29224 45880
rect 30195 45852 30288 45880
rect 29052 45840 29058 45852
rect 30282 45840 30288 45852
rect 30340 45880 30346 45892
rect 30834 45880 30840 45892
rect 30340 45852 30840 45880
rect 30340 45840 30346 45852
rect 30834 45840 30840 45852
rect 30892 45840 30898 45892
rect 31294 45880 31300 45892
rect 31255 45852 31300 45880
rect 31294 45840 31300 45852
rect 31352 45840 31358 45892
rect 31662 45880 31668 45892
rect 31404 45852 31668 45880
rect 26844 45784 27568 45812
rect 26844 45772 26850 45784
rect 28902 45772 28908 45824
rect 28960 45812 28966 45824
rect 29546 45812 29552 45824
rect 28960 45784 29552 45812
rect 28960 45772 28966 45784
rect 29546 45772 29552 45784
rect 29604 45772 29610 45824
rect 30006 45772 30012 45824
rect 30064 45812 30070 45824
rect 30193 45815 30251 45821
rect 30193 45812 30205 45815
rect 30064 45784 30205 45812
rect 30064 45772 30070 45784
rect 30193 45781 30205 45784
rect 30239 45812 30251 45815
rect 31018 45812 31024 45824
rect 30239 45784 31024 45812
rect 30239 45781 30251 45784
rect 30193 45775 30251 45781
rect 31018 45772 31024 45784
rect 31076 45772 31082 45824
rect 31205 45815 31263 45821
rect 31205 45781 31217 45815
rect 31251 45812 31263 45815
rect 31404 45812 31432 45852
rect 31662 45840 31668 45852
rect 31720 45840 31726 45892
rect 31846 45880 31852 45892
rect 31807 45852 31852 45880
rect 31846 45840 31852 45852
rect 31904 45840 31910 45892
rect 31251 45784 31432 45812
rect 31251 45781 31263 45784
rect 31205 45775 31263 45781
rect 31478 45772 31484 45824
rect 31536 45812 31542 45824
rect 32140 45812 32168 45988
rect 36541 45985 36553 45988
rect 36587 45985 36599 46019
rect 37918 46016 37924 46028
rect 37879 45988 37924 46016
rect 36541 45979 36599 45985
rect 37918 45976 37924 45988
rect 37976 45976 37982 46028
rect 38286 45976 38292 46028
rect 38344 46016 38350 46028
rect 38657 46019 38715 46025
rect 38657 46016 38669 46019
rect 38344 45988 38669 46016
rect 38344 45976 38350 45988
rect 38657 45985 38669 45988
rect 38703 45985 38715 46019
rect 38657 45979 38715 45985
rect 32309 45951 32367 45957
rect 32309 45917 32321 45951
rect 32355 45948 32367 45951
rect 33134 45948 33140 45960
rect 32355 45920 33140 45948
rect 32355 45917 32367 45920
rect 32309 45911 32367 45917
rect 33134 45908 33140 45920
rect 33192 45948 33198 45960
rect 33781 45951 33839 45957
rect 33781 45948 33793 45951
rect 33192 45920 33793 45948
rect 33192 45908 33198 45920
rect 33781 45917 33793 45920
rect 33827 45917 33839 45951
rect 33962 45948 33968 45960
rect 33923 45920 33968 45948
rect 33781 45911 33839 45917
rect 33962 45908 33968 45920
rect 34020 45908 34026 45960
rect 34330 45948 34336 45960
rect 34291 45920 34336 45948
rect 34330 45908 34336 45920
rect 34388 45908 34394 45960
rect 34606 45908 34612 45960
rect 34664 45948 34670 45960
rect 34974 45948 34980 45960
rect 34664 45920 34980 45948
rect 34664 45908 34670 45920
rect 34974 45908 34980 45920
rect 35032 45908 35038 45960
rect 35526 45908 35532 45960
rect 35584 45948 35590 45960
rect 35805 45951 35863 45957
rect 35584 45936 35664 45948
rect 35704 45939 35762 45945
rect 35704 45936 35716 45939
rect 35584 45920 35716 45936
rect 35584 45908 35590 45920
rect 35636 45908 35716 45920
rect 33318 45880 33324 45892
rect 33279 45852 33324 45880
rect 33318 45840 33324 45852
rect 33376 45840 33382 45892
rect 34422 45840 34428 45892
rect 34480 45880 34486 45892
rect 35544 45880 35572 45908
rect 35704 45905 35716 45908
rect 35750 45905 35762 45939
rect 35805 45917 35817 45951
rect 35851 45917 35863 45951
rect 35805 45911 35863 45917
rect 35704 45899 35762 45905
rect 34480 45852 35572 45880
rect 35820 45880 35848 45911
rect 35894 45908 35900 45960
rect 35952 45948 35958 45960
rect 35989 45951 36047 45957
rect 35989 45948 36001 45951
rect 35952 45920 36001 45948
rect 35952 45908 35958 45920
rect 35989 45917 36001 45920
rect 36035 45917 36047 45951
rect 35989 45911 36047 45917
rect 36078 45908 36084 45960
rect 36136 45948 36142 45960
rect 36136 45920 36181 45948
rect 36136 45908 36142 45920
rect 36354 45908 36360 45960
rect 36412 45948 36418 45960
rect 37737 45951 37795 45957
rect 37737 45948 37749 45951
rect 36412 45920 37749 45948
rect 36412 45908 36418 45920
rect 37737 45917 37749 45920
rect 37783 45948 37795 45951
rect 37783 45920 37964 45948
rect 37783 45917 37795 45920
rect 37737 45911 37795 45917
rect 36262 45880 36268 45892
rect 35820 45852 36268 45880
rect 34480 45840 34486 45852
rect 36262 45840 36268 45852
rect 36320 45840 36326 45892
rect 31536 45784 32168 45812
rect 32217 45815 32275 45821
rect 31536 45772 31542 45784
rect 32217 45781 32229 45815
rect 32263 45812 32275 45815
rect 32582 45812 32588 45824
rect 32263 45784 32588 45812
rect 32263 45781 32275 45784
rect 32217 45775 32275 45781
rect 32582 45772 32588 45784
rect 32640 45772 32646 45824
rect 32858 45812 32864 45824
rect 32819 45784 32864 45812
rect 32858 45772 32864 45784
rect 32916 45772 32922 45824
rect 33594 45772 33600 45824
rect 33652 45812 33658 45824
rect 33965 45815 34023 45821
rect 33965 45812 33977 45815
rect 33652 45784 33977 45812
rect 33652 45772 33658 45784
rect 33965 45781 33977 45784
rect 34011 45781 34023 45815
rect 37090 45812 37096 45824
rect 37051 45784 37096 45812
rect 33965 45775 34023 45781
rect 37090 45772 37096 45784
rect 37148 45772 37154 45824
rect 37936 45812 37964 45920
rect 38378 45908 38384 45960
rect 38436 45948 38442 45960
rect 38749 45951 38807 45957
rect 38749 45948 38761 45951
rect 38436 45920 38761 45948
rect 38436 45908 38442 45920
rect 38749 45917 38761 45920
rect 38795 45917 38807 45951
rect 38749 45911 38807 45917
rect 38838 45908 38844 45960
rect 38896 45948 38902 45960
rect 39025 45951 39083 45957
rect 39025 45948 39037 45951
rect 38896 45920 39037 45948
rect 38896 45908 38902 45920
rect 39025 45917 39037 45920
rect 39071 45917 39083 45951
rect 39206 45948 39212 45960
rect 39167 45920 39212 45948
rect 39025 45911 39083 45917
rect 39206 45908 39212 45920
rect 39264 45908 39270 45960
rect 38010 45840 38016 45892
rect 38068 45880 38074 45892
rect 39390 45880 39396 45892
rect 38068 45852 39396 45880
rect 38068 45840 38074 45852
rect 39390 45840 39396 45852
rect 39448 45840 39454 45892
rect 38746 45812 38752 45824
rect 37936 45784 38752 45812
rect 38746 45772 38752 45784
rect 38804 45772 38810 45824
rect 1104 45722 48852 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 48852 45722
rect 1104 45648 48852 45670
rect 13906 45568 13912 45620
rect 13964 45608 13970 45620
rect 20625 45611 20683 45617
rect 20625 45608 20637 45611
rect 13964 45580 20637 45608
rect 13964 45568 13970 45580
rect 20625 45577 20637 45580
rect 20671 45577 20683 45611
rect 20806 45608 20812 45620
rect 20767 45580 20812 45608
rect 20625 45571 20683 45577
rect 20806 45568 20812 45580
rect 20864 45568 20870 45620
rect 22646 45568 22652 45620
rect 22704 45608 22710 45620
rect 23201 45611 23259 45617
rect 23201 45608 23213 45611
rect 22704 45580 23213 45608
rect 22704 45568 22710 45580
rect 23201 45577 23213 45580
rect 23247 45577 23259 45611
rect 23201 45571 23259 45577
rect 23290 45568 23296 45620
rect 23348 45608 23354 45620
rect 24673 45611 24731 45617
rect 24673 45608 24685 45611
rect 23348 45580 24685 45608
rect 23348 45568 23354 45580
rect 24673 45577 24685 45580
rect 24719 45577 24731 45611
rect 24854 45608 24860 45620
rect 24815 45580 24860 45608
rect 24673 45571 24731 45577
rect 24854 45568 24860 45580
rect 24912 45568 24918 45620
rect 24949 45611 25007 45617
rect 24949 45577 24961 45611
rect 24995 45608 25007 45611
rect 25958 45608 25964 45620
rect 24995 45580 25964 45608
rect 24995 45577 25007 45580
rect 24949 45571 25007 45577
rect 25958 45568 25964 45580
rect 26016 45568 26022 45620
rect 26050 45568 26056 45620
rect 26108 45608 26114 45620
rect 26145 45611 26203 45617
rect 26145 45608 26157 45611
rect 26108 45580 26157 45608
rect 26108 45568 26114 45580
rect 26145 45577 26157 45580
rect 26191 45577 26203 45611
rect 26145 45571 26203 45577
rect 26237 45611 26295 45617
rect 26237 45577 26249 45611
rect 26283 45608 26295 45611
rect 26326 45608 26332 45620
rect 26283 45580 26332 45608
rect 26283 45577 26295 45580
rect 26237 45571 26295 45577
rect 26326 45568 26332 45580
rect 26384 45568 26390 45620
rect 26510 45568 26516 45620
rect 26568 45608 26574 45620
rect 28718 45608 28724 45620
rect 26568 45580 28724 45608
rect 26568 45568 26574 45580
rect 28718 45568 28724 45580
rect 28776 45608 28782 45620
rect 30926 45608 30932 45620
rect 28776 45580 30932 45608
rect 28776 45568 28782 45580
rect 30926 45568 30932 45580
rect 30984 45568 30990 45620
rect 32306 45568 32312 45620
rect 32364 45608 32370 45620
rect 32861 45611 32919 45617
rect 32861 45608 32873 45611
rect 32364 45580 32873 45608
rect 32364 45568 32370 45580
rect 32861 45577 32873 45580
rect 32907 45577 32919 45611
rect 32861 45571 32919 45577
rect 32950 45568 32956 45620
rect 33008 45608 33014 45620
rect 37090 45608 37096 45620
rect 33008 45580 37096 45608
rect 33008 45568 33014 45580
rect 37090 45568 37096 45580
rect 37148 45568 37154 45620
rect 37918 45568 37924 45620
rect 37976 45608 37982 45620
rect 38013 45611 38071 45617
rect 38013 45608 38025 45611
rect 37976 45580 38025 45608
rect 37976 45568 37982 45580
rect 38013 45577 38025 45580
rect 38059 45577 38071 45611
rect 38013 45571 38071 45577
rect 38194 45568 38200 45620
rect 38252 45608 38258 45620
rect 43806 45608 43812 45620
rect 38252 45580 39620 45608
rect 38252 45568 38258 45580
rect 19981 45543 20039 45549
rect 19981 45509 19993 45543
rect 20027 45540 20039 45543
rect 20990 45540 20996 45552
rect 20027 45512 20996 45540
rect 20027 45509 20039 45512
rect 19981 45503 20039 45509
rect 20990 45500 20996 45512
rect 21048 45500 21054 45552
rect 24121 45543 24179 45549
rect 22296 45512 23152 45540
rect 19245 45475 19303 45481
rect 19245 45441 19257 45475
rect 19291 45472 19303 45475
rect 19426 45472 19432 45484
rect 19291 45444 19432 45472
rect 19291 45441 19303 45444
rect 19245 45435 19303 45441
rect 19426 45432 19432 45444
rect 19484 45432 19490 45484
rect 22296 45481 22324 45512
rect 19889 45475 19947 45481
rect 19889 45441 19901 45475
rect 19935 45441 19947 45475
rect 19889 45435 19947 45441
rect 20807 45475 20865 45481
rect 20807 45441 20819 45475
rect 20853 45472 20865 45475
rect 22281 45475 22339 45481
rect 22281 45472 22293 45475
rect 20853 45444 22293 45472
rect 20853 45441 20865 45444
rect 20807 45435 20865 45441
rect 22281 45441 22293 45444
rect 22327 45441 22339 45475
rect 22281 45435 22339 45441
rect 19794 45404 19800 45416
rect 18708 45376 19800 45404
rect 2774 45228 2780 45280
rect 2832 45268 2838 45280
rect 18708 45277 18736 45376
rect 19794 45364 19800 45376
rect 19852 45404 19858 45416
rect 19904 45404 19932 45435
rect 19852 45376 19932 45404
rect 19852 45364 19858 45376
rect 20530 45364 20536 45416
rect 20588 45404 20594 45416
rect 21269 45407 21327 45413
rect 21269 45404 21281 45407
rect 20588 45376 21281 45404
rect 20588 45364 20594 45376
rect 21269 45373 21281 45376
rect 21315 45373 21327 45407
rect 21269 45367 21327 45373
rect 22002 45364 22008 45416
rect 22060 45404 22066 45416
rect 22462 45404 22468 45416
rect 22060 45376 22468 45404
rect 22060 45364 22066 45376
rect 22462 45364 22468 45376
rect 22520 45364 22526 45416
rect 23017 45407 23075 45413
rect 23017 45373 23029 45407
rect 23063 45373 23075 45407
rect 23124 45404 23152 45512
rect 24121 45509 24133 45543
rect 24167 45540 24179 45543
rect 24210 45540 24216 45552
rect 24167 45512 24216 45540
rect 24167 45509 24179 45512
rect 24121 45503 24179 45509
rect 24210 45500 24216 45512
rect 24268 45540 24274 45552
rect 24762 45540 24768 45552
rect 24268 45512 24768 45540
rect 24268 45500 24274 45512
rect 24762 45500 24768 45512
rect 24820 45500 24826 45552
rect 25133 45543 25191 45549
rect 25133 45509 25145 45543
rect 25179 45540 25191 45543
rect 25590 45540 25596 45552
rect 25179 45512 25596 45540
rect 25179 45509 25191 45512
rect 25133 45503 25191 45509
rect 25590 45500 25596 45512
rect 25648 45500 25654 45552
rect 25866 45500 25872 45552
rect 25924 45540 25930 45552
rect 27341 45543 27399 45549
rect 27341 45540 27353 45543
rect 25924 45512 27353 45540
rect 25924 45500 25930 45512
rect 27341 45509 27353 45512
rect 27387 45509 27399 45543
rect 27341 45503 27399 45509
rect 28166 45500 28172 45552
rect 28224 45540 28230 45552
rect 30006 45540 30012 45552
rect 28224 45512 30012 45540
rect 28224 45500 28230 45512
rect 23201 45475 23259 45481
rect 23201 45441 23213 45475
rect 23247 45472 23259 45475
rect 23474 45472 23480 45484
rect 23247 45444 23480 45472
rect 23247 45441 23259 45444
rect 23201 45435 23259 45441
rect 23474 45432 23480 45444
rect 23532 45432 23538 45484
rect 23569 45475 23627 45481
rect 23569 45441 23581 45475
rect 23615 45472 23627 45475
rect 24026 45472 24032 45484
rect 23615 45444 24032 45472
rect 23615 45441 23627 45444
rect 23569 45435 23627 45441
rect 24026 45432 24032 45444
rect 24084 45432 24090 45484
rect 25406 45432 25412 45484
rect 25464 45472 25470 45484
rect 25777 45475 25835 45481
rect 25777 45472 25789 45475
rect 25464 45444 25789 45472
rect 25464 45432 25470 45444
rect 25777 45441 25789 45444
rect 25823 45441 25835 45475
rect 27157 45475 27215 45481
rect 27157 45472 27169 45475
rect 25777 45435 25835 45441
rect 25884 45444 27169 45472
rect 25593 45407 25651 45413
rect 25593 45404 25605 45407
rect 23124 45376 25605 45404
rect 23017 45367 23075 45373
rect 25593 45373 25605 45376
rect 25639 45373 25651 45407
rect 25593 45367 25651 45373
rect 19334 45296 19340 45348
rect 19392 45336 19398 45348
rect 19429 45339 19487 45345
rect 19429 45336 19441 45339
rect 19392 45308 19441 45336
rect 19392 45296 19398 45308
rect 19429 45305 19441 45308
rect 19475 45305 19487 45339
rect 19429 45299 19487 45305
rect 21177 45339 21235 45345
rect 21177 45305 21189 45339
rect 21223 45336 21235 45339
rect 22554 45336 22560 45348
rect 21223 45308 22560 45336
rect 21223 45305 21235 45308
rect 21177 45299 21235 45305
rect 22554 45296 22560 45308
rect 22612 45296 22618 45348
rect 23032 45336 23060 45367
rect 23658 45336 23664 45348
rect 23032 45308 23664 45336
rect 23658 45296 23664 45308
rect 23716 45296 23722 45348
rect 25314 45296 25320 45348
rect 25372 45336 25378 45348
rect 25884 45336 25912 45444
rect 27157 45441 27169 45444
rect 27203 45441 27215 45475
rect 28442 45472 28448 45484
rect 28403 45444 28448 45472
rect 27157 45435 27215 45441
rect 28442 45432 28448 45444
rect 28500 45432 28506 45484
rect 28736 45481 28764 45512
rect 30006 45500 30012 45512
rect 30064 45500 30070 45552
rect 30193 45543 30251 45549
rect 30193 45509 30205 45543
rect 30239 45540 30251 45543
rect 31294 45540 31300 45552
rect 30239 45512 31300 45540
rect 30239 45509 30251 45512
rect 30193 45503 30251 45509
rect 31294 45500 31300 45512
rect 31352 45500 31358 45552
rect 33318 45540 33324 45552
rect 32416 45512 33324 45540
rect 28721 45475 28779 45481
rect 28721 45441 28733 45475
rect 28767 45441 28779 45475
rect 28721 45435 28779 45441
rect 29733 45475 29791 45481
rect 29733 45441 29745 45475
rect 29779 45472 29791 45475
rect 29914 45472 29920 45484
rect 29779 45444 29920 45472
rect 29779 45441 29791 45444
rect 29733 45435 29791 45441
rect 29914 45432 29920 45444
rect 29972 45472 29978 45484
rect 30282 45472 30288 45484
rect 29972 45444 30288 45472
rect 29972 45432 29978 45444
rect 30282 45432 30288 45444
rect 30340 45432 30346 45484
rect 31021 45475 31079 45481
rect 31021 45441 31033 45475
rect 31067 45472 31079 45475
rect 31846 45472 31852 45484
rect 31067 45444 31852 45472
rect 31067 45441 31079 45444
rect 31021 45435 31079 45441
rect 31846 45432 31852 45444
rect 31904 45432 31910 45484
rect 32030 45432 32036 45484
rect 32088 45472 32094 45484
rect 32306 45472 32312 45484
rect 32088 45444 32312 45472
rect 32088 45432 32094 45444
rect 32306 45432 32312 45444
rect 32364 45432 32370 45484
rect 32416 45481 32444 45512
rect 33318 45500 33324 45512
rect 33376 45500 33382 45552
rect 33594 45540 33600 45552
rect 33555 45512 33600 45540
rect 33594 45500 33600 45512
rect 33652 45500 33658 45552
rect 34054 45540 34060 45552
rect 34015 45512 34060 45540
rect 34054 45500 34060 45512
rect 34112 45500 34118 45552
rect 34238 45500 34244 45552
rect 34296 45540 34302 45552
rect 38841 45543 38899 45549
rect 38841 45540 38853 45543
rect 34296 45512 36400 45540
rect 34296 45500 34302 45512
rect 32401 45475 32459 45481
rect 32401 45441 32413 45475
rect 32447 45441 32459 45475
rect 32582 45472 32588 45484
rect 32543 45444 32588 45472
rect 32401 45435 32459 45441
rect 32582 45432 32588 45444
rect 32640 45432 32646 45484
rect 32677 45475 32735 45481
rect 32677 45441 32689 45475
rect 32723 45472 32735 45475
rect 33134 45472 33140 45484
rect 32723 45444 33140 45472
rect 32723 45441 32735 45444
rect 32677 45435 32735 45441
rect 33134 45432 33140 45444
rect 33192 45432 33198 45484
rect 33941 45475 33999 45481
rect 33941 45441 33953 45475
rect 33987 45472 33999 45475
rect 34330 45472 34336 45484
rect 33987 45444 34336 45472
rect 33987 45441 33999 45444
rect 33941 45435 33999 45441
rect 34330 45432 34336 45444
rect 34388 45432 34394 45484
rect 35176 45481 35204 45512
rect 35161 45475 35219 45481
rect 35161 45441 35173 45475
rect 35207 45441 35219 45475
rect 35161 45435 35219 45441
rect 36139 45475 36197 45481
rect 36139 45441 36151 45475
rect 36185 45472 36197 45475
rect 36262 45472 36268 45484
rect 36185 45444 36268 45472
rect 36185 45441 36197 45444
rect 36139 45435 36197 45441
rect 36262 45432 36268 45444
rect 36320 45432 36326 45484
rect 26036 45407 26094 45413
rect 26036 45373 26048 45407
rect 26082 45404 26094 45407
rect 26329 45407 26387 45413
rect 26082 45376 26280 45404
rect 26082 45373 26094 45376
rect 26036 45367 26094 45373
rect 25372 45308 25912 45336
rect 26252 45336 26280 45376
rect 26329 45373 26341 45407
rect 26375 45404 26387 45407
rect 27982 45404 27988 45416
rect 26375 45376 27988 45404
rect 26375 45373 26387 45376
rect 26329 45367 26387 45373
rect 27982 45364 27988 45376
rect 28040 45364 28046 45416
rect 28077 45407 28135 45413
rect 28077 45373 28089 45407
rect 28123 45373 28135 45407
rect 28077 45367 28135 45373
rect 31113 45407 31171 45413
rect 31113 45373 31125 45407
rect 31159 45404 31171 45407
rect 32858 45404 32864 45416
rect 31159 45376 32864 45404
rect 31159 45373 31171 45376
rect 31113 45367 31171 45373
rect 27525 45339 27583 45345
rect 27525 45336 27537 45339
rect 26252 45308 27537 45336
rect 25372 45296 25378 45308
rect 27525 45305 27537 45308
rect 27571 45305 27583 45339
rect 27525 45299 27583 45305
rect 18693 45271 18751 45277
rect 18693 45268 18705 45271
rect 2832 45240 18705 45268
rect 2832 45228 2838 45240
rect 18693 45237 18705 45240
rect 18739 45237 18751 45271
rect 18693 45231 18751 45237
rect 22002 45228 22008 45280
rect 22060 45268 22066 45280
rect 22097 45271 22155 45277
rect 22097 45268 22109 45271
rect 22060 45240 22109 45268
rect 22060 45228 22066 45240
rect 22097 45237 22109 45240
rect 22143 45237 22155 45271
rect 22097 45231 22155 45237
rect 25498 45228 25504 45280
rect 25556 45268 25562 45280
rect 28092 45268 28120 45367
rect 32858 45364 32864 45376
rect 32916 45364 32922 45416
rect 33686 45364 33692 45416
rect 33744 45404 33750 45416
rect 33853 45407 33911 45413
rect 33853 45404 33865 45407
rect 33744 45376 33865 45404
rect 33744 45364 33750 45376
rect 33853 45373 33865 45376
rect 33899 45373 33911 45407
rect 33853 45367 33911 45373
rect 34149 45407 34207 45413
rect 34149 45373 34161 45407
rect 34195 45404 34207 45407
rect 34514 45404 34520 45416
rect 34195 45376 34520 45404
rect 34195 45373 34207 45376
rect 34149 45367 34207 45373
rect 34514 45364 34520 45376
rect 34572 45364 34578 45416
rect 31754 45296 31760 45348
rect 31812 45336 31818 45348
rect 32950 45336 32956 45348
rect 31812 45308 32956 45336
rect 31812 45296 31818 45308
rect 32950 45296 32956 45308
rect 33008 45296 33014 45348
rect 35802 45296 35808 45348
rect 35860 45336 35866 45348
rect 36280 45336 36308 45432
rect 36372 45404 36400 45512
rect 37568 45512 38853 45540
rect 36538 45472 36544 45484
rect 36451 45444 36544 45472
rect 36538 45432 36544 45444
rect 36596 45472 36602 45484
rect 37568 45481 37596 45512
rect 38841 45509 38853 45512
rect 38887 45540 38899 45543
rect 39206 45540 39212 45552
rect 38887 45512 39212 45540
rect 38887 45509 38899 45512
rect 38841 45503 38899 45509
rect 39206 45500 39212 45512
rect 39264 45500 39270 45552
rect 37553 45475 37611 45481
rect 37553 45472 37565 45475
rect 36596 45444 37565 45472
rect 36596 45432 36602 45444
rect 37553 45441 37565 45444
rect 37599 45441 37611 45475
rect 37553 45435 37611 45441
rect 37642 45432 37648 45484
rect 37700 45472 37706 45484
rect 37829 45475 37887 45481
rect 37700 45444 37745 45472
rect 37700 45432 37706 45444
rect 37829 45441 37841 45475
rect 37875 45472 37887 45475
rect 37918 45472 37924 45484
rect 37875 45444 37924 45472
rect 37875 45441 37887 45444
rect 37829 45435 37887 45441
rect 37918 45432 37924 45444
rect 37976 45472 37982 45484
rect 39022 45472 39028 45484
rect 37976 45444 38884 45472
rect 38983 45444 39028 45472
rect 37976 45432 37982 45444
rect 36446 45404 36452 45416
rect 36372 45376 36452 45404
rect 36446 45364 36452 45376
rect 36504 45404 36510 45416
rect 37274 45404 37280 45416
rect 36504 45376 37280 45404
rect 36504 45364 36510 45376
rect 37274 45364 37280 45376
rect 37332 45404 37338 45416
rect 37733 45407 37791 45413
rect 37733 45404 37745 45407
rect 37332 45376 37745 45404
rect 37332 45364 37338 45376
rect 37733 45373 37745 45376
rect 37779 45404 37791 45407
rect 38010 45404 38016 45416
rect 37779 45376 38016 45404
rect 37779 45373 37791 45376
rect 37733 45367 37791 45373
rect 38010 45364 38016 45376
rect 38068 45364 38074 45416
rect 38749 45407 38807 45413
rect 38749 45373 38761 45407
rect 38795 45373 38807 45407
rect 38856 45404 38884 45444
rect 39022 45432 39028 45444
rect 39080 45432 39086 45484
rect 39592 45481 39620 45580
rect 41432 45580 43812 45608
rect 39577 45475 39635 45481
rect 39577 45441 39589 45475
rect 39623 45441 39635 45475
rect 39577 45435 39635 45441
rect 39758 45404 39764 45416
rect 38856 45376 39764 45404
rect 38749 45367 38807 45373
rect 37642 45336 37648 45348
rect 35860 45308 37648 45336
rect 35860 45296 35866 45308
rect 37642 45296 37648 45308
rect 37700 45296 37706 45348
rect 38764 45336 38792 45367
rect 39758 45364 39764 45376
rect 39816 45364 39822 45416
rect 41432 45404 41460 45580
rect 43806 45568 43812 45580
rect 43864 45568 43870 45620
rect 41340 45376 41460 45404
rect 38930 45336 38936 45348
rect 38764 45308 38936 45336
rect 38930 45296 38936 45308
rect 38988 45336 38994 45348
rect 39942 45336 39948 45348
rect 38988 45308 39948 45336
rect 38988 45296 38994 45308
rect 39942 45296 39948 45308
rect 40000 45336 40006 45348
rect 41340 45345 41368 45376
rect 40221 45339 40279 45345
rect 40221 45336 40233 45339
rect 40000 45308 40233 45336
rect 40000 45296 40006 45308
rect 40221 45305 40233 45308
rect 40267 45336 40279 45339
rect 40773 45339 40831 45345
rect 40773 45336 40785 45339
rect 40267 45308 40785 45336
rect 40267 45305 40279 45308
rect 40221 45299 40279 45305
rect 40773 45305 40785 45308
rect 40819 45336 40831 45339
rect 41325 45339 41383 45345
rect 41325 45336 41337 45339
rect 40819 45308 41337 45336
rect 40819 45305 40831 45308
rect 40773 45299 40831 45305
rect 41325 45305 41337 45308
rect 41371 45305 41383 45339
rect 41325 45299 41383 45305
rect 33410 45268 33416 45280
rect 25556 45240 28120 45268
rect 33371 45240 33416 45268
rect 25556 45228 25562 45240
rect 33410 45228 33416 45240
rect 33468 45228 33474 45280
rect 34606 45228 34612 45280
rect 34664 45268 34670 45280
rect 34701 45271 34759 45277
rect 34701 45268 34713 45271
rect 34664 45240 34713 45268
rect 34664 45228 34670 45240
rect 34701 45237 34713 45240
rect 34747 45237 34759 45271
rect 34701 45231 34759 45237
rect 34790 45228 34796 45280
rect 34848 45268 34854 45280
rect 34885 45271 34943 45277
rect 34885 45268 34897 45271
rect 34848 45240 34897 45268
rect 34848 45228 34854 45240
rect 34885 45237 34897 45240
rect 34931 45237 34943 45271
rect 35986 45268 35992 45280
rect 35947 45240 35992 45268
rect 34885 45231 34943 45237
rect 35986 45228 35992 45240
rect 36044 45228 36050 45280
rect 41966 45268 41972 45280
rect 41879 45240 41972 45268
rect 41966 45228 41972 45240
rect 42024 45268 42030 45280
rect 42613 45271 42671 45277
rect 42613 45268 42625 45271
rect 42024 45240 42625 45268
rect 42024 45228 42030 45240
rect 42613 45237 42625 45240
rect 42659 45237 42671 45271
rect 42613 45231 42671 45237
rect 1104 45178 48852 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 48852 45178
rect 1104 45104 48852 45126
rect 17954 45024 17960 45076
rect 18012 45064 18018 45076
rect 18785 45067 18843 45073
rect 18785 45064 18797 45067
rect 18012 45036 18797 45064
rect 18012 45024 18018 45036
rect 18785 45033 18797 45036
rect 18831 45064 18843 45067
rect 20162 45064 20168 45076
rect 18831 45036 20168 45064
rect 18831 45033 18843 45036
rect 18785 45027 18843 45033
rect 20162 45024 20168 45036
rect 20220 45024 20226 45076
rect 21821 45067 21879 45073
rect 21821 45033 21833 45067
rect 21867 45064 21879 45067
rect 22554 45064 22560 45076
rect 21867 45036 22560 45064
rect 21867 45033 21879 45036
rect 21821 45027 21879 45033
rect 22554 45024 22560 45036
rect 22612 45024 22618 45076
rect 24762 45024 24768 45076
rect 24820 45064 24826 45076
rect 25961 45067 26019 45073
rect 25961 45064 25973 45067
rect 24820 45036 25973 45064
rect 24820 45024 24826 45036
rect 25961 45033 25973 45036
rect 26007 45033 26019 45067
rect 27154 45064 27160 45076
rect 27115 45036 27160 45064
rect 25961 45027 26019 45033
rect 27154 45024 27160 45036
rect 27212 45024 27218 45076
rect 27982 45064 27988 45076
rect 27264 45036 27988 45064
rect 23566 44996 23572 45008
rect 23527 44968 23572 44996
rect 23566 44956 23572 44968
rect 23624 44956 23630 45008
rect 23658 44956 23664 45008
rect 23716 44996 23722 45008
rect 25133 44999 25191 45005
rect 25133 44996 25145 44999
rect 23716 44968 25145 44996
rect 23716 44956 23722 44968
rect 25133 44965 25145 44968
rect 25179 44965 25191 44999
rect 25133 44959 25191 44965
rect 20806 44928 20812 44940
rect 20719 44900 20812 44928
rect 19794 44860 19800 44872
rect 19755 44832 19800 44860
rect 19794 44820 19800 44832
rect 19852 44860 19858 44872
rect 19978 44860 19984 44872
rect 19852 44832 19984 44860
rect 19852 44820 19858 44832
rect 19978 44820 19984 44832
rect 20036 44860 20042 44872
rect 20732 44869 20760 44900
rect 20806 44888 20812 44900
rect 20864 44928 20870 44940
rect 27264 44928 27292 45036
rect 27982 45024 27988 45036
rect 28040 45024 28046 45076
rect 28166 45024 28172 45076
rect 28224 45064 28230 45076
rect 28997 45067 29055 45073
rect 28997 45064 29009 45067
rect 28224 45036 29009 45064
rect 28224 45024 28230 45036
rect 28997 45033 29009 45036
rect 29043 45033 29055 45067
rect 28997 45027 29055 45033
rect 29546 45024 29552 45076
rect 29604 45064 29610 45076
rect 30745 45067 30803 45073
rect 30745 45064 30757 45067
rect 29604 45036 30757 45064
rect 29604 45024 29610 45036
rect 30745 45033 30757 45036
rect 30791 45033 30803 45067
rect 30745 45027 30803 45033
rect 31757 45067 31815 45073
rect 31757 45033 31769 45067
rect 31803 45064 31815 45067
rect 32306 45064 32312 45076
rect 31803 45036 32312 45064
rect 31803 45033 31815 45036
rect 31757 45027 31815 45033
rect 32306 45024 32312 45036
rect 32364 45024 32370 45076
rect 34146 45064 34152 45076
rect 34107 45036 34152 45064
rect 34146 45024 34152 45036
rect 34204 45024 34210 45076
rect 34977 45067 35035 45073
rect 34977 45033 34989 45067
rect 35023 45064 35035 45067
rect 35710 45064 35716 45076
rect 35023 45036 35716 45064
rect 35023 45033 35035 45036
rect 34977 45027 35035 45033
rect 35710 45024 35716 45036
rect 35768 45024 35774 45076
rect 35820 45036 36584 45064
rect 29086 44996 29092 45008
rect 20864 44900 27292 44928
rect 27632 44968 29092 44996
rect 20864 44888 20870 44900
rect 20533 44863 20591 44869
rect 20533 44860 20545 44863
rect 20036 44832 20545 44860
rect 20036 44820 20042 44832
rect 20533 44829 20545 44832
rect 20579 44829 20591 44863
rect 20533 44823 20591 44829
rect 20717 44863 20775 44869
rect 20717 44829 20729 44863
rect 20763 44829 20775 44863
rect 22002 44860 22008 44872
rect 21963 44832 22008 44860
rect 20717 44823 20775 44829
rect 22002 44820 22008 44832
rect 22060 44820 22066 44872
rect 22649 44863 22707 44869
rect 22649 44829 22661 44863
rect 22695 44829 22707 44863
rect 22649 44823 22707 44829
rect 22833 44863 22891 44869
rect 22833 44829 22845 44863
rect 22879 44860 22891 44863
rect 24394 44860 24400 44872
rect 22879 44832 24400 44860
rect 22879 44829 22891 44832
rect 22833 44823 22891 44829
rect 22664 44792 22692 44823
rect 24394 44820 24400 44832
rect 24452 44820 24458 44872
rect 24578 44860 24584 44872
rect 24539 44832 24584 44860
rect 24578 44820 24584 44832
rect 24636 44820 24642 44872
rect 24670 44820 24676 44872
rect 24728 44860 24734 44872
rect 24857 44863 24915 44869
rect 24728 44832 24773 44860
rect 24728 44820 24734 44832
rect 24857 44829 24869 44863
rect 24903 44829 24915 44863
rect 24857 44823 24915 44829
rect 24949 44863 25007 44869
rect 24949 44829 24961 44863
rect 24995 44860 25007 44863
rect 25314 44860 25320 44872
rect 24995 44832 25320 44860
rect 24995 44829 25007 44832
rect 24949 44823 25007 44829
rect 23845 44795 23903 44801
rect 22664 44764 23520 44792
rect 19981 44727 20039 44733
rect 19981 44693 19993 44727
rect 20027 44724 20039 44727
rect 20162 44724 20168 44736
rect 20027 44696 20168 44724
rect 20027 44693 20039 44696
rect 19981 44687 20039 44693
rect 20162 44684 20168 44696
rect 20220 44724 20226 44736
rect 20438 44724 20444 44736
rect 20220 44696 20444 44724
rect 20220 44684 20226 44696
rect 20438 44684 20444 44696
rect 20496 44684 20502 44736
rect 20806 44684 20812 44736
rect 20864 44724 20870 44736
rect 20901 44727 20959 44733
rect 20901 44724 20913 44727
rect 20864 44696 20913 44724
rect 20864 44684 20870 44696
rect 20901 44693 20913 44696
rect 20947 44693 20959 44727
rect 22738 44724 22744 44736
rect 22699 44696 22744 44724
rect 20901 44687 20959 44693
rect 22738 44684 22744 44696
rect 22796 44684 22802 44736
rect 23382 44724 23388 44736
rect 23343 44696 23388 44724
rect 23382 44684 23388 44696
rect 23440 44684 23446 44736
rect 23492 44724 23520 44764
rect 23845 44761 23857 44795
rect 23891 44792 23903 44795
rect 24688 44792 24716 44820
rect 23891 44764 24716 44792
rect 23891 44761 23903 44764
rect 23845 44755 23903 44761
rect 24762 44752 24768 44804
rect 24820 44792 24826 44804
rect 24872 44792 24900 44823
rect 25314 44820 25320 44832
rect 25372 44820 25378 44872
rect 25869 44863 25927 44869
rect 25869 44829 25881 44863
rect 25915 44860 25927 44863
rect 25958 44860 25964 44872
rect 25915 44832 25964 44860
rect 25915 44829 25927 44832
rect 25869 44823 25927 44829
rect 25958 44820 25964 44832
rect 26016 44860 26022 44872
rect 27338 44860 27344 44872
rect 26016 44832 27344 44860
rect 26016 44820 26022 44832
rect 27338 44820 27344 44832
rect 27396 44820 27402 44872
rect 27632 44869 27660 44968
rect 29086 44956 29092 44968
rect 29144 44996 29150 45008
rect 29825 44999 29883 45005
rect 29825 44996 29837 44999
rect 29144 44968 29837 44996
rect 29144 44956 29150 44968
rect 29825 44965 29837 44968
rect 29871 44965 29883 44999
rect 33410 44996 33416 45008
rect 29825 44959 29883 44965
rect 31726 44968 33416 44996
rect 27982 44888 27988 44940
rect 28040 44928 28046 44940
rect 31726 44928 31754 44968
rect 33410 44956 33416 44968
rect 33468 44956 33474 45008
rect 35820 44996 35848 45036
rect 36446 44996 36452 45008
rect 33520 44968 35848 44996
rect 36004 44968 36452 44996
rect 32490 44928 32496 44940
rect 28040 44900 31754 44928
rect 31956 44900 32496 44928
rect 28040 44888 28046 44900
rect 27617 44863 27675 44869
rect 27617 44829 27629 44863
rect 27663 44829 27675 44863
rect 27617 44823 27675 44829
rect 27706 44820 27712 44872
rect 27764 44860 27770 44872
rect 28074 44860 28080 44872
rect 27764 44832 27809 44860
rect 28035 44832 28080 44860
rect 27764 44820 27770 44832
rect 28074 44820 28080 44832
rect 28132 44820 28138 44872
rect 28721 44863 28779 44869
rect 28721 44860 28733 44863
rect 28184 44832 28733 44860
rect 24820 44764 24900 44792
rect 24820 44752 24826 44764
rect 26418 44752 26424 44804
rect 26476 44792 26482 44804
rect 27430 44792 27436 44804
rect 26476 44764 27436 44792
rect 26476 44752 26482 44764
rect 27430 44752 27436 44764
rect 27488 44792 27494 44804
rect 28184 44792 28212 44832
rect 28721 44829 28733 44832
rect 28767 44829 28779 44863
rect 29914 44860 29920 44872
rect 29875 44832 29920 44860
rect 28721 44823 28779 44829
rect 29914 44820 29920 44832
rect 29972 44820 29978 44872
rect 30190 44860 30196 44872
rect 30151 44832 30196 44860
rect 30190 44820 30196 44832
rect 30248 44860 30254 44872
rect 31294 44860 31300 44872
rect 30248 44832 31300 44860
rect 30248 44820 30254 44832
rect 31294 44820 31300 44832
rect 31352 44820 31358 44872
rect 31956 44869 31984 44900
rect 32490 44888 32496 44900
rect 32548 44928 32554 44940
rect 33520 44928 33548 44968
rect 32548 44900 33548 44928
rect 32548 44888 32554 44900
rect 31941 44863 31999 44869
rect 31941 44829 31953 44863
rect 31987 44829 31999 44863
rect 31941 44823 31999 44829
rect 32125 44863 32183 44869
rect 32125 44829 32137 44863
rect 32171 44860 32183 44863
rect 32674 44860 32680 44872
rect 32171 44832 32680 44860
rect 32171 44829 32183 44832
rect 32125 44823 32183 44829
rect 32674 44820 32680 44832
rect 32732 44820 32738 44872
rect 33520 44860 33548 44900
rect 33689 44931 33747 44937
rect 33689 44897 33701 44931
rect 33735 44928 33747 44931
rect 33962 44928 33968 44940
rect 33735 44900 33968 44928
rect 33735 44897 33747 44900
rect 33689 44891 33747 44897
rect 33962 44888 33968 44900
rect 34020 44888 34026 44940
rect 33350 44832 33548 44860
rect 34330 44820 34336 44872
rect 34388 44860 34394 44872
rect 35069 44863 35127 44869
rect 35069 44860 35081 44863
rect 34388 44832 35081 44860
rect 34388 44820 34394 44832
rect 35069 44829 35081 44832
rect 35115 44829 35127 44863
rect 35069 44823 35127 44829
rect 35713 44863 35771 44869
rect 35713 44829 35725 44863
rect 35759 44860 35771 44863
rect 35802 44860 35808 44872
rect 35759 44832 35808 44860
rect 35759 44829 35771 44832
rect 35713 44823 35771 44829
rect 27488 44764 28212 44792
rect 28261 44795 28319 44801
rect 27488 44752 27494 44764
rect 28261 44761 28273 44795
rect 28307 44792 28319 44795
rect 28534 44792 28540 44804
rect 28307 44764 28540 44792
rect 28307 44761 28319 44764
rect 28261 44755 28319 44761
rect 28534 44752 28540 44764
rect 28592 44792 28598 44804
rect 28997 44795 29055 44801
rect 28997 44792 29009 44795
rect 28592 44764 29009 44792
rect 28592 44752 28598 44764
rect 28997 44761 29009 44764
rect 29043 44761 29055 44795
rect 28997 44755 29055 44761
rect 29181 44795 29239 44801
rect 29181 44761 29193 44795
rect 29227 44792 29239 44795
rect 29362 44792 29368 44804
rect 29227 44764 29368 44792
rect 29227 44761 29239 44764
rect 29181 44755 29239 44761
rect 29362 44752 29368 44764
rect 29420 44752 29426 44804
rect 24302 44724 24308 44736
rect 23492 44696 24308 44724
rect 24302 44684 24308 44696
rect 24360 44684 24366 44736
rect 26329 44727 26387 44733
rect 26329 44693 26341 44727
rect 26375 44724 26387 44727
rect 26602 44724 26608 44736
rect 26375 44696 26608 44724
rect 26375 44693 26387 44696
rect 26329 44687 26387 44693
rect 26602 44684 26608 44696
rect 26660 44684 26666 44736
rect 35084 44724 35112 44823
rect 35802 44820 35808 44832
rect 35860 44820 35866 44872
rect 35897 44863 35955 44869
rect 35897 44829 35909 44863
rect 35943 44860 35955 44863
rect 36004 44860 36032 44968
rect 36446 44956 36452 44968
rect 36504 44956 36510 45008
rect 36354 44928 36360 44940
rect 36315 44900 36360 44928
rect 36354 44888 36360 44900
rect 36412 44888 36418 44940
rect 36556 44928 36584 45036
rect 37826 45024 37832 45076
rect 37884 45064 37890 45076
rect 38381 45067 38439 45073
rect 38381 45064 38393 45067
rect 37884 45036 38393 45064
rect 37884 45024 37890 45036
rect 38381 45033 38393 45036
rect 38427 45033 38439 45067
rect 38381 45027 38439 45033
rect 39758 45024 39764 45076
rect 39816 45064 39822 45076
rect 40589 45067 40647 45073
rect 40589 45064 40601 45067
rect 39816 45036 40601 45064
rect 39816 45024 39822 45036
rect 40589 45033 40601 45036
rect 40635 45064 40647 45067
rect 41141 45067 41199 45073
rect 41141 45064 41153 45067
rect 40635 45036 41153 45064
rect 40635 45033 40647 45036
rect 40589 45027 40647 45033
rect 41141 45033 41153 45036
rect 41187 45033 41199 45067
rect 41141 45027 41199 45033
rect 41230 45024 41236 45076
rect 41288 45064 41294 45076
rect 41785 45067 41843 45073
rect 41785 45064 41797 45067
rect 41288 45036 41797 45064
rect 41288 45024 41294 45036
rect 41785 45033 41797 45036
rect 41831 45064 41843 45067
rect 44174 45064 44180 45076
rect 41831 45036 44180 45064
rect 41831 45033 41843 45036
rect 41785 45027 41843 45033
rect 44174 45024 44180 45036
rect 44232 45024 44238 45076
rect 39117 44999 39175 45005
rect 39117 44965 39129 44999
rect 39163 44996 39175 44999
rect 40218 44996 40224 45008
rect 39163 44968 40224 44996
rect 39163 44965 39175 44968
rect 39117 44959 39175 44965
rect 40218 44956 40224 44968
rect 40276 44956 40282 45008
rect 36817 44931 36875 44937
rect 36817 44928 36829 44931
rect 36556 44900 36829 44928
rect 36817 44897 36829 44900
rect 36863 44897 36875 44931
rect 37550 44928 37556 44940
rect 37511 44900 37556 44928
rect 36817 44891 36875 44897
rect 37550 44888 37556 44900
rect 37608 44888 37614 44940
rect 37642 44888 37648 44940
rect 37700 44928 37706 44940
rect 41966 44928 41972 44940
rect 37700 44900 41972 44928
rect 37700 44888 37706 44900
rect 41966 44888 41972 44900
rect 42024 44888 42030 44940
rect 35943 44832 36032 44860
rect 36173 44863 36231 44869
rect 35943 44829 35955 44832
rect 35897 44823 35955 44829
rect 36173 44829 36185 44863
rect 36219 44860 36231 44863
rect 36538 44860 36544 44872
rect 36219 44832 36544 44860
rect 36219 44829 36231 44832
rect 36173 44823 36231 44829
rect 36538 44820 36544 44832
rect 36596 44820 36602 44872
rect 37458 44860 37464 44872
rect 37371 44832 37464 44860
rect 37458 44820 37464 44832
rect 37516 44860 37522 44872
rect 37918 44860 37924 44872
rect 37516 44832 37924 44860
rect 37516 44820 37522 44832
rect 37918 44820 37924 44832
rect 37976 44820 37982 44872
rect 35434 44752 35440 44804
rect 35492 44792 35498 44804
rect 40037 44795 40095 44801
rect 40037 44792 40049 44795
rect 35492 44764 40049 44792
rect 35492 44752 35498 44764
rect 40037 44761 40049 44764
rect 40083 44761 40095 44795
rect 40037 44755 40095 44761
rect 38102 44724 38108 44736
rect 35084 44696 38108 44724
rect 38102 44684 38108 44696
rect 38160 44684 38166 44736
rect 1104 44634 48852 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 48852 44634
rect 1104 44560 48852 44582
rect 19705 44523 19763 44529
rect 19705 44489 19717 44523
rect 19751 44520 19763 44523
rect 19978 44520 19984 44532
rect 19751 44492 19984 44520
rect 19751 44489 19763 44492
rect 19705 44483 19763 44489
rect 19978 44480 19984 44492
rect 20036 44520 20042 44532
rect 20257 44523 20315 44529
rect 20257 44520 20269 44523
rect 20036 44492 20269 44520
rect 20036 44480 20042 44492
rect 20257 44489 20269 44492
rect 20303 44489 20315 44523
rect 20257 44483 20315 44489
rect 20530 44480 20536 44532
rect 20588 44520 20594 44532
rect 20993 44523 21051 44529
rect 20993 44520 21005 44523
rect 20588 44492 21005 44520
rect 20588 44480 20594 44492
rect 20993 44489 21005 44492
rect 21039 44489 21051 44523
rect 23198 44520 23204 44532
rect 23159 44492 23204 44520
rect 20993 44483 21051 44489
rect 23198 44480 23204 44492
rect 23256 44480 23262 44532
rect 25406 44520 25412 44532
rect 25367 44492 25412 44520
rect 25406 44480 25412 44492
rect 25464 44480 25470 44532
rect 25498 44480 25504 44532
rect 25556 44520 25562 44532
rect 28629 44523 28687 44529
rect 28629 44520 28641 44523
rect 25556 44492 28641 44520
rect 25556 44480 25562 44492
rect 28629 44489 28641 44492
rect 28675 44489 28687 44523
rect 30374 44520 30380 44532
rect 28629 44483 28687 44489
rect 29288 44492 30380 44520
rect 22097 44455 22155 44461
rect 22097 44421 22109 44455
rect 22143 44452 22155 44455
rect 22370 44452 22376 44464
rect 22143 44424 22376 44452
rect 22143 44421 22155 44424
rect 22097 44415 22155 44421
rect 22370 44412 22376 44424
rect 22428 44452 22434 44464
rect 26142 44452 26148 44464
rect 22428 44424 26148 44452
rect 22428 44412 22434 44424
rect 26142 44412 26148 44424
rect 26200 44412 26206 44464
rect 26513 44455 26571 44461
rect 26513 44421 26525 44455
rect 26559 44421 26571 44455
rect 28074 44452 28080 44464
rect 26513 44415 26571 44421
rect 27540 44424 28080 44452
rect 20806 44384 20812 44396
rect 20767 44356 20812 44384
rect 20806 44344 20812 44356
rect 20864 44344 20870 44396
rect 23382 44344 23388 44396
rect 23440 44384 23446 44396
rect 23569 44387 23627 44393
rect 23569 44384 23581 44387
rect 23440 44356 23581 44384
rect 23440 44344 23446 44356
rect 23569 44353 23581 44356
rect 23615 44353 23627 44387
rect 23934 44384 23940 44396
rect 23895 44356 23940 44384
rect 23569 44347 23627 44353
rect 23934 44344 23940 44356
rect 23992 44344 23998 44396
rect 24854 44344 24860 44396
rect 24912 44384 24918 44396
rect 25041 44387 25099 44393
rect 25041 44384 25053 44387
rect 24912 44356 25053 44384
rect 24912 44344 24918 44356
rect 25041 44353 25053 44356
rect 25087 44353 25099 44387
rect 25041 44347 25099 44353
rect 25409 44387 25467 44393
rect 25409 44353 25421 44387
rect 25455 44384 25467 44387
rect 25866 44384 25872 44396
rect 25455 44356 25872 44384
rect 25455 44353 25467 44356
rect 25409 44347 25467 44353
rect 25866 44344 25872 44356
rect 25924 44344 25930 44396
rect 26329 44387 26387 44393
rect 26329 44353 26341 44387
rect 26375 44384 26387 44387
rect 26418 44384 26424 44396
rect 26375 44356 26424 44384
rect 26375 44353 26387 44356
rect 26329 44347 26387 44353
rect 26418 44344 26424 44356
rect 26476 44344 26482 44396
rect 25314 44276 25320 44328
rect 25372 44316 25378 44328
rect 25593 44319 25651 44325
rect 25593 44316 25605 44319
rect 25372 44288 25605 44316
rect 25372 44276 25378 44288
rect 25593 44285 25605 44288
rect 25639 44316 25651 44319
rect 25639 44288 26188 44316
rect 25639 44285 25651 44288
rect 25593 44279 25651 44285
rect 22741 44251 22799 44257
rect 22741 44217 22753 44251
rect 22787 44248 22799 44251
rect 24486 44248 24492 44260
rect 22787 44220 24492 44248
rect 22787 44217 22799 44220
rect 22741 44211 22799 44217
rect 24486 44208 24492 44220
rect 24544 44208 24550 44260
rect 26160 44257 26188 44288
rect 26145 44251 26203 44257
rect 26145 44217 26157 44251
rect 26191 44217 26203 44251
rect 26528 44248 26556 44415
rect 26602 44344 26608 44396
rect 26660 44384 26666 44396
rect 27540 44393 27568 44424
rect 28074 44412 28080 44424
rect 28132 44412 28138 44464
rect 28166 44412 28172 44464
rect 28224 44452 28230 44464
rect 28224 44424 28269 44452
rect 28224 44412 28230 44424
rect 27525 44387 27583 44393
rect 26660 44356 26705 44384
rect 26660 44344 26666 44356
rect 27525 44353 27537 44387
rect 27571 44353 27583 44387
rect 27525 44347 27583 44353
rect 27706 44344 27712 44396
rect 27764 44384 27770 44396
rect 29288 44393 29316 44492
rect 30374 44480 30380 44492
rect 30432 44520 30438 44532
rect 30926 44520 30932 44532
rect 30432 44492 30932 44520
rect 30432 44480 30438 44492
rect 30926 44480 30932 44492
rect 30984 44480 30990 44532
rect 32677 44523 32735 44529
rect 32677 44489 32689 44523
rect 32723 44520 32735 44523
rect 33318 44520 33324 44532
rect 32723 44492 33324 44520
rect 32723 44489 32735 44492
rect 32677 44483 32735 44489
rect 33318 44480 33324 44492
rect 33376 44480 33382 44532
rect 36173 44523 36231 44529
rect 36173 44489 36185 44523
rect 36219 44520 36231 44523
rect 36354 44520 36360 44532
rect 36219 44492 36360 44520
rect 36219 44489 36231 44492
rect 36173 44483 36231 44489
rect 36354 44480 36360 44492
rect 36412 44480 36418 44532
rect 37550 44520 37556 44532
rect 37511 44492 37556 44520
rect 37550 44480 37556 44492
rect 37608 44480 37614 44532
rect 37734 44480 37740 44532
rect 37792 44480 37798 44532
rect 38102 44480 38108 44532
rect 38160 44520 38166 44532
rect 38565 44523 38623 44529
rect 38565 44520 38577 44523
rect 38160 44492 38577 44520
rect 38160 44480 38166 44492
rect 38565 44489 38577 44492
rect 38611 44520 38623 44523
rect 39022 44520 39028 44532
rect 38611 44492 39028 44520
rect 38611 44489 38623 44492
rect 38565 44483 38623 44489
rect 39022 44480 39028 44492
rect 39080 44520 39086 44532
rect 40773 44523 40831 44529
rect 40773 44520 40785 44523
rect 39080 44492 40785 44520
rect 39080 44480 39086 44492
rect 40773 44489 40785 44492
rect 40819 44520 40831 44523
rect 41230 44520 41236 44532
rect 40819 44492 41236 44520
rect 40819 44489 40831 44492
rect 40773 44483 40831 44489
rect 41230 44480 41236 44492
rect 41288 44480 41294 44532
rect 30650 44412 30656 44464
rect 30708 44452 30714 44464
rect 30745 44455 30803 44461
rect 30745 44452 30757 44455
rect 30708 44424 30757 44452
rect 30708 44412 30714 44424
rect 30745 44421 30757 44424
rect 30791 44421 30803 44455
rect 30745 44415 30803 44421
rect 33134 44412 33140 44464
rect 33192 44452 33198 44464
rect 33597 44455 33655 44461
rect 33597 44452 33609 44455
rect 33192 44424 33609 44452
rect 33192 44412 33198 44424
rect 33597 44421 33609 44424
rect 33643 44421 33655 44455
rect 33597 44415 33655 44421
rect 33965 44455 34023 44461
rect 33965 44421 33977 44455
rect 34011 44452 34023 44455
rect 35434 44452 35440 44464
rect 34011 44424 35440 44452
rect 34011 44421 34023 44424
rect 33965 44415 34023 44421
rect 35434 44412 35440 44424
rect 35492 44412 35498 44464
rect 35986 44412 35992 44464
rect 36044 44452 36050 44464
rect 36081 44455 36139 44461
rect 36081 44452 36093 44455
rect 36044 44424 36093 44452
rect 36044 44412 36050 44424
rect 36081 44421 36093 44424
rect 36127 44421 36139 44455
rect 36906 44452 36912 44464
rect 36081 44415 36139 44421
rect 36372 44424 36912 44452
rect 27985 44387 28043 44393
rect 27764 44356 27857 44384
rect 27764 44344 27770 44356
rect 27985 44353 27997 44387
rect 28031 44353 28043 44387
rect 27985 44347 28043 44353
rect 29273 44387 29331 44393
rect 29273 44353 29285 44387
rect 29319 44353 29331 44387
rect 29638 44384 29644 44396
rect 29599 44356 29644 44384
rect 29273 44347 29331 44353
rect 27338 44276 27344 44328
rect 27396 44316 27402 44328
rect 27724 44316 27752 44344
rect 27396 44288 27752 44316
rect 28000 44316 28028 44347
rect 29638 44344 29644 44356
rect 29696 44344 29702 44396
rect 32493 44387 32551 44393
rect 32493 44353 32505 44387
rect 32539 44384 32551 44387
rect 32950 44384 32956 44396
rect 32539 44356 32956 44384
rect 32539 44353 32551 44356
rect 32493 44347 32551 44353
rect 32950 44344 32956 44356
rect 33008 44344 33014 44396
rect 33781 44387 33839 44393
rect 33781 44353 33793 44387
rect 33827 44353 33839 44387
rect 33781 44347 33839 44353
rect 34057 44387 34115 44393
rect 34057 44353 34069 44387
rect 34103 44384 34115 44387
rect 34606 44384 34612 44396
rect 34103 44356 34612 44384
rect 34103 44353 34115 44356
rect 34057 44347 34115 44353
rect 29086 44316 29092 44328
rect 28000 44288 29092 44316
rect 27396 44276 27402 44288
rect 29086 44276 29092 44288
rect 29144 44276 29150 44328
rect 30098 44276 30104 44328
rect 30156 44316 30162 44328
rect 30193 44319 30251 44325
rect 30193 44316 30205 44319
rect 30156 44288 30205 44316
rect 30156 44276 30162 44288
rect 30193 44285 30205 44288
rect 30239 44285 30251 44319
rect 30193 44279 30251 44285
rect 30837 44319 30895 44325
rect 30837 44285 30849 44319
rect 30883 44316 30895 44319
rect 31389 44319 31447 44325
rect 31389 44316 31401 44319
rect 30883 44288 31401 44316
rect 30883 44285 30895 44288
rect 30837 44279 30895 44285
rect 31389 44285 31401 44288
rect 31435 44285 31447 44319
rect 31389 44279 31447 44285
rect 32214 44276 32220 44328
rect 32272 44316 32278 44328
rect 32309 44319 32367 44325
rect 32309 44316 32321 44319
rect 32272 44288 32321 44316
rect 32272 44276 32278 44288
rect 32309 44285 32321 44288
rect 32355 44316 32367 44319
rect 33226 44316 33232 44328
rect 32355 44288 33232 44316
rect 32355 44285 32367 44288
rect 32309 44279 32367 44285
rect 33226 44276 33232 44288
rect 33284 44276 33290 44328
rect 33796 44316 33824 44347
rect 34606 44344 34612 44356
rect 34664 44344 34670 44396
rect 34790 44384 34796 44396
rect 34751 44356 34796 44384
rect 34790 44344 34796 44356
rect 34848 44344 34854 44396
rect 35621 44387 35679 44393
rect 35621 44353 35633 44387
rect 35667 44384 35679 44387
rect 36170 44384 36176 44396
rect 35667 44356 36176 44384
rect 35667 44353 35679 44356
rect 35621 44347 35679 44353
rect 36170 44344 36176 44356
rect 36228 44344 36234 44396
rect 36372 44393 36400 44424
rect 36906 44412 36912 44424
rect 36964 44452 36970 44464
rect 37752 44452 37780 44480
rect 36964 44424 37780 44452
rect 39117 44455 39175 44461
rect 36964 44412 36970 44424
rect 39117 44421 39129 44455
rect 39163 44452 39175 44455
rect 39669 44455 39727 44461
rect 39669 44452 39681 44455
rect 39163 44424 39681 44452
rect 39163 44421 39175 44424
rect 39117 44415 39175 44421
rect 39669 44421 39681 44424
rect 39715 44452 39727 44455
rect 40218 44452 40224 44464
rect 39715 44424 40224 44452
rect 39715 44421 39727 44424
rect 39669 44415 39727 44421
rect 36357 44387 36415 44393
rect 36357 44353 36369 44387
rect 36403 44353 36415 44387
rect 36357 44347 36415 44353
rect 36538 44344 36544 44396
rect 36596 44384 36602 44396
rect 37737 44387 37795 44393
rect 37737 44384 37749 44387
rect 36596 44356 37749 44384
rect 36596 44344 36602 44356
rect 37737 44353 37749 44356
rect 37783 44353 37795 44387
rect 38010 44384 38016 44396
rect 37923 44356 38016 44384
rect 37737 44347 37795 44353
rect 38010 44344 38016 44356
rect 38068 44384 38074 44396
rect 39132 44384 39160 44415
rect 40218 44412 40224 44424
rect 40276 44412 40282 44464
rect 38068 44356 39160 44384
rect 38068 44344 38074 44356
rect 35342 44316 35348 44328
rect 33796 44288 35348 44316
rect 35342 44276 35348 44288
rect 35400 44276 35406 44328
rect 37642 44276 37648 44328
rect 37700 44316 37706 44328
rect 37921 44319 37979 44325
rect 37921 44316 37933 44319
rect 37700 44288 37933 44316
rect 37700 44276 37706 44288
rect 37921 44285 37933 44288
rect 37967 44285 37979 44319
rect 37921 44279 37979 44285
rect 28074 44248 28080 44260
rect 26528 44220 28080 44248
rect 26145 44211 26203 44217
rect 28074 44208 28080 44220
rect 28132 44208 28138 44260
rect 35434 44140 35440 44192
rect 35492 44180 35498 44192
rect 36541 44183 36599 44189
rect 36541 44180 36553 44183
rect 35492 44152 36553 44180
rect 35492 44140 35498 44152
rect 36541 44149 36553 44152
rect 36587 44149 36599 44183
rect 36541 44143 36599 44149
rect 1104 44090 48852 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 48852 44090
rect 1104 44016 48852 44038
rect 22370 43976 22376 43988
rect 22331 43948 22376 43976
rect 22370 43936 22376 43948
rect 22428 43936 22434 43988
rect 23017 43979 23075 43985
rect 23017 43945 23029 43979
rect 23063 43976 23075 43979
rect 24210 43976 24216 43988
rect 23063 43948 24216 43976
rect 23063 43945 23075 43948
rect 23017 43939 23075 43945
rect 24210 43936 24216 43948
rect 24268 43936 24274 43988
rect 28074 43976 28080 43988
rect 28035 43948 28080 43976
rect 28074 43936 28080 43948
rect 28132 43936 28138 43988
rect 29178 43976 29184 43988
rect 29139 43948 29184 43976
rect 29178 43936 29184 43948
rect 29236 43936 29242 43988
rect 29638 43936 29644 43988
rect 29696 43976 29702 43988
rect 29825 43979 29883 43985
rect 29825 43976 29837 43979
rect 29696 43948 29837 43976
rect 29696 43936 29702 43948
rect 29825 43945 29837 43948
rect 29871 43945 29883 43979
rect 29825 43939 29883 43945
rect 30190 43936 30196 43988
rect 30248 43976 30254 43988
rect 30745 43979 30803 43985
rect 30745 43976 30757 43979
rect 30248 43948 30757 43976
rect 30248 43936 30254 43948
rect 30745 43945 30757 43948
rect 30791 43945 30803 43979
rect 31386 43976 31392 43988
rect 31347 43948 31392 43976
rect 30745 43939 30803 43945
rect 31386 43936 31392 43948
rect 31444 43936 31450 43988
rect 32309 43979 32367 43985
rect 32309 43945 32321 43979
rect 32355 43976 32367 43979
rect 32582 43976 32588 43988
rect 32355 43948 32588 43976
rect 32355 43945 32367 43948
rect 32309 43939 32367 43945
rect 32582 43936 32588 43948
rect 32640 43936 32646 43988
rect 33686 43976 33692 43988
rect 33647 43948 33692 43976
rect 33686 43936 33692 43948
rect 33744 43936 33750 43988
rect 34790 43936 34796 43988
rect 34848 43976 34854 43988
rect 34977 43979 35035 43985
rect 34977 43976 34989 43979
rect 34848 43948 34989 43976
rect 34848 43936 34854 43948
rect 34977 43945 34989 43948
rect 35023 43945 35035 43979
rect 35342 43976 35348 43988
rect 35303 43948 35348 43976
rect 34977 43939 35035 43945
rect 35342 43936 35348 43948
rect 35400 43976 35406 43988
rect 35989 43979 36047 43985
rect 35989 43976 36001 43979
rect 35400 43948 36001 43976
rect 35400 43936 35406 43948
rect 35989 43945 36001 43948
rect 36035 43945 36047 43979
rect 35989 43939 36047 43945
rect 36173 43979 36231 43985
rect 36173 43945 36185 43979
rect 36219 43976 36231 43979
rect 36354 43976 36360 43988
rect 36219 43948 36360 43976
rect 36219 43945 36231 43948
rect 36173 43939 36231 43945
rect 36354 43936 36360 43948
rect 36412 43936 36418 43988
rect 36906 43976 36912 43988
rect 36867 43948 36912 43976
rect 36906 43936 36912 43948
rect 36964 43936 36970 43988
rect 37642 43936 37648 43988
rect 37700 43976 37706 43988
rect 38473 43979 38531 43985
rect 38473 43976 38485 43979
rect 37700 43948 38485 43976
rect 37700 43936 37706 43948
rect 38473 43945 38485 43948
rect 38519 43976 38531 43979
rect 39025 43979 39083 43985
rect 39025 43976 39037 43979
rect 38519 43948 39037 43976
rect 38519 43945 38531 43948
rect 38473 43939 38531 43945
rect 39025 43945 39037 43948
rect 39071 43945 39083 43979
rect 39025 43939 39083 43945
rect 39942 43936 39948 43988
rect 40000 43976 40006 43988
rect 40037 43979 40095 43985
rect 40037 43976 40049 43979
rect 40000 43948 40049 43976
rect 40000 43936 40006 43948
rect 40037 43945 40049 43948
rect 40083 43976 40095 43979
rect 40589 43979 40647 43985
rect 40589 43976 40601 43979
rect 40083 43948 40601 43976
rect 40083 43945 40095 43948
rect 40037 43939 40095 43945
rect 40589 43945 40601 43948
rect 40635 43945 40647 43979
rect 40589 43939 40647 43945
rect 23934 43908 23940 43920
rect 23895 43880 23940 43908
rect 23934 43868 23940 43880
rect 23992 43868 23998 43920
rect 26694 43908 26700 43920
rect 25056 43880 26700 43908
rect 24029 43843 24087 43849
rect 24029 43809 24041 43843
rect 24075 43840 24087 43843
rect 24578 43840 24584 43852
rect 24075 43812 24584 43840
rect 24075 43809 24087 43812
rect 24029 43803 24087 43809
rect 24578 43800 24584 43812
rect 24636 43800 24642 43852
rect 25056 43849 25084 43880
rect 26694 43868 26700 43880
rect 26752 43868 26758 43920
rect 29362 43908 29368 43920
rect 28276 43880 29368 43908
rect 25041 43843 25099 43849
rect 25041 43809 25053 43843
rect 25087 43809 25099 43843
rect 25866 43840 25872 43852
rect 25827 43812 25872 43840
rect 25041 43803 25099 43809
rect 25866 43800 25872 43812
rect 25924 43800 25930 43852
rect 26602 43840 26608 43852
rect 26563 43812 26608 43840
rect 26602 43800 26608 43812
rect 26660 43800 26666 43852
rect 27522 43840 27528 43852
rect 27483 43812 27528 43840
rect 27522 43800 27528 43812
rect 27580 43800 27586 43852
rect 25504 43784 25556 43790
rect 23477 43775 23535 43781
rect 23477 43741 23489 43775
rect 23523 43741 23535 43775
rect 23477 43735 23535 43741
rect 23661 43775 23719 43781
rect 23661 43741 23673 43775
rect 23707 43772 23719 43775
rect 24762 43772 24768 43784
rect 23707 43744 24768 43772
rect 23707 43741 23719 43744
rect 23661 43735 23719 43741
rect 20714 43704 20720 43716
rect 20675 43676 20720 43704
rect 20714 43664 20720 43676
rect 20772 43664 20778 43716
rect 23492 43704 23520 43735
rect 24762 43732 24768 43744
rect 24820 43732 24826 43784
rect 26881 43775 26939 43781
rect 26881 43741 26893 43775
rect 26927 43772 26939 43775
rect 27246 43772 27252 43784
rect 26927 43744 27252 43772
rect 26927 43741 26939 43744
rect 26881 43735 26939 43741
rect 27246 43732 27252 43744
rect 27304 43732 27310 43784
rect 28276 43781 28304 43880
rect 29362 43868 29368 43880
rect 29420 43868 29426 43920
rect 34698 43868 34704 43920
rect 34756 43908 34762 43920
rect 37369 43911 37427 43917
rect 37369 43908 37381 43911
rect 34756 43880 37381 43908
rect 34756 43868 34762 43880
rect 37369 43877 37381 43880
rect 37415 43877 37427 43911
rect 38010 43908 38016 43920
rect 37971 43880 38016 43908
rect 37369 43871 37427 43877
rect 38010 43868 38016 43880
rect 38068 43868 38074 43920
rect 29086 43800 29092 43852
rect 29144 43840 29150 43852
rect 30009 43843 30067 43849
rect 30009 43840 30021 43843
rect 29144 43812 30021 43840
rect 29144 43800 29150 43812
rect 30009 43809 30021 43812
rect 30055 43809 30067 43843
rect 30009 43803 30067 43809
rect 33226 43800 33232 43852
rect 33284 43840 33290 43852
rect 34333 43843 34391 43849
rect 34333 43840 34345 43843
rect 33284 43812 34345 43840
rect 33284 43800 33290 43812
rect 34333 43809 34345 43812
rect 34379 43840 34391 43843
rect 36630 43840 36636 43852
rect 34379 43812 36636 43840
rect 34379 43809 34391 43812
rect 34333 43803 34391 43809
rect 36630 43800 36636 43812
rect 36688 43800 36694 43852
rect 28261 43775 28319 43781
rect 28261 43741 28273 43775
rect 28307 43741 28319 43775
rect 28534 43772 28540 43784
rect 28495 43744 28540 43772
rect 28261 43735 28319 43741
rect 28534 43732 28540 43744
rect 28592 43732 28598 43784
rect 29730 43732 29736 43784
rect 29788 43772 29794 43784
rect 30193 43775 30251 43781
rect 30193 43772 30205 43775
rect 29788 43744 30205 43772
rect 29788 43732 29794 43744
rect 30193 43741 30205 43744
rect 30239 43741 30251 43775
rect 30193 43735 30251 43741
rect 30282 43732 30288 43784
rect 30340 43772 30346 43784
rect 31478 43772 31484 43784
rect 30340 43744 31484 43772
rect 30340 43732 30346 43744
rect 31478 43732 31484 43744
rect 31536 43732 31542 43784
rect 32490 43732 32496 43784
rect 32548 43772 32554 43784
rect 32585 43775 32643 43781
rect 32585 43772 32597 43775
rect 32548 43744 32597 43772
rect 32548 43732 32554 43744
rect 32585 43741 32597 43744
rect 32631 43741 32643 43775
rect 32585 43735 32643 43741
rect 33134 43732 33140 43784
rect 33192 43772 33198 43784
rect 33413 43775 33471 43781
rect 33413 43772 33425 43775
rect 33192 43744 33425 43772
rect 33192 43732 33198 43744
rect 33413 43741 33425 43744
rect 33459 43741 33471 43775
rect 33413 43735 33471 43741
rect 33597 43775 33655 43781
rect 33597 43741 33609 43775
rect 33643 43772 33655 43775
rect 33962 43772 33968 43784
rect 33643 43744 33968 43772
rect 33643 43741 33655 43744
rect 33597 43735 33655 43741
rect 33962 43732 33968 43744
rect 34020 43732 34026 43784
rect 35434 43772 35440 43784
rect 35395 43744 35440 43772
rect 35434 43732 35440 43744
rect 35492 43732 35498 43784
rect 35986 43732 35992 43784
rect 36044 43732 36050 43784
rect 25504 43726 25556 43732
rect 25314 43704 25320 43716
rect 23492 43676 25320 43704
rect 25314 43664 25320 43676
rect 25372 43664 25378 43716
rect 28166 43664 28172 43716
rect 28224 43704 28230 43716
rect 28445 43707 28503 43713
rect 28445 43704 28457 43707
rect 28224 43676 28457 43704
rect 28224 43664 28230 43676
rect 28445 43673 28457 43676
rect 28491 43673 28503 43707
rect 28445 43667 28503 43673
rect 32401 43707 32459 43713
rect 32401 43673 32413 43707
rect 32447 43704 32459 43707
rect 32674 43704 32680 43716
rect 32447 43676 32680 43704
rect 32447 43673 32459 43676
rect 32401 43667 32459 43673
rect 32674 43664 32680 43676
rect 32732 43664 32738 43716
rect 36004 43704 36032 43732
rect 36173 43707 36231 43713
rect 36173 43704 36185 43707
rect 36004 43676 36185 43704
rect 36173 43673 36185 43676
rect 36219 43673 36231 43707
rect 36173 43667 36231 43673
rect 36357 43707 36415 43713
rect 36357 43673 36369 43707
rect 36403 43704 36415 43707
rect 36538 43704 36544 43716
rect 36403 43676 36544 43704
rect 36403 43673 36415 43676
rect 36357 43667 36415 43673
rect 36538 43664 36544 43676
rect 36596 43704 36602 43716
rect 36906 43704 36912 43716
rect 36596 43676 36912 43704
rect 36596 43664 36602 43676
rect 36906 43664 36912 43676
rect 36964 43664 36970 43716
rect 20438 43596 20444 43648
rect 20496 43636 20502 43648
rect 21177 43639 21235 43645
rect 21177 43636 21189 43639
rect 20496 43608 21189 43636
rect 20496 43596 20502 43608
rect 21177 43605 21189 43608
rect 21223 43636 21235 43639
rect 21821 43639 21879 43645
rect 21821 43636 21833 43639
rect 21223 43608 21833 43636
rect 21223 43605 21235 43608
rect 21177 43599 21235 43605
rect 21821 43605 21833 43608
rect 21867 43636 21879 43639
rect 22462 43636 22468 43648
rect 21867 43608 22468 43636
rect 21867 43605 21879 43608
rect 21821 43599 21879 43605
rect 22462 43596 22468 43608
rect 22520 43636 22526 43648
rect 22830 43636 22836 43648
rect 22520 43608 22836 43636
rect 22520 43596 22526 43608
rect 22830 43596 22836 43608
rect 22888 43596 22894 43648
rect 1104 43546 48852 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 48852 43546
rect 1104 43472 48852 43494
rect 22830 43432 22836 43444
rect 22791 43404 22836 43432
rect 22830 43392 22836 43404
rect 22888 43392 22894 43444
rect 24578 43432 24584 43444
rect 24539 43404 24584 43432
rect 24578 43392 24584 43404
rect 24636 43392 24642 43444
rect 26145 43435 26203 43441
rect 26145 43401 26157 43435
rect 26191 43432 26203 43435
rect 26694 43432 26700 43444
rect 26191 43404 26700 43432
rect 26191 43401 26203 43404
rect 26145 43395 26203 43401
rect 24946 43364 24952 43376
rect 24780 43336 24952 43364
rect 24780 43305 24808 43336
rect 24946 43324 24952 43336
rect 25004 43364 25010 43376
rect 25498 43364 25504 43376
rect 25004 43336 25504 43364
rect 25004 43324 25010 43336
rect 25498 43324 25504 43336
rect 25556 43324 25562 43376
rect 24765 43299 24823 43305
rect 24765 43265 24777 43299
rect 24811 43265 24823 43299
rect 24765 43259 24823 43265
rect 25038 43256 25044 43308
rect 25096 43296 25102 43308
rect 25409 43299 25467 43305
rect 25409 43296 25421 43299
rect 25096 43268 25421 43296
rect 25096 43256 25102 43268
rect 25409 43265 25421 43268
rect 25455 43265 25467 43299
rect 25409 43259 25467 43265
rect 20714 43188 20720 43240
rect 20772 43228 20778 43240
rect 23477 43231 23535 43237
rect 23477 43228 23489 43231
rect 20772 43200 23489 43228
rect 20772 43188 20778 43200
rect 23477 43197 23489 43200
rect 23523 43228 23535 43231
rect 24118 43228 24124 43240
rect 23523 43200 24124 43228
rect 23523 43197 23535 43200
rect 23477 43191 23535 43197
rect 24118 43188 24124 43200
rect 24176 43228 24182 43240
rect 24854 43228 24860 43240
rect 24176 43200 24860 43228
rect 24176 43188 24182 43200
rect 24854 43188 24860 43200
rect 24912 43188 24918 43240
rect 24949 43231 25007 43237
rect 24949 43197 24961 43231
rect 24995 43228 25007 43231
rect 26160 43228 26188 43395
rect 26694 43392 26700 43404
rect 26752 43392 26758 43444
rect 27246 43432 27252 43444
rect 27207 43404 27252 43432
rect 27246 43392 27252 43404
rect 27304 43392 27310 43444
rect 27706 43392 27712 43444
rect 27764 43432 27770 43444
rect 28813 43435 28871 43441
rect 28813 43432 28825 43435
rect 27764 43404 28825 43432
rect 27764 43392 27770 43404
rect 28813 43401 28825 43404
rect 28859 43432 28871 43435
rect 28902 43432 28908 43444
rect 28859 43404 28908 43432
rect 28859 43401 28871 43404
rect 28813 43395 28871 43401
rect 28902 43392 28908 43404
rect 28960 43432 28966 43444
rect 29365 43435 29423 43441
rect 29365 43432 29377 43435
rect 28960 43404 29377 43432
rect 28960 43392 28966 43404
rect 29365 43401 29377 43404
rect 29411 43432 29423 43435
rect 29917 43435 29975 43441
rect 29917 43432 29929 43435
rect 29411 43404 29929 43432
rect 29411 43401 29423 43404
rect 29365 43395 29423 43401
rect 29917 43401 29929 43404
rect 29963 43432 29975 43435
rect 30282 43432 30288 43444
rect 29963 43404 30288 43432
rect 29963 43401 29975 43404
rect 29917 43395 29975 43401
rect 30282 43392 30288 43404
rect 30340 43392 30346 43444
rect 30374 43392 30380 43444
rect 30432 43432 30438 43444
rect 32309 43435 32367 43441
rect 32309 43432 32321 43435
rect 30432 43404 32321 43432
rect 30432 43392 30438 43404
rect 32309 43401 32321 43404
rect 32355 43401 32367 43435
rect 32309 43395 32367 43401
rect 32674 43392 32680 43444
rect 32732 43432 32738 43444
rect 32861 43435 32919 43441
rect 32861 43432 32873 43435
rect 32732 43404 32873 43432
rect 32732 43392 32738 43404
rect 32861 43401 32873 43404
rect 32907 43401 32919 43435
rect 32861 43395 32919 43401
rect 35437 43435 35495 43441
rect 35437 43401 35449 43435
rect 35483 43432 35495 43435
rect 35526 43432 35532 43444
rect 35483 43404 35532 43432
rect 35483 43401 35495 43404
rect 35437 43395 35495 43401
rect 35526 43392 35532 43404
rect 35584 43392 35590 43444
rect 36538 43432 36544 43444
rect 36499 43404 36544 43432
rect 36538 43392 36544 43404
rect 36596 43392 36602 43444
rect 37553 43435 37611 43441
rect 37553 43401 37565 43435
rect 37599 43432 37611 43435
rect 37642 43432 37648 43444
rect 37599 43404 37648 43432
rect 37599 43401 37611 43404
rect 37553 43395 37611 43401
rect 37642 43392 37648 43404
rect 37700 43392 37706 43444
rect 38010 43392 38016 43444
rect 38068 43432 38074 43444
rect 38565 43435 38623 43441
rect 38565 43432 38577 43435
rect 38068 43404 38577 43432
rect 38068 43392 38074 43404
rect 38565 43401 38577 43404
rect 38611 43401 38623 43435
rect 38565 43395 38623 43401
rect 38654 43392 38660 43444
rect 38712 43432 38718 43444
rect 39117 43435 39175 43441
rect 39117 43432 39129 43435
rect 38712 43404 39129 43432
rect 38712 43392 38718 43404
rect 39117 43401 39129 43404
rect 39163 43401 39175 43435
rect 39117 43395 39175 43401
rect 34514 43364 34520 43376
rect 34475 43336 34520 43364
rect 34514 43324 34520 43336
rect 34572 43324 34578 43376
rect 34701 43367 34759 43373
rect 34701 43333 34713 43367
rect 34747 43364 34759 43367
rect 35897 43367 35955 43373
rect 35897 43364 35909 43367
rect 34747 43336 35909 43364
rect 34747 43333 34759 43336
rect 34701 43327 34759 43333
rect 35897 43333 35909 43336
rect 35943 43364 35955 43367
rect 38105 43367 38163 43373
rect 38105 43364 38117 43367
rect 35943 43336 38117 43364
rect 35943 43333 35955 43336
rect 35897 43327 35955 43333
rect 38105 43333 38117 43336
rect 38151 43364 38163 43367
rect 39942 43364 39948 43376
rect 38151 43336 39948 43364
rect 38151 43333 38163 43336
rect 38105 43327 38163 43333
rect 39942 43324 39948 43336
rect 40000 43324 40006 43376
rect 27709 43299 27767 43305
rect 27709 43265 27721 43299
rect 27755 43296 27767 43299
rect 28074 43296 28080 43308
rect 27755 43268 28080 43296
rect 27755 43265 27767 43268
rect 27709 43259 27767 43265
rect 28074 43256 28080 43268
rect 28132 43256 28138 43308
rect 29914 43256 29920 43308
rect 29972 43296 29978 43308
rect 30466 43296 30472 43308
rect 29972 43268 30472 43296
rect 29972 43256 29978 43268
rect 30466 43256 30472 43268
rect 30524 43256 30530 43308
rect 31570 43296 31576 43308
rect 31531 43268 31576 43296
rect 31570 43256 31576 43268
rect 31628 43256 31634 43308
rect 33778 43296 33784 43308
rect 33739 43268 33784 43296
rect 33778 43256 33784 43268
rect 33836 43256 33842 43308
rect 34606 43256 34612 43308
rect 34664 43296 34670 43308
rect 34885 43299 34943 43305
rect 34885 43296 34897 43299
rect 34664 43268 34897 43296
rect 34664 43256 34670 43268
rect 34885 43265 34897 43268
rect 34931 43296 34943 43299
rect 35526 43296 35532 43308
rect 34931 43268 35532 43296
rect 34931 43265 34943 43268
rect 34885 43259 34943 43265
rect 35526 43256 35532 43268
rect 35584 43256 35590 43308
rect 24995 43200 26188 43228
rect 24995 43197 25007 43200
rect 24949 43191 25007 43197
rect 27890 43188 27896 43240
rect 27948 43228 27954 43240
rect 28169 43231 28227 43237
rect 28169 43228 28181 43231
rect 27948 43200 28181 43228
rect 27948 43188 27954 43200
rect 28169 43197 28181 43200
rect 28215 43197 28227 43231
rect 28169 43191 28227 43197
rect 24029 43095 24087 43101
rect 24029 43061 24041 43095
rect 24075 43092 24087 43095
rect 26234 43092 26240 43104
rect 24075 43064 26240 43092
rect 24075 43061 24087 43064
rect 24029 43055 24087 43061
rect 26234 43052 26240 43064
rect 26292 43052 26298 43104
rect 27430 43092 27436 43104
rect 27391 43064 27436 43092
rect 27430 43052 27436 43064
rect 27488 43052 27494 43104
rect 39666 43092 39672 43104
rect 39627 43064 39672 43092
rect 39666 43052 39672 43064
rect 39724 43052 39730 43104
rect 1104 43002 48852 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 48852 43002
rect 1104 42928 48852 42950
rect 24673 42891 24731 42897
rect 24673 42857 24685 42891
rect 24719 42888 24731 42891
rect 24762 42888 24768 42900
rect 24719 42860 24768 42888
rect 24719 42857 24731 42860
rect 24673 42851 24731 42857
rect 24762 42848 24768 42860
rect 24820 42848 24826 42900
rect 24854 42848 24860 42900
rect 24912 42888 24918 42900
rect 25590 42888 25596 42900
rect 24912 42860 25596 42888
rect 24912 42848 24918 42860
rect 25590 42848 25596 42860
rect 25648 42888 25654 42900
rect 25961 42891 26019 42897
rect 25961 42888 25973 42891
rect 25648 42860 25973 42888
rect 25648 42848 25654 42860
rect 25961 42857 25973 42860
rect 26007 42857 26019 42891
rect 25961 42851 26019 42857
rect 26234 42848 26240 42900
rect 26292 42888 26298 42900
rect 26605 42891 26663 42897
rect 26605 42888 26617 42891
rect 26292 42860 26617 42888
rect 26292 42848 26298 42860
rect 26605 42857 26617 42860
rect 26651 42888 26663 42891
rect 27706 42888 27712 42900
rect 26651 42860 27712 42888
rect 26651 42857 26663 42860
rect 26605 42851 26663 42857
rect 27706 42848 27712 42860
rect 27764 42848 27770 42900
rect 27893 42891 27951 42897
rect 27893 42857 27905 42891
rect 27939 42888 27951 42891
rect 29362 42888 29368 42900
rect 27939 42860 29368 42888
rect 27939 42857 27951 42860
rect 27893 42851 27951 42857
rect 29362 42848 29368 42860
rect 29420 42848 29426 42900
rect 29730 42888 29736 42900
rect 29691 42860 29736 42888
rect 29730 42848 29736 42860
rect 29788 42848 29794 42900
rect 30374 42888 30380 42900
rect 30335 42860 30380 42888
rect 30374 42848 30380 42860
rect 30432 42848 30438 42900
rect 30466 42848 30472 42900
rect 30524 42888 30530 42900
rect 31941 42891 31999 42897
rect 31941 42888 31953 42891
rect 30524 42860 31953 42888
rect 30524 42848 30530 42860
rect 31941 42857 31953 42860
rect 31987 42857 31999 42891
rect 31941 42851 31999 42857
rect 32585 42891 32643 42897
rect 32585 42857 32597 42891
rect 32631 42888 32643 42891
rect 32674 42888 32680 42900
rect 32631 42860 32680 42888
rect 32631 42857 32643 42860
rect 32585 42851 32643 42857
rect 32674 42848 32680 42860
rect 32732 42888 32738 42900
rect 33873 42891 33931 42897
rect 33873 42888 33885 42891
rect 32732 42860 33885 42888
rect 32732 42848 32738 42860
rect 33873 42857 33885 42860
rect 33919 42888 33931 42891
rect 34606 42888 34612 42900
rect 33919 42860 34612 42888
rect 33919 42857 33931 42860
rect 33873 42851 33931 42857
rect 34606 42848 34612 42860
rect 34664 42848 34670 42900
rect 36633 42891 36691 42897
rect 36633 42857 36645 42891
rect 36679 42888 36691 42891
rect 37642 42888 37648 42900
rect 36679 42860 37648 42888
rect 36679 42857 36691 42860
rect 36633 42851 36691 42857
rect 37642 42848 37648 42860
rect 37700 42848 37706 42900
rect 28902 42780 28908 42832
rect 28960 42820 28966 42832
rect 29089 42823 29147 42829
rect 29089 42820 29101 42823
rect 28960 42792 29101 42820
rect 28960 42780 28966 42792
rect 29089 42789 29101 42792
rect 29135 42789 29147 42823
rect 29089 42783 29147 42789
rect 23014 42752 23020 42764
rect 22975 42724 23020 42752
rect 23014 42712 23020 42724
rect 23072 42712 23078 42764
rect 24029 42755 24087 42761
rect 24029 42721 24041 42755
rect 24075 42752 24087 42755
rect 24210 42752 24216 42764
rect 24075 42724 24216 42752
rect 24075 42721 24087 42724
rect 24029 42715 24087 42721
rect 24210 42712 24216 42724
rect 24268 42712 24274 42764
rect 25130 42752 25136 42764
rect 24780 42724 25136 42752
rect 24780 42693 24808 42724
rect 25130 42712 25136 42724
rect 25188 42752 25194 42764
rect 25501 42755 25559 42761
rect 25501 42752 25513 42755
rect 25188 42724 25513 42752
rect 25188 42712 25194 42724
rect 25501 42721 25513 42724
rect 25547 42752 25559 42755
rect 26694 42752 26700 42764
rect 25547 42724 26700 42752
rect 25547 42721 25559 42724
rect 25501 42715 25559 42721
rect 26694 42712 26700 42724
rect 26752 42752 26758 42764
rect 27065 42755 27123 42761
rect 27065 42752 27077 42755
rect 26752 42724 27077 42752
rect 26752 42712 26758 42724
rect 27065 42721 27077 42724
rect 27111 42721 27123 42755
rect 28994 42752 29000 42764
rect 28907 42724 29000 42752
rect 27065 42715 27123 42721
rect 28966 42712 29000 42724
rect 29052 42752 29058 42764
rect 29748 42752 29776 42848
rect 30837 42755 30895 42761
rect 30837 42752 30849 42755
rect 29052 42724 30849 42752
rect 29052 42712 29058 42724
rect 30837 42721 30849 42724
rect 30883 42721 30895 42755
rect 30837 42715 30895 42721
rect 31294 42712 31300 42764
rect 31352 42752 31358 42764
rect 31389 42755 31447 42761
rect 31389 42752 31401 42755
rect 31352 42724 31401 42752
rect 31352 42712 31358 42724
rect 31389 42721 31401 42724
rect 31435 42752 31447 42755
rect 33045 42755 33103 42761
rect 33045 42752 33057 42755
rect 31435 42724 33057 42752
rect 31435 42721 31447 42724
rect 31389 42715 31447 42721
rect 33045 42721 33057 42724
rect 33091 42721 33103 42755
rect 33045 42715 33103 42721
rect 34330 42712 34336 42764
rect 34388 42752 34394 42764
rect 34885 42755 34943 42761
rect 34885 42752 34897 42755
rect 34388 42724 34897 42752
rect 34388 42712 34394 42724
rect 34885 42721 34897 42724
rect 34931 42752 34943 42755
rect 35437 42755 35495 42761
rect 35437 42752 35449 42755
rect 34931 42724 35449 42752
rect 34931 42721 34943 42724
rect 34885 42715 34943 42721
rect 35437 42721 35449 42724
rect 35483 42721 35495 42755
rect 35437 42715 35495 42721
rect 37185 42755 37243 42761
rect 37185 42721 37197 42755
rect 37231 42752 37243 42755
rect 38746 42752 38752 42764
rect 37231 42724 38752 42752
rect 37231 42721 37243 42724
rect 37185 42715 37243 42721
rect 38746 42712 38752 42724
rect 38804 42752 38810 42764
rect 39666 42752 39672 42764
rect 38804 42724 39672 42752
rect 38804 42712 38810 42724
rect 39666 42712 39672 42724
rect 39724 42712 39730 42764
rect 24765 42687 24823 42693
rect 24765 42653 24777 42687
rect 24811 42653 24823 42687
rect 24946 42684 24952 42696
rect 24907 42656 24952 42684
rect 24765 42647 24823 42653
rect 24946 42644 24952 42656
rect 25004 42644 25010 42696
rect 28537 42687 28595 42693
rect 28537 42653 28549 42687
rect 28583 42684 28595 42687
rect 28966 42684 28994 42712
rect 28583 42656 28994 42684
rect 28583 42653 28595 42656
rect 28537 42647 28595 42653
rect 36081 42619 36139 42625
rect 36081 42585 36093 42619
rect 36127 42616 36139 42619
rect 38010 42616 38016 42628
rect 36127 42588 38016 42616
rect 36127 42585 36139 42588
rect 36081 42579 36139 42585
rect 38010 42576 38016 42588
rect 38068 42576 38074 42628
rect 1104 42458 48852 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 48852 42458
rect 1104 42384 48852 42406
rect 24118 42344 24124 42356
rect 24079 42316 24124 42344
rect 24118 42304 24124 42316
rect 24176 42304 24182 42356
rect 25130 42344 25136 42356
rect 25091 42316 25136 42344
rect 25130 42304 25136 42316
rect 25188 42304 25194 42356
rect 25590 42344 25596 42356
rect 25551 42316 25596 42344
rect 25590 42304 25596 42316
rect 25648 42304 25654 42356
rect 26142 42304 26148 42356
rect 26200 42344 26206 42356
rect 26237 42347 26295 42353
rect 26237 42344 26249 42347
rect 26200 42316 26249 42344
rect 26200 42304 26206 42316
rect 26237 42313 26249 42316
rect 26283 42313 26295 42347
rect 26237 42307 26295 42313
rect 28629 42347 28687 42353
rect 28629 42313 28641 42347
rect 28675 42344 28687 42347
rect 28994 42344 29000 42356
rect 28675 42316 29000 42344
rect 28675 42313 28687 42316
rect 28629 42307 28687 42313
rect 28994 42304 29000 42316
rect 29052 42304 29058 42356
rect 29181 42347 29239 42353
rect 29181 42313 29193 42347
rect 29227 42344 29239 42347
rect 29362 42344 29368 42356
rect 29227 42316 29368 42344
rect 29227 42313 29239 42316
rect 29181 42307 29239 42313
rect 29362 42304 29368 42316
rect 29420 42304 29426 42356
rect 29638 42304 29644 42356
rect 29696 42344 29702 42356
rect 29733 42347 29791 42353
rect 29733 42344 29745 42347
rect 29696 42316 29745 42344
rect 29696 42304 29702 42316
rect 29733 42313 29745 42316
rect 29779 42344 29791 42347
rect 30006 42344 30012 42356
rect 29779 42316 30012 42344
rect 29779 42313 29791 42316
rect 29733 42307 29791 42313
rect 30006 42304 30012 42316
rect 30064 42344 30070 42356
rect 30929 42347 30987 42353
rect 30929 42344 30941 42347
rect 30064 42316 30941 42344
rect 30064 42304 30070 42316
rect 30929 42313 30941 42316
rect 30975 42313 30987 42347
rect 30929 42307 30987 42313
rect 32401 42347 32459 42353
rect 32401 42313 32413 42347
rect 32447 42344 32459 42347
rect 33226 42344 33232 42356
rect 32447 42316 33232 42344
rect 32447 42313 32459 42316
rect 32401 42307 32459 42313
rect 33226 42304 33232 42316
rect 33284 42304 33290 42356
rect 33597 42347 33655 42353
rect 33597 42313 33609 42347
rect 33643 42344 33655 42347
rect 34517 42347 34575 42353
rect 34517 42344 34529 42347
rect 33643 42316 34529 42344
rect 33643 42313 33655 42316
rect 33597 42307 33655 42313
rect 34517 42313 34529 42316
rect 34563 42344 34575 42347
rect 34698 42344 34704 42356
rect 34563 42316 34704 42344
rect 34563 42313 34575 42316
rect 34517 42307 34575 42313
rect 34698 42304 34704 42316
rect 34756 42344 34762 42356
rect 35713 42347 35771 42353
rect 35713 42344 35725 42347
rect 34756 42316 35725 42344
rect 34756 42304 34762 42316
rect 35713 42313 35725 42316
rect 35759 42313 35771 42347
rect 35713 42307 35771 42313
rect 36357 42347 36415 42353
rect 36357 42313 36369 42347
rect 36403 42344 36415 42347
rect 37458 42344 37464 42356
rect 36403 42316 37464 42344
rect 36403 42313 36415 42316
rect 36357 42307 36415 42313
rect 37458 42304 37464 42316
rect 37516 42304 37522 42356
rect 27249 42279 27307 42285
rect 27249 42245 27261 42279
rect 27295 42276 27307 42279
rect 30374 42276 30380 42288
rect 27295 42248 30380 42276
rect 27295 42245 27307 42248
rect 27249 42239 27307 42245
rect 30374 42236 30380 42248
rect 30432 42236 30438 42288
rect 30466 42236 30472 42288
rect 30524 42276 30530 42288
rect 31481 42279 31539 42285
rect 31481 42276 31493 42279
rect 30524 42248 31493 42276
rect 30524 42236 30530 42248
rect 31481 42245 31493 42248
rect 31527 42245 31539 42279
rect 31481 42239 31539 42245
rect 33045 42279 33103 42285
rect 33045 42245 33057 42279
rect 33091 42276 33103 42279
rect 34330 42276 34336 42288
rect 33091 42248 34336 42276
rect 33091 42245 33103 42248
rect 33045 42239 33103 42245
rect 34330 42236 34336 42248
rect 34388 42276 34394 42288
rect 34977 42279 35035 42285
rect 34977 42276 34989 42279
rect 34388 42248 34989 42276
rect 34388 42236 34394 42248
rect 34977 42245 34989 42248
rect 35023 42245 35035 42279
rect 34977 42239 35035 42245
rect 27706 42004 27712 42016
rect 27667 41976 27712 42004
rect 27706 41964 27712 41976
rect 27764 42004 27770 42016
rect 30466 42004 30472 42016
rect 27764 41976 30472 42004
rect 27764 41964 27770 41976
rect 30466 41964 30472 41976
rect 30524 41964 30530 42016
rect 1104 41914 48852 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 48852 41914
rect 1104 41840 48852 41862
rect 24210 41760 24216 41812
rect 24268 41800 24274 41812
rect 25317 41803 25375 41809
rect 25317 41800 25329 41803
rect 24268 41772 25329 41800
rect 24268 41760 24274 41772
rect 25317 41769 25329 41772
rect 25363 41769 25375 41803
rect 26234 41800 26240 41812
rect 26195 41772 26240 41800
rect 25317 41763 25375 41769
rect 26234 41760 26240 41772
rect 26292 41760 26298 41812
rect 26694 41760 26700 41812
rect 26752 41800 26758 41812
rect 27985 41803 28043 41809
rect 27985 41800 27997 41803
rect 26752 41772 27997 41800
rect 26752 41760 26758 41772
rect 27985 41769 27997 41772
rect 28031 41769 28043 41803
rect 29730 41800 29736 41812
rect 29691 41772 29736 41800
rect 27985 41763 28043 41769
rect 29730 41760 29736 41772
rect 29788 41800 29794 41812
rect 30837 41803 30895 41809
rect 30837 41800 30849 41803
rect 29788 41772 30849 41800
rect 29788 41760 29794 41772
rect 30837 41769 30849 41772
rect 30883 41769 30895 41803
rect 30837 41763 30895 41769
rect 26973 41735 27031 41741
rect 26973 41701 26985 41735
rect 27019 41732 27031 41735
rect 27706 41732 27712 41744
rect 27019 41704 27712 41732
rect 27019 41701 27031 41704
rect 26973 41695 27031 41701
rect 27706 41692 27712 41704
rect 27764 41732 27770 41744
rect 28629 41735 28687 41741
rect 28629 41732 28641 41735
rect 27764 41704 28641 41732
rect 27764 41692 27770 41704
rect 28629 41701 28641 41704
rect 28675 41701 28687 41735
rect 28629 41695 28687 41701
rect 29362 41692 29368 41744
rect 29420 41732 29426 41744
rect 30285 41735 30343 41741
rect 30285 41732 30297 41735
rect 29420 41704 30297 41732
rect 29420 41692 29426 41704
rect 30285 41701 30297 41704
rect 30331 41701 30343 41735
rect 30285 41695 30343 41701
rect 1104 41370 48852 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 48852 41370
rect 1104 41296 48852 41318
rect 28629 41259 28687 41265
rect 28629 41225 28641 41259
rect 28675 41256 28687 41259
rect 29638 41256 29644 41268
rect 28675 41228 29644 41256
rect 28675 41225 28687 41228
rect 28629 41219 28687 41225
rect 29638 41216 29644 41228
rect 29696 41216 29702 41268
rect 1104 40826 48852 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 48852 40826
rect 1104 40752 48852 40774
rect 1104 40282 48852 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 48852 40282
rect 1104 40208 48852 40230
rect 1104 39738 48852 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 48852 39738
rect 1104 39664 48852 39686
rect 1104 39194 48852 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 48852 39194
rect 1104 39120 48852 39142
rect 1104 38650 48852 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 48852 38650
rect 1104 38576 48852 38598
rect 1104 38106 48852 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 48852 38106
rect 1104 38032 48852 38054
rect 1104 37562 48852 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 48852 37562
rect 1104 37488 48852 37510
rect 1104 37018 48852 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 48852 37018
rect 1104 36944 48852 36966
rect 1104 36474 48852 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 48852 36474
rect 1104 36400 48852 36422
rect 1104 35930 48852 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 48852 35930
rect 1104 35856 48852 35878
rect 1104 35386 48852 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 48852 35386
rect 1104 35312 48852 35334
rect 1104 34842 48852 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 48852 34842
rect 1104 34768 48852 34790
rect 1104 34298 48852 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 48852 34298
rect 1104 34224 48852 34246
rect 1104 33754 48852 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 48852 33754
rect 1104 33680 48852 33702
rect 1104 33210 48852 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 48852 33210
rect 1104 33136 48852 33158
rect 1104 32666 48852 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 48852 32666
rect 1104 32592 48852 32614
rect 1104 32122 48852 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 48852 32122
rect 1104 32048 48852 32070
rect 1104 31578 48852 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 48852 31578
rect 1104 31504 48852 31526
rect 1104 31034 48852 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 48852 31034
rect 1104 30960 48852 30982
rect 1104 30490 48852 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 48852 30490
rect 1104 30416 48852 30438
rect 1104 29946 48852 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 48852 29946
rect 1104 29872 48852 29894
rect 1104 29402 48852 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 48852 29402
rect 1104 29328 48852 29350
rect 1104 28858 48852 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 48852 28858
rect 1104 28784 48852 28806
rect 1104 28314 48852 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 48852 28314
rect 1104 28240 48852 28262
rect 1104 27770 48852 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 48852 27770
rect 1104 27696 48852 27718
rect 1104 27226 48852 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 48852 27226
rect 1104 27152 48852 27174
rect 1104 26682 48852 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 48852 26682
rect 1104 26608 48852 26630
rect 1104 26138 48852 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 48852 26138
rect 1104 26064 48852 26086
rect 1104 25594 48852 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 48852 25594
rect 1104 25520 48852 25542
rect 1104 25050 48852 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 48852 25050
rect 1104 24976 48852 24998
rect 1104 24506 48852 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 48852 24506
rect 1104 24432 48852 24454
rect 1104 23962 48852 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 48852 23962
rect 1104 23888 48852 23910
rect 1104 23418 48852 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 48852 23418
rect 1104 23344 48852 23366
rect 1104 22874 48852 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 48852 22874
rect 1104 22800 48852 22822
rect 1104 22330 48852 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 48852 22330
rect 1104 22256 48852 22278
rect 1104 21786 48852 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 48852 21786
rect 1104 21712 48852 21734
rect 1104 21242 48852 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 48852 21242
rect 1104 21168 48852 21190
rect 1104 20698 48852 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 48852 20698
rect 1104 20624 48852 20646
rect 1104 20154 48852 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 48852 20154
rect 1104 20080 48852 20102
rect 1104 19610 48852 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 48852 19610
rect 1104 19536 48852 19558
rect 1104 19066 48852 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 48852 19066
rect 1104 18992 48852 19014
rect 1104 18522 48852 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 48852 18522
rect 1104 18448 48852 18470
rect 1104 17978 48852 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 48852 17978
rect 1104 17904 48852 17926
rect 1104 17434 48852 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 48852 17434
rect 1104 17360 48852 17382
rect 1104 16890 48852 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 48852 16890
rect 1104 16816 48852 16838
rect 1104 16346 48852 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 48852 16346
rect 1104 16272 48852 16294
rect 1104 15802 48852 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 48852 15802
rect 1104 15728 48852 15750
rect 1104 15258 48852 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 48852 15258
rect 1104 15184 48852 15206
rect 1104 14714 48852 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 48852 14714
rect 1104 14640 48852 14662
rect 1104 14170 48852 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 48852 14170
rect 1104 14096 48852 14118
rect 1104 13626 48852 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 48852 13626
rect 1104 13552 48852 13574
rect 1104 13082 48852 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 48852 13082
rect 1104 13008 48852 13030
rect 1104 12538 48852 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 48852 12538
rect 1104 12464 48852 12486
rect 1104 11994 48852 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 48852 11994
rect 1104 11920 48852 11942
rect 1104 11450 48852 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 48852 11450
rect 1104 11376 48852 11398
rect 1104 10906 48852 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 48852 10906
rect 1104 10832 48852 10854
rect 1104 10362 48852 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 48852 10362
rect 1104 10288 48852 10310
rect 1104 9818 48852 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 48852 9818
rect 1104 9744 48852 9766
rect 1104 9274 48852 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 48852 9274
rect 1104 9200 48852 9222
rect 1104 8730 48852 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 48852 8730
rect 1104 8656 48852 8678
rect 1104 8186 48852 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 48852 8186
rect 1104 8112 48852 8134
rect 1104 7642 48852 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 48852 7642
rect 1104 7568 48852 7590
rect 1104 7098 48852 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 48852 7098
rect 1104 7024 48852 7046
rect 22922 6780 22928 6792
rect 22883 6752 22928 6780
rect 22922 6740 22928 6752
rect 22980 6740 22986 6792
rect 25317 6783 25375 6789
rect 25317 6749 25329 6783
rect 25363 6749 25375 6783
rect 25317 6743 25375 6749
rect 20530 6672 20536 6724
rect 20588 6712 20594 6724
rect 25332 6712 25360 6743
rect 25777 6715 25835 6721
rect 25777 6712 25789 6715
rect 20588 6684 25789 6712
rect 20588 6672 20594 6684
rect 25777 6681 25789 6684
rect 25823 6712 25835 6715
rect 27154 6712 27160 6724
rect 25823 6684 27160 6712
rect 25823 6681 25835 6684
rect 25777 6675 25835 6681
rect 27154 6672 27160 6684
rect 27212 6672 27218 6724
rect 23017 6647 23075 6653
rect 23017 6613 23029 6647
rect 23063 6644 23075 6647
rect 23198 6644 23204 6656
rect 23063 6616 23204 6644
rect 23063 6613 23075 6616
rect 23017 6607 23075 6613
rect 23198 6604 23204 6616
rect 23256 6604 23262 6656
rect 24762 6604 24768 6656
rect 24820 6644 24826 6656
rect 25133 6647 25191 6653
rect 25133 6644 25145 6647
rect 24820 6616 25145 6644
rect 24820 6604 24826 6616
rect 25133 6613 25145 6616
rect 25179 6613 25191 6647
rect 25133 6607 25191 6613
rect 1104 6554 48852 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 48852 6554
rect 1104 6480 48852 6502
rect 20530 6440 20536 6452
rect 20491 6412 20536 6440
rect 20530 6400 20536 6412
rect 20588 6400 20594 6452
rect 27154 6440 27160 6452
rect 27115 6412 27160 6440
rect 27154 6400 27160 6412
rect 27212 6400 27218 6452
rect 23753 6375 23811 6381
rect 23753 6341 23765 6375
rect 23799 6372 23811 6375
rect 24489 6375 24547 6381
rect 24489 6372 24501 6375
rect 23799 6344 24501 6372
rect 23799 6341 23811 6344
rect 23753 6335 23811 6341
rect 24489 6341 24501 6344
rect 24535 6341 24547 6375
rect 24489 6335 24547 6341
rect 25038 6332 25044 6384
rect 25096 6372 25102 6384
rect 25961 6375 26019 6381
rect 25961 6372 25973 6375
rect 25096 6344 25973 6372
rect 25096 6332 25102 6344
rect 25961 6341 25973 6344
rect 26007 6341 26019 6375
rect 25961 6335 26019 6341
rect 21082 6264 21088 6316
rect 21140 6304 21146 6316
rect 22281 6307 22339 6313
rect 22281 6304 22293 6307
rect 21140 6276 22293 6304
rect 21140 6264 21146 6276
rect 22281 6273 22293 6276
rect 22327 6304 22339 6307
rect 22922 6304 22928 6316
rect 22327 6276 22928 6304
rect 22327 6273 22339 6276
rect 22281 6267 22339 6273
rect 22922 6264 22928 6276
rect 22980 6264 22986 6316
rect 23661 6307 23719 6313
rect 23661 6273 23673 6307
rect 23707 6273 23719 6307
rect 23661 6267 23719 6273
rect 23676 6168 23704 6267
rect 24026 6196 24032 6248
rect 24084 6236 24090 6248
rect 24397 6239 24455 6245
rect 24397 6236 24409 6239
rect 24084 6208 24409 6236
rect 24084 6196 24090 6208
rect 24397 6205 24409 6208
rect 24443 6205 24455 6239
rect 25866 6236 25872 6248
rect 25827 6208 25872 6236
rect 24397 6199 24455 6205
rect 25866 6196 25872 6208
rect 25924 6196 25930 6248
rect 26513 6239 26571 6245
rect 26513 6205 26525 6239
rect 26559 6236 26571 6239
rect 26602 6236 26608 6248
rect 26559 6208 26608 6236
rect 26559 6205 26571 6208
rect 26513 6199 26571 6205
rect 26602 6196 26608 6208
rect 26660 6196 26666 6248
rect 24762 6168 24768 6180
rect 23676 6140 24768 6168
rect 24762 6128 24768 6140
rect 24820 6128 24826 6180
rect 24946 6168 24952 6180
rect 24907 6140 24952 6168
rect 24946 6128 24952 6140
rect 25004 6128 25010 6180
rect 22373 6103 22431 6109
rect 22373 6069 22385 6103
rect 22419 6100 22431 6103
rect 22554 6100 22560 6112
rect 22419 6072 22560 6100
rect 22419 6069 22431 6072
rect 22373 6063 22431 6069
rect 22554 6060 22560 6072
rect 22612 6060 22618 6112
rect 23017 6103 23075 6109
rect 23017 6069 23029 6103
rect 23063 6100 23075 6103
rect 23106 6100 23112 6112
rect 23063 6072 23112 6100
rect 23063 6069 23075 6072
rect 23017 6063 23075 6069
rect 23106 6060 23112 6072
rect 23164 6060 23170 6112
rect 1104 6010 48852 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 48852 6010
rect 1104 5936 48852 5958
rect 19521 5899 19579 5905
rect 19521 5865 19533 5899
rect 19567 5896 19579 5899
rect 20530 5896 20536 5908
rect 19567 5868 20536 5896
rect 19567 5865 19579 5868
rect 19521 5859 19579 5865
rect 20530 5856 20536 5868
rect 20588 5856 20594 5908
rect 24026 5896 24032 5908
rect 23987 5868 24032 5896
rect 24026 5856 24032 5868
rect 24084 5856 24090 5908
rect 25038 5896 25044 5908
rect 24999 5868 25044 5896
rect 25038 5856 25044 5868
rect 25096 5856 25102 5908
rect 24762 5788 24768 5840
rect 24820 5828 24826 5840
rect 24820 5800 26832 5828
rect 24820 5788 24826 5800
rect 21913 5763 21971 5769
rect 21913 5729 21925 5763
rect 21959 5760 21971 5763
rect 22465 5763 22523 5769
rect 22465 5760 22477 5763
rect 21959 5732 22477 5760
rect 21959 5729 21971 5732
rect 21913 5723 21971 5729
rect 22465 5729 22477 5732
rect 22511 5729 22523 5763
rect 22922 5760 22928 5772
rect 22883 5732 22928 5760
rect 22465 5723 22523 5729
rect 22922 5720 22928 5732
rect 22980 5720 22986 5772
rect 20165 5695 20223 5701
rect 20165 5661 20177 5695
rect 20211 5692 20223 5695
rect 20254 5692 20260 5704
rect 20211 5664 20260 5692
rect 20211 5661 20223 5664
rect 20165 5655 20223 5661
rect 20254 5652 20260 5664
rect 20312 5652 20318 5704
rect 21082 5692 21088 5704
rect 21043 5664 21088 5692
rect 21082 5652 21088 5664
rect 21140 5652 21146 5704
rect 24964 5701 24992 5800
rect 25961 5763 26019 5769
rect 25961 5729 25973 5763
rect 26007 5760 26019 5763
rect 26234 5760 26240 5772
rect 26007 5732 26240 5760
rect 26007 5729 26019 5732
rect 25961 5723 26019 5729
rect 26234 5720 26240 5732
rect 26292 5720 26298 5772
rect 26804 5701 26832 5800
rect 24949 5695 25007 5701
rect 24949 5661 24961 5695
rect 24995 5661 25007 5695
rect 24949 5655 25007 5661
rect 26789 5695 26847 5701
rect 26789 5661 26801 5695
rect 26835 5661 26847 5695
rect 26789 5655 26847 5661
rect 27617 5695 27675 5701
rect 27617 5661 27629 5695
rect 27663 5692 27675 5695
rect 28077 5695 28135 5701
rect 28077 5692 28089 5695
rect 27663 5664 28089 5692
rect 27663 5661 27675 5664
rect 27617 5655 27675 5661
rect 28077 5661 28089 5664
rect 28123 5661 28135 5695
rect 28077 5655 28135 5661
rect 28905 5695 28963 5701
rect 28905 5661 28917 5695
rect 28951 5692 28963 5695
rect 28994 5692 29000 5704
rect 28951 5664 29000 5692
rect 28951 5661 28963 5664
rect 28905 5655 28963 5661
rect 22554 5624 22560 5636
rect 22515 5596 22560 5624
rect 22554 5584 22560 5596
rect 22612 5584 22618 5636
rect 26145 5627 26203 5633
rect 26145 5593 26157 5627
rect 26191 5593 26203 5627
rect 26145 5587 26203 5593
rect 21177 5559 21235 5565
rect 21177 5525 21189 5559
rect 21223 5556 21235 5559
rect 21726 5556 21732 5568
rect 21223 5528 21732 5556
rect 21223 5525 21235 5528
rect 21177 5519 21235 5525
rect 21726 5516 21732 5528
rect 21784 5516 21790 5568
rect 26160 5556 26188 5587
rect 26234 5584 26240 5636
rect 26292 5624 26298 5636
rect 26292 5596 26337 5624
rect 26292 5584 26298 5596
rect 26694 5584 26700 5636
rect 26752 5624 26758 5636
rect 27632 5624 27660 5655
rect 26752 5596 27660 5624
rect 28092 5624 28120 5655
rect 28994 5652 29000 5664
rect 29052 5652 29058 5704
rect 29086 5624 29092 5636
rect 28092 5596 29092 5624
rect 26752 5584 26758 5596
rect 29086 5584 29092 5596
rect 29144 5584 29150 5636
rect 26881 5559 26939 5565
rect 26881 5556 26893 5559
rect 26160 5528 26893 5556
rect 26881 5525 26893 5528
rect 26927 5525 26939 5559
rect 26881 5519 26939 5525
rect 27338 5516 27344 5568
rect 27396 5556 27402 5568
rect 27525 5559 27583 5565
rect 27525 5556 27537 5559
rect 27396 5528 27537 5556
rect 27396 5516 27402 5528
rect 27525 5525 27537 5528
rect 27571 5525 27583 5559
rect 27525 5519 27583 5525
rect 28169 5559 28227 5565
rect 28169 5525 28181 5559
rect 28215 5556 28227 5559
rect 28534 5556 28540 5568
rect 28215 5528 28540 5556
rect 28215 5525 28227 5528
rect 28169 5519 28227 5525
rect 28534 5516 28540 5528
rect 28592 5516 28598 5568
rect 1104 5466 48852 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 48852 5466
rect 1104 5392 48852 5414
rect 20806 5352 20812 5364
rect 20719 5324 20812 5352
rect 20806 5312 20812 5324
rect 20864 5352 20870 5364
rect 21082 5352 21088 5364
rect 20864 5324 21088 5352
rect 20864 5312 20870 5324
rect 21082 5312 21088 5324
rect 21140 5312 21146 5364
rect 23106 5284 23112 5296
rect 23067 5256 23112 5284
rect 23106 5244 23112 5256
rect 23164 5244 23170 5296
rect 24578 5284 24584 5296
rect 24539 5256 24584 5284
rect 24578 5244 24584 5256
rect 24636 5244 24642 5296
rect 27338 5284 27344 5296
rect 27299 5256 27344 5284
rect 27338 5244 27344 5256
rect 27396 5244 27402 5296
rect 28534 5284 28540 5296
rect 28495 5256 28540 5284
rect 28534 5244 28540 5256
rect 28592 5244 28598 5296
rect 29086 5244 29092 5296
rect 29144 5244 29150 5296
rect 19981 5219 20039 5225
rect 19981 5185 19993 5219
rect 20027 5216 20039 5219
rect 20530 5216 20536 5228
rect 20027 5188 20536 5216
rect 20027 5185 20039 5188
rect 19981 5179 20039 5185
rect 20530 5176 20536 5188
rect 20588 5216 20594 5228
rect 20625 5219 20683 5225
rect 20625 5216 20637 5219
rect 20588 5188 20637 5216
rect 20588 5176 20594 5188
rect 20625 5185 20637 5188
rect 20671 5185 20683 5219
rect 20625 5179 20683 5185
rect 25777 5219 25835 5225
rect 25777 5185 25789 5219
rect 25823 5216 25835 5219
rect 25866 5216 25872 5228
rect 25823 5188 25872 5216
rect 25823 5185 25835 5188
rect 25777 5179 25835 5185
rect 25866 5176 25872 5188
rect 25924 5176 25930 5228
rect 26234 5176 26240 5228
rect 26292 5216 26298 5228
rect 26421 5219 26479 5225
rect 26421 5216 26433 5219
rect 26292 5188 26433 5216
rect 26292 5176 26298 5188
rect 26421 5185 26433 5188
rect 26467 5185 26479 5219
rect 29104 5216 29132 5244
rect 29733 5219 29791 5225
rect 29733 5216 29745 5219
rect 29104 5188 29745 5216
rect 26421 5179 26479 5185
rect 29733 5185 29745 5188
rect 29779 5216 29791 5219
rect 29822 5216 29828 5228
rect 29779 5188 29828 5216
rect 29779 5185 29791 5188
rect 29733 5179 29791 5185
rect 29822 5176 29828 5188
rect 29880 5176 29886 5228
rect 21453 5151 21511 5157
rect 21453 5117 21465 5151
rect 21499 5148 21511 5151
rect 23017 5151 23075 5157
rect 23017 5148 23029 5151
rect 21499 5120 23029 5148
rect 21499 5117 21511 5120
rect 21453 5111 21511 5117
rect 23017 5117 23029 5120
rect 23063 5117 23075 5151
rect 24489 5151 24547 5157
rect 24489 5148 24501 5151
rect 23017 5111 23075 5117
rect 23492 5120 24501 5148
rect 22465 5083 22523 5089
rect 22465 5049 22477 5083
rect 22511 5080 22523 5083
rect 23492 5080 23520 5120
rect 24489 5117 24501 5120
rect 24535 5117 24547 5151
rect 24489 5111 24547 5117
rect 25133 5151 25191 5157
rect 25133 5117 25145 5151
rect 25179 5148 25191 5151
rect 25222 5148 25228 5160
rect 25179 5120 25228 5148
rect 25179 5117 25191 5120
rect 25133 5111 25191 5117
rect 25222 5108 25228 5120
rect 25280 5108 25286 5160
rect 27249 5151 27307 5157
rect 27249 5117 27261 5151
rect 27295 5148 27307 5151
rect 27338 5148 27344 5160
rect 27295 5120 27344 5148
rect 27295 5117 27307 5120
rect 27249 5111 27307 5117
rect 27338 5108 27344 5120
rect 27396 5108 27402 5160
rect 28442 5148 28448 5160
rect 28403 5120 28448 5148
rect 28442 5108 28448 5120
rect 28500 5108 28506 5160
rect 29089 5151 29147 5157
rect 29089 5117 29101 5151
rect 29135 5148 29147 5151
rect 29178 5148 29184 5160
rect 29135 5120 29184 5148
rect 29135 5117 29147 5120
rect 29089 5111 29147 5117
rect 29178 5108 29184 5120
rect 29236 5108 29242 5160
rect 22511 5052 23520 5080
rect 23569 5083 23627 5089
rect 22511 5049 22523 5052
rect 22465 5043 22523 5049
rect 23569 5049 23581 5083
rect 23615 5049 23627 5083
rect 27798 5080 27804 5092
rect 27759 5052 27804 5080
rect 23569 5043 23627 5049
rect 19426 5012 19432 5024
rect 19387 4984 19432 5012
rect 19426 4972 19432 4984
rect 19484 4972 19490 5024
rect 20073 5015 20131 5021
rect 20073 4981 20085 5015
rect 20119 5012 20131 5015
rect 20346 5012 20352 5024
rect 20119 4984 20352 5012
rect 20119 4981 20131 4984
rect 20073 4975 20131 4981
rect 20346 4972 20352 4984
rect 20404 4972 20410 5024
rect 23474 4972 23480 5024
rect 23532 5012 23538 5024
rect 23584 5012 23612 5043
rect 27798 5040 27804 5052
rect 27856 5040 27862 5092
rect 23532 4984 23612 5012
rect 23532 4972 23538 4984
rect 29086 4972 29092 5024
rect 29144 5012 29150 5024
rect 29641 5015 29699 5021
rect 29641 5012 29653 5015
rect 29144 4984 29653 5012
rect 29144 4972 29150 4984
rect 29641 4981 29653 4984
rect 29687 4981 29699 5015
rect 29641 4975 29699 4981
rect 1104 4922 48852 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 48852 4922
rect 1104 4848 48852 4870
rect 27338 4808 27344 4820
rect 27299 4780 27344 4808
rect 27338 4768 27344 4780
rect 27396 4768 27402 4820
rect 19705 4743 19763 4749
rect 19705 4709 19717 4743
rect 19751 4740 19763 4743
rect 22186 4740 22192 4752
rect 19751 4712 21680 4740
rect 22147 4712 22192 4740
rect 19751 4709 19763 4712
rect 19705 4703 19763 4709
rect 20254 4672 20260 4684
rect 20215 4644 20260 4672
rect 20254 4632 20260 4644
rect 20312 4632 20318 4684
rect 21652 4681 21680 4712
rect 22186 4700 22192 4712
rect 22244 4700 22250 4752
rect 21637 4675 21695 4681
rect 21637 4641 21649 4675
rect 21683 4641 21695 4675
rect 23566 4672 23572 4684
rect 23527 4644 23572 4672
rect 21637 4635 21695 4641
rect 23566 4632 23572 4644
rect 23624 4632 23630 4684
rect 25041 4675 25099 4681
rect 25041 4641 25053 4675
rect 25087 4672 25099 4675
rect 25593 4675 25651 4681
rect 25593 4672 25605 4675
rect 25087 4644 25605 4672
rect 25087 4641 25099 4644
rect 25041 4635 25099 4641
rect 25593 4641 25605 4644
rect 25639 4641 25651 4675
rect 26050 4672 26056 4684
rect 26011 4644 26056 4672
rect 25593 4635 25651 4641
rect 26050 4632 26056 4644
rect 26108 4632 26114 4684
rect 28810 4672 28816 4684
rect 28771 4644 28816 4672
rect 28810 4632 28816 4644
rect 28868 4632 28874 4684
rect 28994 4632 29000 4684
rect 29052 4672 29058 4684
rect 29089 4675 29147 4681
rect 29089 4672 29101 4675
rect 29052 4644 29101 4672
rect 29052 4632 29058 4644
rect 29089 4641 29101 4644
rect 29135 4641 29147 4675
rect 29089 4635 29147 4641
rect 16942 4604 16948 4616
rect 16903 4576 16948 4604
rect 16942 4564 16948 4576
rect 17000 4564 17006 4616
rect 18877 4607 18935 4613
rect 18877 4573 18889 4607
rect 18923 4604 18935 4607
rect 19978 4604 19984 4616
rect 18923 4576 19984 4604
rect 18923 4573 18935 4576
rect 18877 4567 18935 4573
rect 19978 4564 19984 4576
rect 20036 4564 20042 4616
rect 26881 4607 26939 4613
rect 26881 4573 26893 4607
rect 26927 4604 26939 4607
rect 27154 4604 27160 4616
rect 26927 4576 27160 4604
rect 26927 4573 26939 4576
rect 26881 4567 26939 4573
rect 27154 4564 27160 4576
rect 27212 4564 27218 4616
rect 20346 4536 20352 4548
rect 20307 4508 20352 4536
rect 20346 4496 20352 4508
rect 20404 4496 20410 4548
rect 20901 4539 20959 4545
rect 20901 4505 20913 4539
rect 20947 4536 20959 4539
rect 21082 4536 21088 4548
rect 20947 4508 21088 4536
rect 20947 4505 20959 4508
rect 20901 4499 20959 4505
rect 21082 4496 21088 4508
rect 21140 4496 21146 4548
rect 21726 4496 21732 4548
rect 21784 4536 21790 4548
rect 21784 4508 21829 4536
rect 21784 4496 21790 4508
rect 21910 4496 21916 4548
rect 21968 4536 21974 4548
rect 23109 4539 23167 4545
rect 21968 4508 22094 4536
rect 21968 4496 21974 4508
rect 22066 4468 22094 4508
rect 23109 4505 23121 4539
rect 23155 4505 23167 4539
rect 23109 4499 23167 4505
rect 23124 4468 23152 4499
rect 23198 4496 23204 4548
rect 23256 4536 23262 4548
rect 25682 4536 25688 4548
rect 23256 4508 23301 4536
rect 25643 4508 25688 4536
rect 23256 4496 23262 4508
rect 25682 4496 25688 4508
rect 25740 4496 25746 4548
rect 28994 4536 29000 4548
rect 28955 4508 29000 4536
rect 28994 4496 29000 4508
rect 29052 4496 29058 4548
rect 26694 4468 26700 4480
rect 22066 4440 23152 4468
rect 26655 4440 26700 4468
rect 26694 4428 26700 4440
rect 26752 4428 26758 4480
rect 1104 4378 48852 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 48852 4378
rect 1104 4304 48852 4326
rect 23569 4267 23627 4273
rect 23569 4233 23581 4267
rect 23615 4264 23627 4267
rect 24578 4264 24584 4276
rect 23615 4236 24584 4264
rect 23615 4233 23627 4236
rect 23569 4227 23627 4233
rect 24578 4224 24584 4236
rect 24636 4224 24642 4276
rect 25593 4267 25651 4273
rect 25593 4233 25605 4267
rect 25639 4264 25651 4267
rect 25682 4264 25688 4276
rect 25639 4236 25688 4264
rect 25639 4233 25651 4236
rect 25593 4227 25651 4233
rect 25682 4224 25688 4236
rect 25740 4224 25746 4276
rect 20806 4196 20812 4208
rect 19996 4168 20812 4196
rect 19996 4137 20024 4168
rect 20806 4156 20812 4168
rect 20864 4156 20870 4208
rect 22281 4199 22339 4205
rect 22281 4196 22293 4199
rect 21192 4168 22293 4196
rect 19981 4131 20039 4137
rect 19981 4097 19993 4131
rect 20027 4097 20039 4131
rect 19981 4091 20039 4097
rect 20073 4131 20131 4137
rect 20073 4097 20085 4131
rect 20119 4128 20131 4131
rect 21192 4128 21220 4168
rect 22281 4165 22293 4168
rect 22327 4165 22339 4199
rect 24302 4196 24308 4208
rect 24263 4168 24308 4196
rect 22281 4159 22339 4165
rect 24302 4156 24308 4168
rect 24360 4156 24366 4208
rect 27706 4196 27712 4208
rect 27667 4168 27712 4196
rect 27706 4156 27712 4168
rect 27764 4156 27770 4208
rect 28997 4199 29055 4205
rect 28997 4165 29009 4199
rect 29043 4196 29055 4199
rect 29733 4199 29791 4205
rect 29733 4196 29745 4199
rect 29043 4168 29745 4196
rect 29043 4165 29055 4168
rect 28997 4159 29055 4165
rect 29733 4165 29745 4168
rect 29779 4165 29791 4199
rect 29733 4159 29791 4165
rect 20119 4100 21220 4128
rect 23477 4131 23535 4137
rect 20119 4097 20131 4100
rect 20073 4091 20131 4097
rect 23477 4097 23489 4131
rect 23523 4128 23535 4131
rect 23658 4128 23664 4140
rect 23523 4100 23664 4128
rect 23523 4097 23535 4100
rect 23477 4091 23535 4097
rect 23658 4088 23664 4100
rect 23716 4088 23722 4140
rect 24854 4088 24860 4140
rect 24912 4128 24918 4140
rect 25501 4131 25559 4137
rect 25501 4128 25513 4131
rect 24912 4100 25513 4128
rect 24912 4088 24918 4100
rect 25501 4097 25513 4100
rect 25547 4097 25559 4131
rect 29822 4128 29828 4140
rect 29783 4100 29828 4128
rect 25501 4091 25559 4097
rect 29822 4088 29828 4100
rect 29880 4088 29886 4140
rect 19521 4063 19579 4069
rect 19521 4029 19533 4063
rect 19567 4060 19579 4063
rect 22189 4063 22247 4069
rect 22189 4060 22201 4063
rect 19567 4032 22201 4060
rect 19567 4029 19579 4032
rect 19521 4023 19579 4029
rect 22189 4029 22201 4032
rect 22235 4029 22247 4063
rect 22462 4060 22468 4072
rect 22423 4032 22468 4060
rect 22189 4023 22247 4029
rect 22462 4020 22468 4032
rect 22520 4020 22526 4072
rect 24213 4063 24271 4069
rect 24213 4029 24225 4063
rect 24259 4029 24271 4063
rect 24670 4060 24676 4072
rect 24631 4032 24676 4060
rect 24213 4023 24271 4029
rect 18233 3995 18291 4001
rect 18233 3961 18245 3995
rect 18279 3992 18291 3995
rect 19150 3992 19156 4004
rect 18279 3964 19156 3992
rect 18279 3961 18291 3964
rect 18233 3955 18291 3961
rect 19150 3952 19156 3964
rect 19208 3952 19214 4004
rect 21453 3995 21511 4001
rect 21453 3961 21465 3995
rect 21499 3992 21511 3995
rect 24228 3992 24256 4023
rect 24670 4020 24676 4032
rect 24728 4020 24734 4072
rect 27430 4060 27436 4072
rect 27391 4032 27436 4060
rect 27430 4020 27436 4032
rect 27488 4020 27494 4072
rect 27801 4063 27859 4069
rect 27801 4029 27813 4063
rect 27847 4060 27859 4063
rect 28902 4060 28908 4072
rect 27847 4032 28908 4060
rect 27847 4029 27859 4032
rect 27801 4023 27859 4029
rect 28902 4020 28908 4032
rect 28960 4020 28966 4072
rect 29089 4063 29147 4069
rect 29089 4029 29101 4063
rect 29135 4060 29147 4063
rect 29730 4060 29736 4072
rect 29135 4032 29736 4060
rect 29135 4029 29147 4032
rect 29089 4023 29147 4029
rect 29730 4020 29736 4032
rect 29788 4020 29794 4072
rect 21499 3964 24256 3992
rect 26605 3995 26663 4001
rect 21499 3961 21511 3964
rect 21453 3955 21511 3961
rect 26605 3961 26617 3995
rect 26651 3992 26663 3995
rect 28442 3992 28448 4004
rect 26651 3964 28448 3992
rect 26651 3961 26663 3964
rect 26605 3955 26663 3961
rect 28442 3952 28448 3964
rect 28500 3952 28506 4004
rect 28537 3995 28595 4001
rect 28537 3961 28549 3995
rect 28583 3992 28595 3995
rect 28583 3964 29132 3992
rect 28583 3961 28595 3964
rect 28537 3955 28595 3961
rect 29104 3936 29132 3964
rect 15010 3924 15016 3936
rect 14971 3896 15016 3924
rect 15010 3884 15016 3896
rect 15068 3884 15074 3936
rect 16114 3924 16120 3936
rect 16075 3896 16120 3924
rect 16114 3884 16120 3896
rect 16172 3884 16178 3936
rect 17589 3927 17647 3933
rect 17589 3893 17601 3927
rect 17635 3924 17647 3927
rect 18046 3924 18052 3936
rect 17635 3896 18052 3924
rect 17635 3893 17647 3896
rect 17589 3887 17647 3893
rect 18046 3884 18052 3896
rect 18104 3884 18110 3936
rect 18874 3924 18880 3936
rect 18835 3896 18880 3924
rect 18874 3884 18880 3896
rect 18932 3884 18938 3936
rect 20809 3927 20867 3933
rect 20809 3893 20821 3927
rect 20855 3924 20867 3927
rect 21910 3924 21916 3936
rect 20855 3896 21916 3924
rect 20855 3893 20867 3896
rect 20809 3887 20867 3893
rect 21910 3884 21916 3896
rect 21968 3884 21974 3936
rect 23658 3884 23664 3936
rect 23716 3924 23722 3936
rect 24762 3924 24768 3936
rect 23716 3896 24768 3924
rect 23716 3884 23722 3896
rect 24762 3884 24768 3896
rect 24820 3884 24826 3936
rect 29086 3884 29092 3936
rect 29144 3884 29150 3936
rect 29914 3884 29920 3936
rect 29972 3924 29978 3936
rect 30285 3927 30343 3933
rect 30285 3924 30297 3927
rect 29972 3896 30297 3924
rect 29972 3884 29978 3896
rect 30285 3893 30297 3896
rect 30331 3893 30343 3927
rect 30285 3887 30343 3893
rect 1104 3834 48852 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 48852 3834
rect 1104 3760 48852 3782
rect 18233 3723 18291 3729
rect 18233 3689 18245 3723
rect 18279 3720 18291 3723
rect 20806 3720 20812 3732
rect 18279 3692 20812 3720
rect 18279 3689 18291 3692
rect 18233 3683 18291 3689
rect 20806 3680 20812 3692
rect 20864 3680 20870 3732
rect 23293 3723 23351 3729
rect 23293 3689 23305 3723
rect 23339 3720 23351 3723
rect 25314 3720 25320 3732
rect 23339 3692 25320 3720
rect 23339 3689 23351 3692
rect 23293 3683 23351 3689
rect 25314 3680 25320 3692
rect 25372 3680 25378 3732
rect 26881 3723 26939 3729
rect 26881 3689 26893 3723
rect 26927 3720 26939 3723
rect 27706 3720 27712 3732
rect 26927 3692 27712 3720
rect 26927 3689 26939 3692
rect 26881 3683 26939 3689
rect 27706 3680 27712 3692
rect 27764 3680 27770 3732
rect 28902 3720 28908 3732
rect 28863 3692 28908 3720
rect 28902 3680 28908 3692
rect 28960 3680 28966 3732
rect 29730 3720 29736 3732
rect 29691 3692 29736 3720
rect 29730 3680 29736 3692
rect 29788 3680 29794 3732
rect 16301 3655 16359 3661
rect 16301 3621 16313 3655
rect 16347 3652 16359 3655
rect 17218 3652 17224 3664
rect 16347 3624 17224 3652
rect 16347 3621 16359 3624
rect 16301 3615 16359 3621
rect 17218 3612 17224 3624
rect 17276 3612 17282 3664
rect 17589 3655 17647 3661
rect 17589 3621 17601 3655
rect 17635 3652 17647 3655
rect 20254 3652 20260 3664
rect 17635 3624 20260 3652
rect 17635 3621 17647 3624
rect 17589 3615 17647 3621
rect 20254 3612 20260 3624
rect 20312 3612 20318 3664
rect 20625 3655 20683 3661
rect 20625 3621 20637 3655
rect 20671 3652 20683 3655
rect 24118 3652 24124 3664
rect 20671 3624 24124 3652
rect 20671 3621 20683 3624
rect 20625 3615 20683 3621
rect 24118 3612 24124 3624
rect 24176 3612 24182 3664
rect 24964 3624 25268 3652
rect 15013 3587 15071 3593
rect 15013 3553 15025 3587
rect 15059 3584 15071 3587
rect 15838 3584 15844 3596
rect 15059 3556 15844 3584
rect 15059 3553 15071 3556
rect 15013 3547 15071 3553
rect 15838 3544 15844 3556
rect 15896 3544 15902 3596
rect 16945 3587 17003 3593
rect 16945 3553 16957 3587
rect 16991 3584 17003 3587
rect 18598 3584 18604 3596
rect 16991 3556 18604 3584
rect 16991 3553 17003 3556
rect 16945 3547 17003 3553
rect 18598 3544 18604 3556
rect 18656 3544 18662 3596
rect 18874 3544 18880 3596
rect 18932 3584 18938 3596
rect 21177 3587 21235 3593
rect 21177 3584 21189 3587
rect 18932 3556 21189 3584
rect 18932 3544 18938 3556
rect 21177 3553 21189 3556
rect 21223 3553 21235 3587
rect 21177 3547 21235 3553
rect 21358 3544 21364 3596
rect 21416 3584 21422 3596
rect 21453 3587 21511 3593
rect 21453 3584 21465 3587
rect 21416 3556 21465 3584
rect 21416 3544 21422 3556
rect 21453 3553 21465 3556
rect 21499 3553 21511 3587
rect 21453 3547 21511 3553
rect 22741 3587 22799 3593
rect 22741 3553 22753 3587
rect 22787 3584 22799 3587
rect 24964 3584 24992 3624
rect 25240 3593 25268 3624
rect 27982 3612 27988 3664
rect 28040 3652 28046 3664
rect 29178 3652 29184 3664
rect 28040 3624 29184 3652
rect 28040 3612 28046 3624
rect 29178 3612 29184 3624
rect 29236 3612 29242 3664
rect 32950 3612 32956 3664
rect 33008 3652 33014 3664
rect 33597 3655 33655 3661
rect 33597 3652 33609 3655
rect 33008 3624 33609 3652
rect 33008 3612 33014 3624
rect 33597 3621 33609 3624
rect 33643 3621 33655 3655
rect 33597 3615 33655 3621
rect 36814 3612 36820 3664
rect 36872 3652 36878 3664
rect 37461 3655 37519 3661
rect 37461 3652 37473 3655
rect 36872 3624 37473 3652
rect 36872 3612 36878 3624
rect 37461 3621 37473 3624
rect 37507 3621 37519 3655
rect 37461 3615 37519 3621
rect 22787 3556 24992 3584
rect 25225 3587 25283 3593
rect 22787 3553 22799 3556
rect 22741 3547 22799 3553
rect 25225 3553 25237 3587
rect 25271 3553 25283 3587
rect 25498 3584 25504 3596
rect 25459 3556 25504 3584
rect 25225 3547 25283 3553
rect 25498 3544 25504 3556
rect 25556 3544 25562 3596
rect 28077 3587 28135 3593
rect 28077 3553 28089 3587
rect 28123 3584 28135 3587
rect 28258 3584 28264 3596
rect 28123 3556 28264 3584
rect 28123 3553 28135 3556
rect 28077 3547 28135 3553
rect 28258 3544 28264 3556
rect 28316 3544 28322 3596
rect 30190 3544 30196 3596
rect 30248 3584 30254 3596
rect 31021 3587 31079 3593
rect 31021 3584 31033 3587
rect 30248 3556 31033 3584
rect 30248 3544 30254 3556
rect 31021 3553 31033 3556
rect 31067 3553 31079 3587
rect 31021 3547 31079 3553
rect 34790 3544 34796 3596
rect 34848 3584 34854 3596
rect 35529 3587 35587 3593
rect 35529 3584 35541 3587
rect 34848 3556 35541 3584
rect 34848 3544 34854 3556
rect 35529 3553 35541 3556
rect 35575 3553 35587 3587
rect 35529 3547 35587 3553
rect 4154 3476 4160 3528
rect 4212 3516 4218 3528
rect 4249 3519 4307 3525
rect 4249 3516 4261 3519
rect 4212 3488 4261 3516
rect 4212 3476 4218 3488
rect 4249 3485 4261 3488
rect 4295 3485 4307 3519
rect 5166 3516 5172 3528
rect 5127 3488 5172 3516
rect 4249 3479 4307 3485
rect 5166 3476 5172 3488
rect 5224 3476 5230 3528
rect 5994 3516 6000 3528
rect 5955 3488 6000 3516
rect 5994 3476 6000 3488
rect 6052 3476 6058 3528
rect 6822 3516 6828 3528
rect 6783 3488 6828 3516
rect 6822 3476 6828 3488
rect 6880 3476 6886 3528
rect 7650 3516 7656 3528
rect 7611 3488 7656 3516
rect 7650 3476 7656 3488
rect 7708 3476 7714 3528
rect 8478 3516 8484 3528
rect 8439 3488 8484 3516
rect 8478 3476 8484 3488
rect 8536 3476 8542 3528
rect 9306 3516 9312 3528
rect 9267 3488 9312 3516
rect 9306 3476 9312 3488
rect 9364 3476 9370 3528
rect 10134 3516 10140 3528
rect 10095 3488 10140 3516
rect 10134 3476 10140 3488
rect 10192 3476 10198 3528
rect 10962 3516 10968 3528
rect 10923 3488 10968 3516
rect 10962 3476 10968 3488
rect 11020 3476 11026 3528
rect 11701 3519 11759 3525
rect 11701 3485 11713 3519
rect 11747 3516 11759 3519
rect 11790 3516 11796 3528
rect 11747 3488 11796 3516
rect 11747 3485 11759 3488
rect 11701 3479 11759 3485
rect 11790 3476 11796 3488
rect 11848 3476 11854 3528
rect 12345 3519 12403 3525
rect 12345 3485 12357 3519
rect 12391 3516 12403 3519
rect 12526 3516 12532 3528
rect 12391 3488 12532 3516
rect 12391 3485 12403 3488
rect 12345 3479 12403 3485
rect 12526 3476 12532 3488
rect 12584 3476 12590 3528
rect 12989 3519 13047 3525
rect 12989 3485 13001 3519
rect 13035 3516 13047 3519
rect 13078 3516 13084 3528
rect 13035 3488 13084 3516
rect 13035 3485 13047 3488
rect 12989 3479 13047 3485
rect 13078 3476 13084 3488
rect 13136 3476 13142 3528
rect 13630 3516 13636 3528
rect 13591 3488 13636 3516
rect 13630 3476 13636 3488
rect 13688 3476 13694 3528
rect 15657 3519 15715 3525
rect 15657 3485 15669 3519
rect 15703 3516 15715 3519
rect 16390 3516 16396 3528
rect 15703 3488 16396 3516
rect 15703 3485 15715 3488
rect 15657 3479 15715 3485
rect 16390 3476 16396 3488
rect 16448 3476 16454 3528
rect 18693 3519 18751 3525
rect 18693 3485 18705 3519
rect 18739 3516 18751 3519
rect 19242 3516 19248 3528
rect 18739 3488 19248 3516
rect 18739 3485 18751 3488
rect 18693 3479 18751 3485
rect 19242 3476 19248 3488
rect 19300 3516 19306 3528
rect 19797 3519 19855 3525
rect 19797 3516 19809 3519
rect 19300 3488 19809 3516
rect 19300 3476 19306 3488
rect 19797 3485 19809 3488
rect 19843 3516 19855 3519
rect 20714 3516 20720 3528
rect 19843 3488 20720 3516
rect 19843 3485 19855 3488
rect 19797 3479 19855 3485
rect 20714 3476 20720 3488
rect 20772 3476 20778 3528
rect 23201 3519 23259 3525
rect 23201 3485 23213 3519
rect 23247 3516 23259 3519
rect 23658 3516 23664 3528
rect 23247 3488 23664 3516
rect 23247 3485 23259 3488
rect 23201 3479 23259 3485
rect 23658 3476 23664 3488
rect 23716 3476 23722 3528
rect 24029 3519 24087 3525
rect 24029 3485 24041 3519
rect 24075 3485 24087 3519
rect 24029 3479 24087 3485
rect 18785 3451 18843 3457
rect 18785 3417 18797 3451
rect 18831 3448 18843 3451
rect 21269 3451 21327 3457
rect 21269 3448 21281 3451
rect 18831 3420 21281 3448
rect 18831 3417 18843 3420
rect 18785 3411 18843 3417
rect 21269 3417 21281 3420
rect 21315 3417 21327 3451
rect 24044 3448 24072 3479
rect 26694 3476 26700 3528
rect 26752 3516 26758 3528
rect 26789 3519 26847 3525
rect 26789 3516 26801 3519
rect 26752 3488 26801 3516
rect 26752 3476 26758 3488
rect 26789 3485 26801 3488
rect 26835 3485 26847 3519
rect 30282 3516 30288 3528
rect 26789 3479 26847 3485
rect 28828 3488 30288 3516
rect 24044 3420 25268 3448
rect 21269 3411 21327 3417
rect 19889 3383 19947 3389
rect 19889 3349 19901 3383
rect 19935 3380 19947 3383
rect 23014 3380 23020 3392
rect 19935 3352 23020 3380
rect 19935 3349 19947 3352
rect 19889 3343 19947 3349
rect 23014 3340 23020 3352
rect 23072 3340 23078 3392
rect 23937 3383 23995 3389
rect 23937 3349 23949 3383
rect 23983 3380 23995 3383
rect 25038 3380 25044 3392
rect 23983 3352 25044 3380
rect 23983 3349 23995 3352
rect 23937 3343 23995 3349
rect 25038 3340 25044 3352
rect 25096 3340 25102 3392
rect 25240 3380 25268 3420
rect 25314 3408 25320 3460
rect 25372 3457 25378 3460
rect 25372 3448 25384 3457
rect 25372 3420 25417 3448
rect 25372 3411 25384 3420
rect 25372 3408 25378 3411
rect 26804 3380 26832 3479
rect 28261 3451 28319 3457
rect 28261 3417 28273 3451
rect 28307 3417 28319 3451
rect 28261 3411 28319 3417
rect 25240 3352 26832 3380
rect 28276 3380 28304 3411
rect 28350 3408 28356 3460
rect 28408 3448 28414 3460
rect 28408 3420 28453 3448
rect 28408 3408 28414 3420
rect 28828 3380 28856 3488
rect 30282 3476 30288 3488
rect 30340 3476 30346 3528
rect 30561 3519 30619 3525
rect 30561 3485 30573 3519
rect 30607 3485 30619 3519
rect 30561 3479 30619 3485
rect 29822 3408 29828 3460
rect 29880 3448 29886 3460
rect 30576 3448 30604 3479
rect 31110 3476 31116 3528
rect 31168 3516 31174 3528
rect 31665 3519 31723 3525
rect 31665 3516 31677 3519
rect 31168 3488 31677 3516
rect 31168 3476 31174 3488
rect 31665 3485 31677 3488
rect 31711 3485 31723 3519
rect 31665 3479 31723 3485
rect 31846 3476 31852 3528
rect 31904 3516 31910 3528
rect 32309 3519 32367 3525
rect 32309 3516 32321 3519
rect 31904 3488 32321 3516
rect 31904 3476 31910 3488
rect 32309 3485 32321 3488
rect 32355 3485 32367 3519
rect 32309 3479 32367 3485
rect 32398 3476 32404 3528
rect 32456 3516 32462 3528
rect 32953 3519 33011 3525
rect 32953 3516 32965 3519
rect 32456 3488 32965 3516
rect 32456 3476 32462 3488
rect 32953 3485 32965 3488
rect 32999 3485 33011 3519
rect 32953 3479 33011 3485
rect 34330 3476 34336 3528
rect 34388 3516 34394 3528
rect 34885 3519 34943 3525
rect 34885 3516 34897 3519
rect 34388 3488 34897 3516
rect 34388 3476 34394 3488
rect 34885 3485 34897 3488
rect 34931 3485 34943 3519
rect 34885 3479 34943 3485
rect 35710 3476 35716 3528
rect 35768 3516 35774 3528
rect 36173 3519 36231 3525
rect 36173 3516 36185 3519
rect 35768 3488 36185 3516
rect 35768 3476 35774 3488
rect 36173 3485 36185 3488
rect 36219 3485 36231 3519
rect 36173 3479 36231 3485
rect 36262 3476 36268 3528
rect 36320 3516 36326 3528
rect 36817 3519 36875 3525
rect 36817 3516 36829 3519
rect 36320 3488 36829 3516
rect 36320 3476 36326 3488
rect 36817 3485 36829 3488
rect 36863 3485 36875 3519
rect 36817 3479 36875 3485
rect 37642 3476 37648 3528
rect 37700 3516 37706 3528
rect 38105 3519 38163 3525
rect 38105 3516 38117 3519
rect 37700 3488 38117 3516
rect 37700 3476 37706 3488
rect 38105 3485 38117 3488
rect 38151 3485 38163 3519
rect 38105 3479 38163 3485
rect 38194 3476 38200 3528
rect 38252 3516 38258 3528
rect 38749 3519 38807 3525
rect 38749 3516 38761 3519
rect 38252 3488 38761 3516
rect 38252 3476 38258 3488
rect 38749 3485 38761 3488
rect 38795 3485 38807 3519
rect 38749 3479 38807 3485
rect 39574 3476 39580 3528
rect 39632 3516 39638 3528
rect 40037 3519 40095 3525
rect 40037 3516 40049 3519
rect 39632 3488 40049 3516
rect 39632 3476 39638 3488
rect 40037 3485 40049 3488
rect 40083 3485 40095 3519
rect 40037 3479 40095 3485
rect 40402 3476 40408 3528
rect 40460 3516 40466 3528
rect 40681 3519 40739 3525
rect 40681 3516 40693 3519
rect 40460 3488 40693 3516
rect 40460 3476 40466 3488
rect 40681 3485 40693 3488
rect 40727 3485 40739 3519
rect 40681 3479 40739 3485
rect 40954 3476 40960 3528
rect 41012 3516 41018 3528
rect 41325 3519 41383 3525
rect 41325 3516 41337 3519
rect 41012 3488 41337 3516
rect 41012 3476 41018 3488
rect 41325 3485 41337 3488
rect 41371 3485 41383 3519
rect 41325 3479 41383 3485
rect 41506 3476 41512 3528
rect 41564 3516 41570 3528
rect 41969 3519 42027 3525
rect 41969 3516 41981 3519
rect 41564 3488 41981 3516
rect 41564 3476 41570 3488
rect 41969 3485 41981 3488
rect 42015 3485 42027 3519
rect 42886 3516 42892 3528
rect 42847 3488 42892 3516
rect 41969 3479 42027 3485
rect 42886 3476 42892 3488
rect 42944 3476 42950 3528
rect 43162 3476 43168 3528
rect 43220 3516 43226 3528
rect 43349 3519 43407 3525
rect 43349 3516 43361 3519
rect 43220 3488 43361 3516
rect 43220 3476 43226 3488
rect 43349 3485 43361 3488
rect 43395 3485 43407 3519
rect 43349 3479 43407 3485
rect 44818 3476 44824 3528
rect 44876 3516 44882 3528
rect 45189 3519 45247 3525
rect 45189 3516 45201 3519
rect 44876 3488 45201 3516
rect 44876 3476 44882 3488
rect 45189 3485 45201 3488
rect 45235 3485 45247 3519
rect 45189 3479 45247 3485
rect 45646 3476 45652 3528
rect 45704 3516 45710 3528
rect 45833 3519 45891 3525
rect 45833 3516 45845 3519
rect 45704 3488 45845 3516
rect 45704 3476 45710 3488
rect 45833 3485 45845 3488
rect 45879 3485 45891 3519
rect 46474 3516 46480 3528
rect 46435 3488 46480 3516
rect 45833 3479 45891 3485
rect 46474 3476 46480 3488
rect 46532 3476 46538 3528
rect 46750 3476 46756 3528
rect 46808 3516 46814 3528
rect 47121 3519 47179 3525
rect 47121 3516 47133 3519
rect 46808 3488 47133 3516
rect 46808 3476 46814 3488
rect 47121 3485 47133 3488
rect 47167 3485 47179 3519
rect 47121 3479 47179 3485
rect 47302 3476 47308 3528
rect 47360 3516 47366 3528
rect 47765 3519 47823 3525
rect 47765 3516 47777 3519
rect 47360 3488 47777 3516
rect 47360 3476 47366 3488
rect 47765 3485 47777 3488
rect 47811 3485 47823 3519
rect 47765 3479 47823 3485
rect 30926 3448 30932 3460
rect 29880 3420 30932 3448
rect 29880 3408 29886 3420
rect 30926 3408 30932 3420
rect 30984 3408 30990 3460
rect 28276 3352 28856 3380
rect 28902 3340 28908 3392
rect 28960 3380 28966 3392
rect 30469 3383 30527 3389
rect 30469 3380 30481 3383
rect 28960 3352 30481 3380
rect 28960 3340 28966 3352
rect 30469 3349 30481 3352
rect 30515 3349 30527 3383
rect 30469 3343 30527 3349
rect 1104 3290 48852 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 48852 3290
rect 1104 3216 48852 3238
rect 20070 3176 20076 3188
rect 17052 3148 20076 3176
rect 15013 3043 15071 3049
rect 15013 3009 15025 3043
rect 15059 3040 15071 3043
rect 16666 3040 16672 3052
rect 15059 3012 16672 3040
rect 15059 3009 15071 3012
rect 15013 3003 15071 3009
rect 16666 3000 16672 3012
rect 16724 3000 16730 3052
rect 17052 3049 17080 3148
rect 20070 3136 20076 3148
rect 20128 3136 20134 3188
rect 20165 3179 20223 3185
rect 20165 3145 20177 3179
rect 20211 3176 20223 3179
rect 20211 3148 24256 3176
rect 20211 3145 20223 3148
rect 20165 3139 20223 3145
rect 18233 3111 18291 3117
rect 18233 3077 18245 3111
rect 18279 3108 18291 3111
rect 20901 3111 20959 3117
rect 20901 3108 20913 3111
rect 18279 3080 20913 3108
rect 18279 3077 18291 3080
rect 18233 3071 18291 3077
rect 20901 3077 20913 3080
rect 20947 3077 20959 3111
rect 23014 3108 23020 3120
rect 22975 3080 23020 3108
rect 20901 3071 20959 3077
rect 23014 3068 23020 3080
rect 23072 3068 23078 3120
rect 24118 3108 24124 3120
rect 24079 3080 24124 3108
rect 24118 3068 24124 3080
rect 24176 3068 24182 3120
rect 24228 3117 24256 3148
rect 25038 3136 25044 3188
rect 25096 3176 25102 3188
rect 31018 3176 31024 3188
rect 25096 3148 27384 3176
rect 25096 3136 25102 3148
rect 27356 3117 27384 3148
rect 29012 3148 31024 3176
rect 24213 3111 24271 3117
rect 24213 3077 24225 3111
rect 24259 3077 24271 3111
rect 25961 3111 26019 3117
rect 25961 3108 25973 3111
rect 24213 3071 24271 3077
rect 24780 3080 25973 3108
rect 17037 3043 17095 3049
rect 17037 3009 17049 3043
rect 17083 3009 17095 3043
rect 17037 3003 17095 3009
rect 18325 3043 18383 3049
rect 18325 3009 18337 3043
rect 18371 3040 18383 3043
rect 18414 3040 18420 3052
rect 18371 3012 18420 3040
rect 18371 3009 18383 3012
rect 18325 3003 18383 3009
rect 18414 3000 18420 3012
rect 18472 3040 18478 3052
rect 19242 3040 19248 3052
rect 18472 3012 19248 3040
rect 18472 3000 18478 3012
rect 19242 3000 19248 3012
rect 19300 3040 19306 3052
rect 19429 3043 19487 3049
rect 19429 3040 19441 3043
rect 19300 3012 19441 3040
rect 19300 3000 19306 3012
rect 19429 3009 19441 3012
rect 19475 3009 19487 3043
rect 19429 3003 19487 3009
rect 20073 3043 20131 3049
rect 20073 3009 20085 3043
rect 20119 3040 20131 3043
rect 20162 3040 20168 3052
rect 20119 3012 20168 3040
rect 20119 3009 20131 3012
rect 20073 3003 20131 3009
rect 20162 3000 20168 3012
rect 20220 3040 20226 3052
rect 20622 3040 20628 3052
rect 20220 3012 20628 3040
rect 20220 3000 20226 3012
rect 20622 3000 20628 3012
rect 20680 3000 20686 3052
rect 22189 3043 22247 3049
rect 22189 3009 22201 3043
rect 22235 3009 22247 3043
rect 22189 3003 22247 3009
rect 4709 2975 4767 2981
rect 4709 2941 4721 2975
rect 4755 2972 4767 2975
rect 5442 2972 5448 2984
rect 4755 2944 5448 2972
rect 4755 2941 4767 2944
rect 4709 2935 4767 2941
rect 5442 2932 5448 2944
rect 5500 2932 5506 2984
rect 7285 2975 7343 2981
rect 7285 2941 7297 2975
rect 7331 2972 7343 2975
rect 7926 2972 7932 2984
rect 7331 2944 7932 2972
rect 7331 2941 7343 2944
rect 7285 2935 7343 2941
rect 7926 2932 7932 2944
rect 7984 2932 7990 2984
rect 9217 2975 9275 2981
rect 9217 2941 9229 2975
rect 9263 2972 9275 2975
rect 9858 2972 9864 2984
rect 9263 2944 9864 2972
rect 9263 2941 9275 2944
rect 9217 2935 9275 2941
rect 9858 2932 9864 2944
rect 9916 2932 9922 2984
rect 16301 2975 16359 2981
rect 16301 2941 16313 2975
rect 16347 2972 16359 2975
rect 17681 2975 17739 2981
rect 16347 2944 17632 2972
rect 16347 2941 16359 2944
rect 16301 2935 16359 2941
rect 4065 2907 4123 2913
rect 4065 2873 4077 2907
rect 4111 2904 4123 2907
rect 4890 2904 4896 2916
rect 4111 2876 4896 2904
rect 4111 2873 4123 2876
rect 4065 2867 4123 2873
rect 4890 2864 4896 2876
rect 4948 2864 4954 2916
rect 5353 2907 5411 2913
rect 5353 2873 5365 2907
rect 5399 2904 5411 2907
rect 6270 2904 6276 2916
rect 5399 2876 6276 2904
rect 5399 2873 5411 2876
rect 5353 2867 5411 2873
rect 6270 2864 6276 2876
rect 6328 2864 6334 2916
rect 8754 2904 8760 2916
rect 7944 2876 8760 2904
rect 2777 2839 2835 2845
rect 2777 2805 2789 2839
rect 2823 2836 2835 2839
rect 3142 2836 3148 2848
rect 2823 2808 3148 2836
rect 2823 2805 2835 2808
rect 2777 2799 2835 2805
rect 3142 2796 3148 2808
rect 3200 2796 3206 2848
rect 3421 2839 3479 2845
rect 3421 2805 3433 2839
rect 3467 2836 3479 2839
rect 3878 2836 3884 2848
rect 3467 2808 3884 2836
rect 3467 2805 3479 2808
rect 3421 2799 3479 2805
rect 3878 2796 3884 2808
rect 3936 2796 3942 2848
rect 5997 2839 6055 2845
rect 5997 2805 6009 2839
rect 6043 2836 6055 2839
rect 6546 2836 6552 2848
rect 6043 2808 6552 2836
rect 6043 2805 6055 2808
rect 5997 2799 6055 2805
rect 6546 2796 6552 2808
rect 6604 2796 6610 2848
rect 7944 2845 7972 2876
rect 8754 2864 8760 2876
rect 8812 2864 8818 2916
rect 10505 2907 10563 2913
rect 10505 2873 10517 2907
rect 10551 2904 10563 2907
rect 11238 2904 11244 2916
rect 10551 2876 11244 2904
rect 10551 2873 10563 2876
rect 10505 2867 10563 2873
rect 11238 2864 11244 2876
rect 11296 2864 11302 2916
rect 12437 2907 12495 2913
rect 12437 2873 12449 2907
rect 12483 2904 12495 2907
rect 13354 2904 13360 2916
rect 12483 2876 13360 2904
rect 12483 2873 12495 2876
rect 12437 2867 12495 2873
rect 13354 2864 13360 2876
rect 13412 2864 13418 2916
rect 13725 2907 13783 2913
rect 13725 2873 13737 2907
rect 13771 2904 13783 2907
rect 14458 2904 14464 2916
rect 13771 2876 14464 2904
rect 13771 2873 13783 2876
rect 13725 2867 13783 2873
rect 14458 2864 14464 2876
rect 14516 2864 14522 2916
rect 15657 2907 15715 2913
rect 15657 2873 15669 2907
rect 15703 2904 15715 2907
rect 17494 2904 17500 2916
rect 15703 2876 17500 2904
rect 15703 2873 15715 2876
rect 15657 2867 15715 2873
rect 17494 2864 17500 2876
rect 17552 2864 17558 2916
rect 17604 2904 17632 2944
rect 17681 2941 17693 2975
rect 17727 2972 17739 2975
rect 20809 2975 20867 2981
rect 20809 2972 20821 2975
rect 17727 2944 20821 2972
rect 17727 2941 17739 2944
rect 17681 2935 17739 2941
rect 20809 2941 20821 2944
rect 20855 2941 20867 2975
rect 20809 2935 20867 2941
rect 21453 2975 21511 2981
rect 21453 2941 21465 2975
rect 21499 2972 21511 2975
rect 21634 2972 21640 2984
rect 21499 2944 21640 2972
rect 21499 2941 21511 2944
rect 21453 2935 21511 2941
rect 21634 2932 21640 2944
rect 21692 2932 21698 2984
rect 18782 2904 18788 2916
rect 17604 2876 18788 2904
rect 18782 2864 18788 2876
rect 18840 2864 18846 2916
rect 19521 2907 19579 2913
rect 19521 2873 19533 2907
rect 19567 2904 19579 2907
rect 22002 2904 22008 2916
rect 19567 2876 22008 2904
rect 19567 2873 19579 2876
rect 19521 2867 19579 2873
rect 22002 2864 22008 2876
rect 22060 2864 22066 2916
rect 7929 2839 7987 2845
rect 7929 2805 7941 2839
rect 7975 2805 7987 2839
rect 7929 2799 7987 2805
rect 8573 2839 8631 2845
rect 8573 2805 8585 2839
rect 8619 2836 8631 2839
rect 9030 2836 9036 2848
rect 8619 2808 9036 2836
rect 8619 2805 8631 2808
rect 8573 2799 8631 2805
rect 9030 2796 9036 2808
rect 9088 2796 9094 2848
rect 9861 2839 9919 2845
rect 9861 2805 9873 2839
rect 9907 2836 9919 2839
rect 10686 2836 10692 2848
rect 9907 2808 10692 2836
rect 9907 2805 9919 2808
rect 9861 2799 9919 2805
rect 10686 2796 10692 2808
rect 10744 2796 10750 2848
rect 11149 2839 11207 2845
rect 11149 2805 11161 2839
rect 11195 2836 11207 2839
rect 12066 2836 12072 2848
rect 11195 2808 12072 2836
rect 11195 2805 11207 2808
rect 11149 2799 11207 2805
rect 12066 2796 12072 2808
rect 12124 2796 12130 2848
rect 13081 2839 13139 2845
rect 13081 2805 13093 2839
rect 13127 2836 13139 2839
rect 13906 2836 13912 2848
rect 13127 2808 13912 2836
rect 13127 2805 13139 2808
rect 13081 2799 13139 2805
rect 13906 2796 13912 2808
rect 13964 2796 13970 2848
rect 14369 2839 14427 2845
rect 14369 2805 14381 2839
rect 14415 2836 14427 2839
rect 15286 2836 15292 2848
rect 14415 2808 15292 2836
rect 14415 2805 14427 2808
rect 14369 2799 14427 2805
rect 15286 2796 15292 2808
rect 15344 2796 15350 2848
rect 15378 2796 15384 2848
rect 15436 2836 15442 2848
rect 17770 2836 17776 2848
rect 15436 2808 17776 2836
rect 15436 2796 15442 2808
rect 17770 2796 17776 2808
rect 17828 2796 17834 2848
rect 18966 2836 18972 2848
rect 18927 2808 18972 2836
rect 18966 2796 18972 2808
rect 19024 2796 19030 2848
rect 20070 2796 20076 2848
rect 20128 2836 20134 2848
rect 20530 2836 20536 2848
rect 20128 2808 20536 2836
rect 20128 2796 20134 2808
rect 20530 2796 20536 2808
rect 20588 2796 20594 2848
rect 20622 2796 20628 2848
rect 20680 2836 20686 2848
rect 22204 2836 22232 3003
rect 22370 2932 22376 2984
rect 22428 2972 22434 2984
rect 22925 2975 22983 2981
rect 22925 2972 22937 2975
rect 22428 2944 22937 2972
rect 22428 2932 22434 2944
rect 22925 2941 22937 2944
rect 22971 2941 22983 2975
rect 22925 2935 22983 2941
rect 23569 2975 23627 2981
rect 23569 2941 23581 2975
rect 23615 2972 23627 2975
rect 23842 2972 23848 2984
rect 23615 2944 23848 2972
rect 23615 2941 23627 2944
rect 23569 2935 23627 2941
rect 23842 2932 23848 2944
rect 23900 2932 23906 2984
rect 24394 2972 24400 2984
rect 24355 2944 24400 2972
rect 24394 2932 24400 2944
rect 24452 2932 24458 2984
rect 22281 2907 22339 2913
rect 22281 2873 22293 2907
rect 22327 2904 22339 2907
rect 24780 2904 24808 3080
rect 25961 3077 25973 3080
rect 26007 3077 26019 3111
rect 25961 3071 26019 3077
rect 27341 3111 27399 3117
rect 27341 3077 27353 3111
rect 27387 3077 27399 3111
rect 28902 3108 28908 3120
rect 28863 3080 28908 3108
rect 27341 3071 27399 3077
rect 28902 3068 28908 3080
rect 28960 3068 28966 3120
rect 29012 3117 29040 3148
rect 31018 3136 31024 3148
rect 31076 3136 31082 3188
rect 28997 3111 29055 3117
rect 28997 3077 29009 3111
rect 29043 3077 29055 3111
rect 28997 3071 29055 3077
rect 30101 3111 30159 3117
rect 30101 3077 30113 3111
rect 30147 3108 30159 3111
rect 31481 3111 31539 3117
rect 31481 3108 31493 3111
rect 30147 3080 31493 3108
rect 30147 3077 30159 3080
rect 30101 3071 30159 3077
rect 31481 3077 31493 3080
rect 31527 3077 31539 3111
rect 31481 3071 31539 3077
rect 30926 3000 30932 3052
rect 30984 3040 30990 3052
rect 31389 3043 31447 3049
rect 31389 3040 31401 3043
rect 30984 3012 31401 3040
rect 30984 3000 30990 3012
rect 31389 3009 31401 3012
rect 31435 3009 31447 3043
rect 31389 3003 31447 3009
rect 32674 3000 32680 3052
rect 32732 3040 32738 3052
rect 34241 3043 34299 3049
rect 34241 3040 34253 3043
rect 32732 3012 34253 3040
rect 32732 3000 32738 3012
rect 34241 3009 34253 3012
rect 34287 3009 34299 3043
rect 34241 3003 34299 3009
rect 25774 2972 25780 2984
rect 25735 2944 25780 2972
rect 25774 2932 25780 2944
rect 25832 2932 25838 2984
rect 26053 2975 26111 2981
rect 26053 2941 26065 2975
rect 26099 2941 26111 2975
rect 27246 2972 27252 2984
rect 27207 2944 27252 2972
rect 26053 2935 26111 2941
rect 22327 2876 24808 2904
rect 22327 2873 22339 2876
rect 22281 2867 22339 2873
rect 23658 2836 23664 2848
rect 20680 2808 23664 2836
rect 20680 2796 20686 2808
rect 23658 2796 23664 2808
rect 23716 2796 23722 2848
rect 26068 2836 26096 2935
rect 27246 2932 27252 2944
rect 27304 2932 27310 2984
rect 27525 2975 27583 2981
rect 27525 2941 27537 2975
rect 27571 2941 27583 2975
rect 28534 2972 28540 2984
rect 28495 2944 28540 2972
rect 27525 2935 27583 2941
rect 26878 2864 26884 2916
rect 26936 2904 26942 2916
rect 27540 2904 27568 2935
rect 28534 2932 28540 2944
rect 28592 2932 28598 2984
rect 29362 2932 29368 2984
rect 29420 2972 29426 2984
rect 29549 2975 29607 2981
rect 29549 2972 29561 2975
rect 29420 2944 29561 2972
rect 29420 2932 29426 2944
rect 29549 2941 29561 2944
rect 29595 2941 29607 2975
rect 29549 2935 29607 2941
rect 30193 2975 30251 2981
rect 30193 2941 30205 2975
rect 30239 2972 30251 2975
rect 31662 2972 31668 2984
rect 30239 2944 31668 2972
rect 30239 2941 30251 2944
rect 30193 2935 30251 2941
rect 31662 2932 31668 2944
rect 31720 2932 31726 2984
rect 32122 2932 32128 2984
rect 32180 2972 32186 2984
rect 33597 2975 33655 2981
rect 33597 2972 33609 2975
rect 32180 2944 33609 2972
rect 32180 2932 32186 2944
rect 33597 2941 33609 2944
rect 33643 2941 33655 2975
rect 33597 2935 33655 2941
rect 34054 2932 34060 2984
rect 34112 2972 34118 2984
rect 35529 2975 35587 2981
rect 35529 2972 35541 2975
rect 34112 2944 35541 2972
rect 34112 2932 34118 2944
rect 35529 2941 35541 2944
rect 35575 2941 35587 2975
rect 35529 2935 35587 2941
rect 37090 2932 37096 2984
rect 37148 2972 37154 2984
rect 38105 2975 38163 2981
rect 38105 2972 38117 2975
rect 37148 2944 38117 2972
rect 37148 2932 37154 2944
rect 38105 2941 38117 2944
rect 38151 2941 38163 2975
rect 38105 2935 38163 2941
rect 38746 2932 38752 2984
rect 38804 2972 38810 2984
rect 39393 2975 39451 2981
rect 39393 2972 39405 2975
rect 38804 2944 39405 2972
rect 38804 2932 38810 2944
rect 39393 2941 39405 2944
rect 39439 2941 39451 2975
rect 39393 2935 39451 2941
rect 40678 2932 40684 2984
rect 40736 2972 40742 2984
rect 41325 2975 41383 2981
rect 41325 2972 41337 2975
rect 40736 2944 41337 2972
rect 40736 2932 40742 2944
rect 41325 2941 41337 2944
rect 41371 2941 41383 2975
rect 41325 2935 41383 2941
rect 42610 2932 42616 2984
rect 42668 2972 42674 2984
rect 43257 2975 43315 2981
rect 43257 2972 43269 2975
rect 42668 2944 43269 2972
rect 42668 2932 42674 2944
rect 43257 2941 43269 2944
rect 43303 2941 43315 2975
rect 43257 2935 43315 2941
rect 44542 2932 44548 2984
rect 44600 2972 44606 2984
rect 45189 2975 45247 2981
rect 45189 2972 45201 2975
rect 44600 2944 45201 2972
rect 44600 2932 44606 2944
rect 45189 2941 45201 2944
rect 45235 2941 45247 2975
rect 45189 2935 45247 2941
rect 26936 2876 27568 2904
rect 26936 2864 26942 2876
rect 28350 2864 28356 2916
rect 28408 2904 28414 2916
rect 30745 2907 30803 2913
rect 30745 2904 30757 2907
rect 28408 2876 30757 2904
rect 28408 2864 28414 2876
rect 30745 2873 30757 2876
rect 30791 2873 30803 2907
rect 30745 2867 30803 2873
rect 30834 2864 30840 2916
rect 30892 2864 30898 2916
rect 31570 2864 31576 2916
rect 31628 2904 31634 2916
rect 32953 2907 33011 2913
rect 32953 2904 32965 2907
rect 31628 2876 32965 2904
rect 31628 2864 31634 2876
rect 32953 2873 32965 2876
rect 32999 2873 33011 2907
rect 32953 2867 33011 2873
rect 33502 2864 33508 2916
rect 33560 2904 33566 2916
rect 34885 2907 34943 2913
rect 34885 2904 34897 2907
rect 33560 2876 34897 2904
rect 33560 2864 33566 2876
rect 34885 2873 34897 2876
rect 34931 2873 34943 2907
rect 34885 2867 34943 2873
rect 35342 2864 35348 2916
rect 35400 2904 35406 2916
rect 36173 2907 36231 2913
rect 36173 2904 36185 2907
rect 35400 2876 36185 2904
rect 35400 2864 35406 2876
rect 36173 2873 36185 2876
rect 36219 2873 36231 2907
rect 36173 2867 36231 2873
rect 37918 2864 37924 2916
rect 37976 2904 37982 2916
rect 37976 2876 38792 2904
rect 37976 2864 37982 2876
rect 29730 2836 29736 2848
rect 26068 2808 29736 2836
rect 29730 2796 29736 2808
rect 29788 2796 29794 2848
rect 30852 2836 30880 2864
rect 32309 2839 32367 2845
rect 32309 2836 32321 2839
rect 30852 2808 32321 2836
rect 32309 2805 32321 2808
rect 32355 2805 32367 2839
rect 32309 2799 32367 2805
rect 35986 2796 35992 2848
rect 36044 2836 36050 2848
rect 38764 2845 38792 2876
rect 37461 2839 37519 2845
rect 37461 2836 37473 2839
rect 36044 2808 37473 2836
rect 36044 2796 36050 2808
rect 37461 2805 37473 2808
rect 37507 2805 37519 2839
rect 37461 2799 37519 2805
rect 38749 2839 38807 2845
rect 38749 2805 38761 2839
rect 38795 2805 38807 2839
rect 38749 2799 38807 2805
rect 39022 2796 39028 2848
rect 39080 2836 39086 2848
rect 40037 2839 40095 2845
rect 40037 2836 40049 2839
rect 39080 2808 40049 2836
rect 39080 2796 39086 2808
rect 40037 2805 40049 2808
rect 40083 2805 40095 2839
rect 40037 2799 40095 2805
rect 40126 2796 40132 2848
rect 40184 2836 40190 2848
rect 40681 2839 40739 2845
rect 40681 2836 40693 2839
rect 40184 2808 40693 2836
rect 40184 2796 40190 2808
rect 40681 2805 40693 2808
rect 40727 2805 40739 2839
rect 40681 2799 40739 2805
rect 42058 2796 42064 2848
rect 42116 2836 42122 2848
rect 42613 2839 42671 2845
rect 42613 2836 42625 2839
rect 42116 2808 42625 2836
rect 42116 2796 42122 2808
rect 42613 2805 42625 2808
rect 42659 2805 42671 2839
rect 42613 2799 42671 2805
rect 43438 2796 43444 2848
rect 43496 2836 43502 2848
rect 43901 2839 43959 2845
rect 43901 2836 43913 2839
rect 43496 2808 43913 2836
rect 43496 2796 43502 2808
rect 43901 2805 43913 2808
rect 43947 2805 43959 2839
rect 43901 2799 43959 2805
rect 43990 2796 43996 2848
rect 44048 2836 44054 2848
rect 44545 2839 44603 2845
rect 44545 2836 44557 2839
rect 44048 2808 44557 2836
rect 44048 2796 44054 2808
rect 44545 2805 44557 2808
rect 44591 2805 44603 2839
rect 44545 2799 44603 2805
rect 45370 2796 45376 2848
rect 45428 2836 45434 2848
rect 45833 2839 45891 2845
rect 45833 2836 45845 2839
rect 45428 2808 45845 2836
rect 45428 2796 45434 2808
rect 45833 2805 45845 2808
rect 45879 2805 45891 2839
rect 45833 2799 45891 2805
rect 45922 2796 45928 2848
rect 45980 2836 45986 2848
rect 46477 2839 46535 2845
rect 46477 2836 46489 2839
rect 45980 2808 46489 2836
rect 45980 2796 45986 2808
rect 46477 2805 46489 2808
rect 46523 2805 46535 2839
rect 46477 2799 46535 2805
rect 47026 2796 47032 2848
rect 47084 2836 47090 2848
rect 47765 2839 47823 2845
rect 47765 2836 47777 2839
rect 47084 2808 47777 2836
rect 47084 2796 47090 2808
rect 47765 2805 47777 2808
rect 47811 2805 47823 2839
rect 47765 2799 47823 2805
rect 1104 2746 48852 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 48852 2746
rect 1104 2672 48852 2694
rect 15013 2635 15071 2641
rect 15013 2601 15025 2635
rect 15059 2632 15071 2635
rect 15378 2632 15384 2644
rect 15059 2604 15384 2632
rect 15059 2601 15071 2604
rect 15013 2595 15071 2601
rect 15378 2592 15384 2604
rect 15436 2592 15442 2644
rect 19613 2635 19671 2641
rect 19613 2601 19625 2635
rect 19659 2632 19671 2635
rect 23937 2635 23995 2641
rect 19659 2604 23244 2632
rect 19659 2601 19671 2604
rect 19613 2595 19671 2601
rect 5353 2567 5411 2573
rect 5353 2533 5365 2567
rect 5399 2564 5411 2567
rect 7098 2564 7104 2576
rect 5399 2536 7104 2564
rect 5399 2533 5411 2536
rect 5353 2527 5411 2533
rect 7098 2524 7104 2536
rect 7156 2524 7162 2576
rect 7929 2567 7987 2573
rect 7929 2533 7941 2567
rect 7975 2564 7987 2567
rect 9582 2564 9588 2576
rect 7975 2536 9588 2564
rect 7975 2533 7987 2536
rect 7929 2527 7987 2533
rect 9582 2524 9588 2536
rect 9640 2524 9646 2576
rect 9861 2567 9919 2573
rect 9861 2533 9873 2567
rect 9907 2564 9919 2567
rect 11514 2564 11520 2576
rect 9907 2536 11520 2564
rect 9907 2533 9919 2536
rect 9861 2527 9919 2533
rect 11514 2524 11520 2536
rect 11572 2524 11578 2576
rect 12437 2567 12495 2573
rect 12437 2533 12449 2567
rect 12483 2564 12495 2567
rect 14182 2564 14188 2576
rect 12483 2536 14188 2564
rect 12483 2533 12495 2536
rect 12437 2527 12495 2533
rect 14182 2524 14188 2536
rect 14240 2524 14246 2576
rect 15657 2567 15715 2573
rect 15657 2533 15669 2567
rect 15703 2564 15715 2567
rect 18322 2564 18328 2576
rect 15703 2536 18328 2564
rect 15703 2533 15715 2536
rect 15657 2527 15715 2533
rect 18322 2524 18328 2536
rect 18380 2524 18386 2576
rect 20165 2567 20223 2573
rect 20165 2533 20177 2567
rect 20211 2564 20223 2567
rect 20211 2536 23152 2564
rect 20211 2533 20223 2536
rect 20165 2527 20223 2533
rect 2777 2499 2835 2505
rect 2777 2465 2789 2499
rect 2823 2496 2835 2499
rect 3510 2496 3516 2508
rect 2823 2468 3516 2496
rect 2823 2465 2835 2468
rect 2777 2459 2835 2465
rect 3510 2456 3516 2468
rect 3568 2456 3574 2508
rect 7285 2499 7343 2505
rect 7285 2465 7297 2499
rect 7331 2496 7343 2499
rect 8202 2496 8208 2508
rect 7331 2468 8208 2496
rect 7331 2465 7343 2468
rect 7285 2459 7343 2465
rect 8202 2456 8208 2468
rect 8260 2456 8266 2508
rect 8573 2499 8631 2505
rect 8573 2465 8585 2499
rect 8619 2496 8631 2499
rect 10410 2496 10416 2508
rect 8619 2468 10416 2496
rect 8619 2465 8631 2468
rect 8573 2459 8631 2465
rect 10410 2456 10416 2468
rect 10468 2456 10474 2508
rect 11149 2499 11207 2505
rect 11149 2465 11161 2499
rect 11195 2496 11207 2499
rect 12802 2496 12808 2508
rect 11195 2468 12808 2496
rect 11195 2465 11207 2468
rect 11149 2459 11207 2465
rect 12802 2456 12808 2468
rect 12860 2456 12866 2508
rect 13081 2499 13139 2505
rect 13081 2465 13093 2499
rect 13127 2496 13139 2499
rect 14734 2496 14740 2508
rect 13127 2468 14740 2496
rect 13127 2465 13139 2468
rect 13081 2459 13139 2465
rect 14734 2456 14740 2468
rect 14792 2456 14798 2508
rect 17589 2499 17647 2505
rect 17589 2465 17601 2499
rect 17635 2496 17647 2499
rect 20809 2499 20867 2505
rect 20809 2496 20821 2499
rect 17635 2468 20821 2496
rect 17635 2465 17647 2468
rect 17589 2459 17647 2465
rect 20809 2465 20821 2468
rect 20855 2465 20867 2499
rect 20809 2459 20867 2465
rect 22278 2456 22284 2508
rect 22336 2496 22342 2508
rect 22465 2499 22523 2505
rect 22465 2496 22477 2499
rect 22336 2468 22477 2496
rect 22336 2456 22342 2468
rect 22465 2465 22477 2468
rect 22511 2465 22523 2499
rect 22738 2496 22744 2508
rect 22699 2468 22744 2496
rect 22465 2459 22523 2465
rect 22738 2456 22744 2468
rect 22796 2456 22802 2508
rect 2133 2431 2191 2437
rect 2133 2397 2145 2431
rect 2179 2428 2191 2431
rect 2590 2428 2596 2440
rect 2179 2400 2596 2428
rect 2179 2397 2191 2400
rect 2133 2391 2191 2397
rect 2590 2388 2596 2400
rect 2648 2388 2654 2440
rect 3421 2431 3479 2437
rect 3421 2397 3433 2431
rect 3467 2428 3479 2431
rect 4614 2428 4620 2440
rect 3467 2400 4620 2428
rect 3467 2397 3479 2400
rect 3421 2391 3479 2397
rect 4614 2388 4620 2400
rect 4672 2388 4678 2440
rect 4709 2431 4767 2437
rect 4709 2397 4721 2431
rect 4755 2428 4767 2431
rect 5718 2428 5724 2440
rect 4755 2400 5724 2428
rect 4755 2397 4767 2400
rect 4709 2391 4767 2397
rect 5718 2388 5724 2400
rect 5776 2388 5782 2440
rect 5997 2431 6055 2437
rect 5997 2397 6009 2431
rect 6043 2428 6055 2431
rect 10505 2431 10563 2437
rect 6043 2400 6914 2428
rect 6043 2397 6055 2400
rect 5997 2391 6055 2397
rect 6886 2360 6914 2400
rect 10505 2397 10517 2431
rect 10551 2428 10563 2431
rect 12250 2428 12256 2440
rect 10551 2400 12256 2428
rect 10551 2397 10563 2400
rect 10505 2391 10563 2397
rect 12250 2388 12256 2400
rect 12308 2388 12314 2440
rect 13725 2431 13783 2437
rect 13725 2397 13737 2431
rect 13771 2428 13783 2431
rect 15562 2428 15568 2440
rect 13771 2400 15568 2428
rect 13771 2397 13783 2400
rect 13725 2391 13783 2397
rect 15562 2388 15568 2400
rect 15620 2388 15626 2440
rect 16298 2428 16304 2440
rect 16259 2400 16304 2428
rect 16298 2388 16304 2400
rect 16356 2388 16362 2440
rect 18233 2431 18291 2437
rect 18233 2397 18245 2431
rect 18279 2428 18291 2431
rect 18414 2428 18420 2440
rect 18279 2400 18420 2428
rect 18279 2397 18291 2400
rect 18233 2391 18291 2397
rect 18414 2388 18420 2400
rect 18472 2388 18478 2440
rect 18874 2428 18880 2440
rect 18835 2400 18880 2428
rect 18874 2388 18880 2400
rect 18932 2388 18938 2440
rect 20073 2431 20131 2437
rect 20073 2397 20085 2431
rect 20119 2428 20131 2431
rect 20162 2428 20168 2440
rect 20119 2400 20168 2428
rect 20119 2397 20131 2400
rect 20073 2391 20131 2397
rect 20162 2388 20168 2400
rect 20220 2388 20226 2440
rect 7374 2360 7380 2372
rect 6886 2332 7380 2360
rect 7374 2320 7380 2332
rect 7432 2320 7438 2372
rect 18141 2363 18199 2369
rect 18141 2329 18153 2363
rect 18187 2360 18199 2363
rect 20901 2363 20959 2369
rect 18187 2332 20760 2360
rect 18187 2329 18199 2332
rect 18141 2323 18199 2329
rect 20732 2292 20760 2332
rect 20901 2329 20913 2363
rect 20947 2329 20959 2363
rect 20901 2323 20959 2329
rect 21453 2363 21511 2369
rect 21453 2329 21465 2363
rect 21499 2360 21511 2363
rect 21910 2360 21916 2372
rect 21499 2332 21916 2360
rect 21499 2329 21511 2332
rect 21453 2323 21511 2329
rect 20916 2292 20944 2323
rect 21910 2320 21916 2332
rect 21968 2320 21974 2372
rect 22557 2363 22615 2369
rect 22557 2329 22569 2363
rect 22603 2329 22615 2363
rect 22557 2323 22615 2329
rect 20732 2264 20944 2292
rect 22002 2252 22008 2304
rect 22060 2292 22066 2304
rect 22572 2292 22600 2323
rect 22060 2264 22600 2292
rect 23124 2292 23152 2536
rect 23216 2360 23244 2604
rect 23937 2601 23949 2635
rect 23983 2632 23995 2635
rect 24302 2632 24308 2644
rect 23983 2604 24308 2632
rect 23983 2601 23995 2604
rect 23937 2595 23995 2601
rect 24302 2592 24308 2604
rect 24360 2592 24366 2644
rect 26329 2635 26387 2641
rect 26329 2601 26341 2635
rect 26375 2632 26387 2635
rect 27246 2632 27252 2644
rect 26375 2604 27252 2632
rect 26375 2601 26387 2604
rect 26329 2595 26387 2601
rect 27246 2592 27252 2604
rect 27304 2592 27310 2644
rect 29730 2632 29736 2644
rect 29691 2604 29736 2632
rect 29730 2592 29736 2604
rect 29788 2592 29794 2644
rect 30282 2592 30288 2644
rect 30340 2632 30346 2644
rect 30469 2635 30527 2641
rect 30469 2632 30481 2635
rect 30340 2604 30481 2632
rect 30340 2592 30346 2604
rect 30469 2601 30481 2604
rect 30515 2601 30527 2635
rect 31018 2632 31024 2644
rect 30979 2604 31024 2632
rect 30469 2595 30527 2601
rect 31018 2592 31024 2604
rect 31076 2592 31082 2644
rect 31662 2592 31668 2644
rect 31720 2632 31726 2644
rect 32309 2635 32367 2641
rect 32309 2632 32321 2635
rect 31720 2604 32321 2632
rect 31720 2592 31726 2604
rect 32309 2601 32321 2604
rect 32355 2601 32367 2635
rect 32309 2595 32367 2601
rect 33226 2524 33232 2576
rect 33284 2564 33290 2576
rect 34885 2567 34943 2573
rect 34885 2564 34897 2567
rect 33284 2536 34897 2564
rect 33284 2524 33290 2536
rect 34885 2533 34897 2536
rect 34931 2533 34943 2567
rect 34885 2527 34943 2533
rect 35434 2524 35440 2576
rect 35492 2564 35498 2576
rect 37461 2567 37519 2573
rect 37461 2564 37473 2567
rect 35492 2536 37473 2564
rect 35492 2524 35498 2536
rect 37461 2533 37473 2536
rect 37507 2533 37519 2567
rect 37461 2527 37519 2533
rect 38470 2524 38476 2576
rect 38528 2564 38534 2576
rect 40037 2567 40095 2573
rect 40037 2564 40049 2567
rect 38528 2536 40049 2564
rect 38528 2524 38534 2536
rect 40037 2533 40049 2536
rect 40083 2533 40095 2567
rect 40037 2527 40095 2533
rect 42334 2524 42340 2576
rect 42392 2564 42398 2576
rect 43901 2567 43959 2573
rect 43901 2564 43913 2567
rect 42392 2536 43913 2564
rect 42392 2524 42398 2536
rect 43901 2533 43913 2536
rect 43947 2533 43959 2567
rect 43901 2527 43959 2533
rect 45094 2524 45100 2576
rect 45152 2564 45158 2576
rect 46477 2567 46535 2573
rect 46477 2564 46489 2567
rect 45152 2536 46489 2564
rect 45152 2524 45158 2536
rect 46477 2533 46489 2536
rect 46523 2533 46535 2567
rect 46477 2527 46535 2533
rect 24118 2456 24124 2508
rect 24176 2496 24182 2508
rect 24949 2499 25007 2505
rect 24949 2496 24961 2499
rect 24176 2468 24961 2496
rect 24176 2456 24182 2468
rect 24949 2465 24961 2468
rect 24995 2465 25007 2499
rect 24949 2459 25007 2465
rect 27801 2499 27859 2505
rect 27801 2465 27813 2499
rect 27847 2496 27859 2499
rect 28353 2499 28411 2505
rect 28353 2496 28365 2499
rect 27847 2468 28365 2496
rect 27847 2465 27859 2468
rect 27801 2459 27859 2465
rect 28353 2465 28365 2468
rect 28399 2465 28411 2499
rect 28353 2459 28411 2465
rect 31294 2456 31300 2508
rect 31352 2496 31358 2508
rect 33597 2499 33655 2505
rect 33597 2496 33609 2499
rect 31352 2468 33609 2496
rect 31352 2456 31358 2468
rect 33597 2465 33609 2468
rect 33643 2465 33655 2499
rect 33597 2459 33655 2465
rect 34606 2456 34612 2508
rect 34664 2496 34670 2508
rect 36173 2499 36231 2505
rect 36173 2496 36185 2499
rect 34664 2468 36185 2496
rect 34664 2456 34670 2468
rect 36173 2465 36185 2468
rect 36219 2465 36231 2499
rect 36173 2459 36231 2465
rect 37366 2456 37372 2508
rect 37424 2496 37430 2508
rect 38749 2499 38807 2505
rect 38749 2496 38761 2499
rect 37424 2468 38761 2496
rect 37424 2456 37430 2468
rect 38749 2465 38761 2468
rect 38795 2465 38807 2499
rect 38749 2459 38807 2465
rect 39298 2456 39304 2508
rect 39356 2496 39362 2508
rect 40681 2499 40739 2505
rect 40681 2496 40693 2499
rect 39356 2468 40693 2496
rect 39356 2456 39362 2468
rect 40681 2465 40693 2468
rect 40727 2465 40739 2499
rect 40681 2459 40739 2465
rect 41230 2456 41236 2508
rect 41288 2496 41294 2508
rect 42613 2499 42671 2505
rect 42613 2496 42625 2499
rect 41288 2468 42625 2496
rect 41288 2456 41294 2468
rect 42613 2465 42625 2468
rect 42659 2465 42671 2499
rect 42613 2459 42671 2465
rect 43714 2456 43720 2508
rect 43772 2496 43778 2508
rect 45189 2499 45247 2505
rect 45189 2496 45201 2499
rect 43772 2468 45201 2496
rect 43772 2456 43778 2468
rect 45189 2465 45201 2468
rect 45235 2465 45247 2499
rect 45189 2459 45247 2465
rect 23658 2388 23664 2440
rect 23716 2428 23722 2440
rect 23845 2431 23903 2437
rect 23845 2428 23857 2431
rect 23716 2400 23857 2428
rect 23716 2388 23722 2400
rect 23845 2397 23857 2400
rect 23891 2397 23903 2431
rect 23845 2391 23903 2397
rect 29181 2431 29239 2437
rect 29181 2397 29193 2431
rect 29227 2428 29239 2431
rect 30561 2431 30619 2437
rect 30561 2428 30573 2431
rect 29227 2400 30573 2428
rect 29227 2397 29239 2400
rect 29181 2391 29239 2397
rect 30561 2397 30573 2400
rect 30607 2428 30619 2431
rect 30834 2428 30840 2440
rect 30607 2400 30840 2428
rect 30607 2397 30619 2400
rect 30561 2391 30619 2397
rect 30834 2388 30840 2400
rect 30892 2388 30898 2440
rect 32953 2431 33011 2437
rect 32953 2397 32965 2431
rect 32999 2397 33011 2431
rect 32953 2391 33011 2397
rect 24673 2363 24731 2369
rect 24673 2360 24685 2363
rect 23216 2332 24685 2360
rect 24673 2329 24685 2332
rect 24719 2329 24731 2363
rect 24673 2323 24731 2329
rect 24765 2363 24823 2369
rect 24765 2329 24777 2363
rect 24811 2329 24823 2363
rect 27154 2360 27160 2372
rect 27115 2332 27160 2360
rect 24765 2323 24823 2329
rect 24780 2292 24808 2323
rect 27154 2320 27160 2332
rect 27212 2320 27218 2372
rect 27709 2363 27767 2369
rect 27709 2329 27721 2363
rect 27755 2360 27767 2363
rect 29089 2363 29147 2369
rect 29089 2360 29101 2363
rect 27755 2332 29101 2360
rect 27755 2329 27767 2332
rect 27709 2323 27767 2329
rect 29089 2329 29101 2332
rect 29135 2329 29147 2363
rect 29089 2323 29147 2329
rect 30466 2320 30472 2372
rect 30524 2360 30530 2372
rect 32968 2360 32996 2391
rect 33778 2388 33784 2440
rect 33836 2428 33842 2440
rect 35529 2431 35587 2437
rect 35529 2428 35541 2431
rect 33836 2400 35541 2428
rect 33836 2388 33842 2400
rect 35529 2397 35541 2400
rect 35575 2397 35587 2431
rect 35529 2391 35587 2397
rect 36538 2388 36544 2440
rect 36596 2428 36602 2440
rect 38105 2431 38163 2437
rect 38105 2428 38117 2431
rect 36596 2400 38117 2428
rect 36596 2388 36602 2400
rect 38105 2397 38117 2400
rect 38151 2397 38163 2431
rect 38105 2391 38163 2397
rect 39850 2388 39856 2440
rect 39908 2428 39914 2440
rect 41325 2431 41383 2437
rect 41325 2428 41337 2431
rect 39908 2400 41337 2428
rect 39908 2388 39914 2400
rect 41325 2397 41337 2400
rect 41371 2397 41383 2431
rect 41325 2391 41383 2397
rect 41782 2388 41788 2440
rect 41840 2428 41846 2440
rect 43257 2431 43315 2437
rect 43257 2428 43269 2431
rect 41840 2400 43269 2428
rect 41840 2388 41846 2400
rect 43257 2397 43269 2400
rect 43303 2397 43315 2431
rect 45833 2431 45891 2437
rect 45833 2428 45845 2431
rect 43257 2391 43315 2397
rect 45526 2400 45845 2428
rect 30524 2332 32996 2360
rect 30524 2320 30530 2332
rect 44266 2320 44272 2372
rect 44324 2360 44330 2372
rect 45526 2360 45554 2400
rect 45833 2397 45845 2400
rect 45879 2397 45891 2431
rect 45833 2391 45891 2397
rect 46198 2388 46204 2440
rect 46256 2428 46262 2440
rect 47765 2431 47823 2437
rect 47765 2428 47777 2431
rect 46256 2400 47777 2428
rect 46256 2388 46262 2400
rect 47765 2397 47777 2400
rect 47811 2397 47823 2431
rect 47765 2391 47823 2397
rect 44324 2332 45554 2360
rect 44324 2320 44330 2332
rect 23124 2264 24808 2292
rect 22060 2252 22066 2264
rect 1104 2202 48852 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 48852 2202
rect 1104 2128 48852 2150
rect 18874 2048 18880 2100
rect 18932 2088 18938 2100
rect 22370 2088 22376 2100
rect 18932 2060 22376 2088
rect 18932 2048 18938 2060
rect 22370 2048 22376 2060
rect 22428 2048 22434 2100
rect 16298 1912 16304 1964
rect 16356 1952 16362 1964
rect 19978 1952 19984 1964
rect 16356 1924 19984 1952
rect 16356 1912 16362 1924
rect 19978 1912 19984 1924
rect 20036 1912 20042 1964
<< via1 >>
rect 29000 47608 29052 47660
rect 32956 47608 33008 47660
rect 19432 47540 19484 47592
rect 20260 47540 20312 47592
rect 21916 47540 21968 47592
rect 22100 47540 22152 47592
rect 26792 47540 26844 47592
rect 28816 47540 28868 47592
rect 19892 47472 19944 47524
rect 33324 47540 33376 47592
rect 34152 47472 34204 47524
rect 37740 47472 37792 47524
rect 38752 47472 38804 47524
rect 38844 47472 38896 47524
rect 40776 47472 40828 47524
rect 18880 47404 18932 47456
rect 23480 47404 23532 47456
rect 24124 47404 24176 47456
rect 30196 47404 30248 47456
rect 35348 47404 35400 47456
rect 39764 47404 39816 47456
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 4712 47243 4764 47252
rect 4712 47209 4721 47243
rect 4721 47209 4755 47243
rect 4755 47209 4764 47243
rect 4712 47200 4764 47209
rect 5816 47200 5868 47252
rect 6000 47243 6052 47252
rect 6000 47209 6009 47243
rect 6009 47209 6043 47243
rect 6043 47209 6052 47243
rect 6000 47200 6052 47209
rect 7104 47243 7156 47252
rect 7104 47209 7113 47243
rect 7113 47209 7147 47243
rect 7147 47209 7156 47243
rect 7104 47200 7156 47209
rect 7748 47243 7800 47252
rect 7748 47209 7757 47243
rect 7757 47209 7791 47243
rect 7791 47209 7800 47243
rect 7748 47200 7800 47209
rect 8392 47243 8444 47252
rect 8392 47209 8401 47243
rect 8401 47209 8435 47243
rect 8435 47209 8444 47243
rect 8392 47200 8444 47209
rect 9128 47243 9180 47252
rect 9128 47209 9137 47243
rect 9137 47209 9171 47243
rect 9171 47209 9180 47243
rect 9128 47200 9180 47209
rect 10232 47243 10284 47252
rect 10232 47209 10241 47243
rect 10241 47209 10275 47243
rect 10275 47209 10284 47243
rect 10232 47200 10284 47209
rect 11152 47243 11204 47252
rect 11152 47209 11161 47243
rect 11161 47209 11195 47243
rect 11195 47209 11204 47243
rect 11152 47200 11204 47209
rect 12440 47243 12492 47252
rect 12440 47209 12449 47243
rect 12449 47209 12483 47243
rect 12483 47209 12492 47243
rect 13544 47243 13596 47252
rect 12440 47200 12492 47209
rect 13544 47209 13553 47243
rect 13553 47209 13587 47243
rect 13587 47209 13596 47243
rect 13544 47200 13596 47209
rect 14648 47243 14700 47252
rect 14648 47209 14657 47243
rect 14657 47209 14691 47243
rect 14691 47209 14700 47243
rect 14648 47200 14700 47209
rect 15660 47243 15712 47252
rect 15660 47209 15669 47243
rect 15669 47209 15703 47243
rect 15703 47209 15712 47243
rect 15660 47200 15712 47209
rect 16856 47200 16908 47252
rect 18880 47243 18932 47252
rect 18880 47209 18889 47243
rect 18889 47209 18923 47243
rect 18923 47209 18932 47243
rect 18880 47200 18932 47209
rect 21272 47200 21324 47252
rect 19432 47132 19484 47184
rect 20536 47132 20588 47184
rect 20168 47064 20220 47116
rect 17868 46996 17920 47048
rect 20352 46996 20404 47048
rect 23112 47132 23164 47184
rect 23848 47107 23900 47116
rect 23848 47073 23857 47107
rect 23857 47073 23891 47107
rect 23891 47073 23900 47107
rect 23848 47064 23900 47073
rect 19340 46928 19392 46980
rect 20168 46928 20220 46980
rect 22192 46996 22244 47048
rect 22468 47039 22520 47048
rect 22468 47005 22477 47039
rect 22477 47005 22511 47039
rect 22511 47005 22520 47039
rect 22468 46996 22520 47005
rect 22744 46996 22796 47048
rect 24032 47132 24084 47184
rect 25964 47175 26016 47184
rect 23204 46928 23256 46980
rect 23388 46971 23440 46980
rect 23388 46937 23397 46971
rect 23397 46937 23431 46971
rect 23431 46937 23440 46971
rect 23388 46928 23440 46937
rect 16948 46903 17000 46912
rect 16948 46869 16957 46903
rect 16957 46869 16991 46903
rect 16991 46869 17000 46903
rect 16948 46860 17000 46869
rect 19892 46903 19944 46912
rect 19892 46869 19901 46903
rect 19901 46869 19935 46903
rect 19935 46869 19944 46903
rect 19892 46860 19944 46869
rect 19984 46860 20036 46912
rect 20444 46860 20496 46912
rect 22284 46860 22336 46912
rect 24124 46996 24176 47048
rect 25504 47064 25556 47116
rect 25228 46996 25280 47048
rect 25964 47141 25973 47175
rect 25973 47141 26007 47175
rect 26007 47141 26016 47175
rect 25964 47132 26016 47141
rect 26240 47200 26292 47252
rect 30840 47200 30892 47252
rect 32680 47200 32732 47252
rect 40684 47200 40736 47252
rect 42800 47200 42852 47252
rect 43352 47200 43404 47252
rect 44824 47200 44876 47252
rect 45836 47243 45888 47252
rect 45836 47209 45845 47243
rect 45845 47209 45879 47243
rect 45879 47209 45888 47243
rect 45836 47200 45888 47209
rect 45928 47200 45980 47252
rect 24676 46971 24728 46980
rect 24676 46937 24685 46971
rect 24685 46937 24719 46971
rect 24719 46937 24728 46971
rect 24676 46928 24728 46937
rect 25596 46971 25648 46980
rect 25596 46937 25605 46971
rect 25605 46937 25639 46971
rect 25639 46937 25648 46971
rect 25596 46928 25648 46937
rect 25872 46996 25924 47048
rect 26148 47064 26200 47116
rect 28356 47132 28408 47184
rect 28724 47132 28776 47184
rect 28816 47132 28868 47184
rect 29920 47132 29972 47184
rect 29092 47064 29144 47116
rect 29736 47064 29788 47116
rect 34612 47132 34664 47184
rect 34704 47132 34756 47184
rect 37096 47132 37148 47184
rect 26424 46996 26476 47048
rect 28172 46996 28224 47048
rect 28448 47039 28500 47048
rect 28448 47005 28457 47039
rect 28457 47005 28491 47039
rect 28491 47005 28500 47039
rect 28448 46996 28500 47005
rect 29368 46996 29420 47048
rect 30564 46996 30616 47048
rect 30748 46971 30800 46980
rect 24216 46860 24268 46912
rect 25964 46860 26016 46912
rect 26240 46860 26292 46912
rect 27712 46860 27764 46912
rect 30748 46937 30757 46971
rect 30757 46937 30791 46971
rect 30791 46937 30800 46971
rect 30748 46928 30800 46937
rect 31024 46996 31076 47048
rect 32404 46928 32456 46980
rect 33600 46996 33652 47048
rect 36544 47064 36596 47116
rect 35164 47039 35216 47048
rect 35164 47005 35173 47039
rect 35173 47005 35207 47039
rect 35207 47005 35216 47039
rect 35164 46996 35216 47005
rect 35256 46996 35308 47048
rect 37280 46996 37332 47048
rect 37740 47039 37792 47048
rect 37740 47005 37749 47039
rect 37749 47005 37783 47039
rect 37783 47005 37792 47039
rect 37740 46996 37792 47005
rect 33232 46928 33284 46980
rect 28540 46860 28592 46912
rect 30288 46860 30340 46912
rect 30380 46860 30432 46912
rect 32588 46903 32640 46912
rect 32588 46869 32597 46903
rect 32597 46869 32631 46903
rect 32631 46869 32640 46903
rect 32588 46860 32640 46869
rect 32772 46860 32824 46912
rect 33324 46860 33376 46912
rect 33600 46903 33652 46912
rect 33600 46869 33609 46903
rect 33609 46869 33643 46903
rect 33643 46869 33652 46903
rect 33600 46860 33652 46869
rect 33876 46860 33928 46912
rect 34060 46928 34112 46980
rect 35440 46971 35492 46980
rect 35440 46937 35449 46971
rect 35449 46937 35483 46971
rect 35483 46937 35492 46971
rect 35440 46928 35492 46937
rect 36084 46928 36136 46980
rect 37648 46928 37700 46980
rect 38568 46996 38620 47048
rect 34428 46860 34480 46912
rect 34704 46860 34756 46912
rect 35532 46860 35584 46912
rect 36544 46860 36596 46912
rect 36636 46860 36688 46912
rect 38568 46860 38620 46912
rect 40224 47064 40276 47116
rect 39120 47039 39172 47048
rect 39120 47005 39129 47039
rect 39129 47005 39163 47039
rect 39163 47005 39172 47039
rect 39120 46996 39172 47005
rect 40132 46996 40184 47048
rect 40684 47039 40736 47048
rect 40684 47005 40693 47039
rect 40693 47005 40727 47039
rect 40727 47005 40736 47039
rect 40684 46996 40736 47005
rect 38752 46928 38804 46980
rect 38936 46860 38988 46912
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 16120 46656 16172 46708
rect 17868 46699 17920 46708
rect 17868 46665 17877 46699
rect 17877 46665 17911 46699
rect 17911 46665 17920 46699
rect 17868 46656 17920 46665
rect 12808 46588 12860 46640
rect 19340 46588 19392 46640
rect 6920 46563 6972 46572
rect 6920 46529 6929 46563
rect 6929 46529 6963 46563
rect 6963 46529 6972 46563
rect 6920 46520 6972 46529
rect 17960 46520 18012 46572
rect 18052 46563 18104 46572
rect 18052 46529 18061 46563
rect 18061 46529 18095 46563
rect 18095 46529 18104 46563
rect 18052 46520 18104 46529
rect 19892 46520 19944 46572
rect 20352 46656 20404 46708
rect 22192 46656 22244 46708
rect 20260 46588 20312 46640
rect 22284 46588 22336 46640
rect 20260 46495 20312 46504
rect 20260 46461 20269 46495
rect 20269 46461 20303 46495
rect 20303 46461 20312 46495
rect 20720 46495 20772 46504
rect 20260 46452 20312 46461
rect 20720 46461 20729 46495
rect 20729 46461 20763 46495
rect 20763 46461 20772 46495
rect 20720 46452 20772 46461
rect 21456 46520 21508 46572
rect 22652 46588 22704 46640
rect 23848 46631 23900 46640
rect 23848 46597 23857 46631
rect 23857 46597 23891 46631
rect 23891 46597 23900 46631
rect 23848 46588 23900 46597
rect 25872 46656 25924 46708
rect 26056 46656 26108 46708
rect 26700 46656 26752 46708
rect 28356 46656 28408 46708
rect 28540 46656 28592 46708
rect 29276 46699 29328 46708
rect 29276 46665 29285 46699
rect 29285 46665 29319 46699
rect 29319 46665 29328 46699
rect 29276 46656 29328 46665
rect 30196 46699 30248 46708
rect 30196 46665 30205 46699
rect 30205 46665 30239 46699
rect 30239 46665 30248 46699
rect 30196 46656 30248 46665
rect 31024 46656 31076 46708
rect 33968 46656 34020 46708
rect 32220 46588 32272 46640
rect 32312 46588 32364 46640
rect 34152 46588 34204 46640
rect 34428 46699 34480 46708
rect 34428 46665 34437 46699
rect 34437 46665 34471 46699
rect 34471 46665 34480 46699
rect 34428 46656 34480 46665
rect 35256 46656 35308 46708
rect 35992 46656 36044 46708
rect 21916 46452 21968 46504
rect 22376 46452 22428 46504
rect 23112 46520 23164 46572
rect 24124 46520 24176 46572
rect 24400 46563 24452 46572
rect 24400 46529 24410 46563
rect 24410 46529 24444 46563
rect 24444 46529 24452 46563
rect 24400 46520 24452 46529
rect 24768 46520 24820 46572
rect 25228 46563 25280 46572
rect 25228 46529 25237 46563
rect 25237 46529 25271 46563
rect 25271 46529 25280 46563
rect 25228 46520 25280 46529
rect 25504 46520 25556 46572
rect 25964 46520 26016 46572
rect 26148 46563 26200 46572
rect 26148 46529 26155 46563
rect 26155 46529 26189 46563
rect 26189 46529 26200 46563
rect 26148 46520 26200 46529
rect 27712 46563 27764 46572
rect 27712 46529 27721 46563
rect 27721 46529 27755 46563
rect 27755 46529 27764 46563
rect 27712 46520 27764 46529
rect 27804 46520 27856 46572
rect 29000 46563 29052 46572
rect 22836 46495 22888 46504
rect 22836 46461 22845 46495
rect 22845 46461 22879 46495
rect 22879 46461 22888 46495
rect 22836 46452 22888 46461
rect 23204 46452 23256 46504
rect 24308 46495 24360 46504
rect 24308 46461 24317 46495
rect 24317 46461 24351 46495
rect 24351 46461 24360 46495
rect 26608 46495 26660 46504
rect 24308 46452 24360 46461
rect 26608 46461 26617 46495
rect 26617 46461 26651 46495
rect 26651 46461 26660 46495
rect 26608 46452 26660 46461
rect 27344 46452 27396 46504
rect 29000 46529 29009 46563
rect 29009 46529 29043 46563
rect 29043 46529 29052 46563
rect 29000 46520 29052 46529
rect 29276 46563 29328 46572
rect 29276 46529 29285 46563
rect 29285 46529 29319 46563
rect 29319 46529 29328 46563
rect 29276 46520 29328 46529
rect 30564 46520 30616 46572
rect 31668 46520 31720 46572
rect 31760 46563 31812 46572
rect 31760 46529 31769 46563
rect 31769 46529 31803 46563
rect 31803 46529 31812 46563
rect 32496 46563 32548 46572
rect 31760 46520 31812 46529
rect 29920 46452 29972 46504
rect 30012 46452 30064 46504
rect 30748 46452 30800 46504
rect 31300 46452 31352 46504
rect 32496 46529 32505 46563
rect 32505 46529 32539 46563
rect 32539 46529 32548 46563
rect 32496 46520 32548 46529
rect 32312 46495 32364 46504
rect 32312 46461 32321 46495
rect 32321 46461 32355 46495
rect 32355 46461 32364 46495
rect 32312 46452 32364 46461
rect 21548 46384 21600 46436
rect 22284 46427 22336 46436
rect 22284 46393 22293 46427
rect 22293 46393 22327 46427
rect 22327 46393 22336 46427
rect 22284 46384 22336 46393
rect 22928 46384 22980 46436
rect 23664 46384 23716 46436
rect 25320 46384 25372 46436
rect 18328 46316 18380 46368
rect 19248 46316 19300 46368
rect 19432 46316 19484 46368
rect 20168 46316 20220 46368
rect 25780 46316 25832 46368
rect 26424 46316 26476 46368
rect 26792 46316 26844 46368
rect 27528 46384 27580 46436
rect 29368 46384 29420 46436
rect 30656 46384 30708 46436
rect 32864 46495 32916 46504
rect 32864 46461 32873 46495
rect 32873 46461 32907 46495
rect 32907 46461 32916 46495
rect 32864 46452 32916 46461
rect 33140 46452 33192 46504
rect 33968 46495 34020 46504
rect 33968 46461 33977 46495
rect 33977 46461 34011 46495
rect 34011 46461 34020 46495
rect 33968 46452 34020 46461
rect 34244 46520 34296 46572
rect 36360 46563 36412 46572
rect 36360 46529 36369 46563
rect 36369 46529 36403 46563
rect 36403 46529 36412 46563
rect 36360 46520 36412 46529
rect 36544 46563 36596 46572
rect 36544 46529 36553 46563
rect 36553 46529 36587 46563
rect 36587 46529 36596 46563
rect 36544 46520 36596 46529
rect 35716 46452 35768 46504
rect 32772 46384 32824 46436
rect 27988 46316 28040 46368
rect 29276 46316 29328 46368
rect 31024 46316 31076 46368
rect 32956 46316 33008 46368
rect 34428 46316 34480 46368
rect 34520 46316 34572 46368
rect 36728 46452 36780 46504
rect 38108 46520 38160 46572
rect 38660 46520 38712 46572
rect 38844 46520 38896 46572
rect 38936 46495 38988 46504
rect 36176 46384 36228 46436
rect 37556 46359 37608 46368
rect 37556 46325 37565 46359
rect 37565 46325 37599 46359
rect 37599 46325 37608 46359
rect 37556 46316 37608 46325
rect 38936 46461 38945 46495
rect 38945 46461 38979 46495
rect 38979 46461 38988 46495
rect 38936 46452 38988 46461
rect 39396 46656 39448 46708
rect 41880 46656 41932 46708
rect 40040 46520 40092 46572
rect 42248 46520 42300 46572
rect 43720 46563 43772 46572
rect 43720 46529 43729 46563
rect 43729 46529 43763 46563
rect 43763 46529 43772 46563
rect 43720 46520 43772 46529
rect 44456 46563 44508 46572
rect 44456 46529 44465 46563
rect 44465 46529 44499 46563
rect 44499 46529 44508 46563
rect 44456 46520 44508 46529
rect 39212 46452 39264 46504
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 16948 46112 17000 46164
rect 17868 46112 17920 46164
rect 18052 46112 18104 46164
rect 19064 46044 19116 46096
rect 19248 46044 19300 46096
rect 20536 46112 20588 46164
rect 22836 46112 22888 46164
rect 25688 46112 25740 46164
rect 27344 46155 27396 46164
rect 27344 46121 27353 46155
rect 27353 46121 27387 46155
rect 27387 46121 27396 46155
rect 27344 46112 27396 46121
rect 28816 46112 28868 46164
rect 30840 46155 30892 46164
rect 30840 46121 30849 46155
rect 30849 46121 30883 46155
rect 30883 46121 30892 46155
rect 30840 46112 30892 46121
rect 32496 46112 32548 46164
rect 19892 46044 19944 46096
rect 11704 45908 11756 45960
rect 19984 45976 20036 46028
rect 22652 46044 22704 46096
rect 25228 46044 25280 46096
rect 26148 46044 26200 46096
rect 27436 46044 27488 46096
rect 27620 46044 27672 46096
rect 19892 45951 19944 45960
rect 17224 45840 17276 45892
rect 19892 45917 19901 45951
rect 19901 45917 19935 45951
rect 19935 45917 19944 45951
rect 19892 45908 19944 45917
rect 20168 45908 20220 45960
rect 21456 45908 21508 45960
rect 22008 45908 22060 45960
rect 22284 45951 22336 45960
rect 22284 45917 22293 45951
rect 22293 45917 22327 45951
rect 22327 45917 22336 45951
rect 22284 45908 22336 45917
rect 26608 45976 26660 46028
rect 27712 45976 27764 46028
rect 28724 46044 28776 46096
rect 22652 45951 22704 45960
rect 20444 45840 20496 45892
rect 21732 45840 21784 45892
rect 21916 45840 21968 45892
rect 22652 45917 22661 45951
rect 22661 45917 22695 45951
rect 22695 45917 22704 45951
rect 22652 45908 22704 45917
rect 22928 45951 22980 45960
rect 22928 45917 22937 45951
rect 22937 45917 22971 45951
rect 22971 45917 22980 45951
rect 22928 45908 22980 45917
rect 23756 45908 23808 45960
rect 20720 45772 20772 45824
rect 20996 45772 21048 45824
rect 24124 45840 24176 45892
rect 24860 45840 24912 45892
rect 23664 45815 23716 45824
rect 23664 45781 23673 45815
rect 23673 45781 23707 45815
rect 23707 45781 23716 45815
rect 23664 45772 23716 45781
rect 24032 45772 24084 45824
rect 24400 45772 24452 45824
rect 25780 45951 25832 45960
rect 25780 45917 25789 45951
rect 25789 45917 25823 45951
rect 25823 45917 25832 45951
rect 26516 45951 26568 45960
rect 25780 45908 25832 45917
rect 26516 45917 26525 45951
rect 26525 45917 26559 45951
rect 26559 45917 26568 45951
rect 26516 45908 26568 45917
rect 26700 45908 26752 45960
rect 26332 45883 26384 45892
rect 26332 45849 26341 45883
rect 26341 45849 26375 45883
rect 26375 45849 26384 45883
rect 26332 45840 26384 45849
rect 27620 45951 27672 45960
rect 27620 45917 27629 45951
rect 27629 45917 27663 45951
rect 27663 45917 27672 45951
rect 28080 45976 28132 46028
rect 31024 46044 31076 46096
rect 31944 46044 31996 46096
rect 27620 45908 27672 45917
rect 26792 45772 26844 45824
rect 27712 45840 27764 45892
rect 28448 45908 28500 45960
rect 28724 45908 28776 45960
rect 29092 45951 29144 45994
rect 29092 45942 29101 45951
rect 29101 45942 29135 45951
rect 29135 45942 29144 45951
rect 29736 45976 29788 46028
rect 32772 46044 32824 46096
rect 33600 46112 33652 46164
rect 34336 46112 34388 46164
rect 36728 46112 36780 46164
rect 37924 46112 37976 46164
rect 38292 46112 38344 46164
rect 39304 46112 39356 46164
rect 41328 46155 41380 46164
rect 41328 46121 41337 46155
rect 41337 46121 41371 46155
rect 41371 46121 41380 46155
rect 41328 46112 41380 46121
rect 41512 46112 41564 46164
rect 43812 46155 43864 46164
rect 43812 46121 43821 46155
rect 43821 46121 43855 46155
rect 43855 46121 43864 46155
rect 43812 46112 43864 46121
rect 37004 46044 37056 46096
rect 40776 46044 40828 46096
rect 28356 45840 28408 45892
rect 29000 45840 29052 45892
rect 30380 45908 30432 45960
rect 30748 45908 30800 45960
rect 32036 45951 32088 45960
rect 32036 45917 32045 45951
rect 32045 45917 32079 45951
rect 32079 45917 32088 45951
rect 32036 45908 32088 45917
rect 30288 45883 30340 45892
rect 30288 45849 30297 45883
rect 30297 45849 30331 45883
rect 30331 45849 30340 45883
rect 30288 45840 30340 45849
rect 30840 45840 30892 45892
rect 31300 45883 31352 45892
rect 31300 45849 31309 45883
rect 31309 45849 31343 45883
rect 31343 45849 31352 45883
rect 31300 45840 31352 45849
rect 28908 45772 28960 45824
rect 29552 45772 29604 45824
rect 30012 45772 30064 45824
rect 31024 45772 31076 45824
rect 31668 45840 31720 45892
rect 31852 45883 31904 45892
rect 31852 45849 31861 45883
rect 31861 45849 31895 45883
rect 31895 45849 31904 45883
rect 31852 45840 31904 45849
rect 31484 45772 31536 45824
rect 37924 46019 37976 46028
rect 37924 45985 37933 46019
rect 37933 45985 37967 46019
rect 37967 45985 37976 46019
rect 37924 45976 37976 45985
rect 38292 45976 38344 46028
rect 33140 45908 33192 45960
rect 33968 45951 34020 45960
rect 33968 45917 33977 45951
rect 33977 45917 34011 45951
rect 34011 45917 34020 45951
rect 33968 45908 34020 45917
rect 34336 45951 34388 45960
rect 34336 45917 34345 45951
rect 34345 45917 34379 45951
rect 34379 45917 34388 45951
rect 34336 45908 34388 45917
rect 34612 45908 34664 45960
rect 34980 45951 35032 45960
rect 34980 45917 34989 45951
rect 34989 45917 35023 45951
rect 35023 45917 35032 45951
rect 34980 45908 35032 45917
rect 35532 45908 35584 45960
rect 33324 45883 33376 45892
rect 33324 45849 33333 45883
rect 33333 45849 33367 45883
rect 33367 45849 33376 45883
rect 33324 45840 33376 45849
rect 34428 45840 34480 45892
rect 35900 45908 35952 45960
rect 36084 45951 36136 45960
rect 36084 45917 36093 45951
rect 36093 45917 36127 45951
rect 36127 45917 36136 45951
rect 36084 45908 36136 45917
rect 36360 45908 36412 45960
rect 36268 45840 36320 45892
rect 32588 45772 32640 45824
rect 32864 45815 32916 45824
rect 32864 45781 32873 45815
rect 32873 45781 32907 45815
rect 32907 45781 32916 45815
rect 32864 45772 32916 45781
rect 33600 45772 33652 45824
rect 37096 45815 37148 45824
rect 37096 45781 37105 45815
rect 37105 45781 37139 45815
rect 37139 45781 37148 45815
rect 37096 45772 37148 45781
rect 38384 45908 38436 45960
rect 38844 45908 38896 45960
rect 39212 45951 39264 45960
rect 39212 45917 39221 45951
rect 39221 45917 39255 45951
rect 39255 45917 39264 45951
rect 39212 45908 39264 45917
rect 38016 45840 38068 45892
rect 39396 45840 39448 45892
rect 38752 45772 38804 45824
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 13912 45568 13964 45620
rect 20812 45611 20864 45620
rect 20812 45577 20821 45611
rect 20821 45577 20855 45611
rect 20855 45577 20864 45611
rect 20812 45568 20864 45577
rect 22652 45568 22704 45620
rect 23296 45568 23348 45620
rect 24860 45611 24912 45620
rect 24860 45577 24869 45611
rect 24869 45577 24903 45611
rect 24903 45577 24912 45611
rect 24860 45568 24912 45577
rect 25964 45568 26016 45620
rect 26056 45568 26108 45620
rect 26332 45568 26384 45620
rect 26516 45568 26568 45620
rect 28724 45568 28776 45620
rect 30932 45568 30984 45620
rect 32312 45568 32364 45620
rect 32956 45568 33008 45620
rect 37096 45568 37148 45620
rect 37924 45568 37976 45620
rect 38200 45568 38252 45620
rect 20996 45500 21048 45552
rect 19432 45432 19484 45484
rect 2780 45228 2832 45280
rect 19800 45364 19852 45416
rect 20536 45364 20588 45416
rect 22008 45364 22060 45416
rect 22468 45407 22520 45416
rect 22468 45373 22477 45407
rect 22477 45373 22511 45407
rect 22511 45373 22520 45407
rect 22468 45364 22520 45373
rect 24216 45500 24268 45552
rect 24768 45543 24820 45552
rect 24768 45509 24777 45543
rect 24777 45509 24811 45543
rect 24811 45509 24820 45543
rect 24768 45500 24820 45509
rect 25596 45500 25648 45552
rect 25872 45500 25924 45552
rect 28172 45500 28224 45552
rect 23480 45432 23532 45484
rect 24032 45432 24084 45484
rect 25412 45432 25464 45484
rect 19340 45296 19392 45348
rect 22560 45296 22612 45348
rect 23664 45296 23716 45348
rect 25320 45296 25372 45348
rect 28448 45475 28500 45484
rect 28448 45441 28457 45475
rect 28457 45441 28491 45475
rect 28491 45441 28500 45475
rect 28448 45432 28500 45441
rect 30012 45500 30064 45552
rect 31300 45500 31352 45552
rect 29920 45432 29972 45484
rect 30288 45432 30340 45484
rect 31852 45432 31904 45484
rect 32036 45432 32088 45484
rect 32312 45475 32364 45484
rect 32312 45441 32321 45475
rect 32321 45441 32355 45475
rect 32355 45441 32364 45475
rect 32312 45432 32364 45441
rect 33324 45500 33376 45552
rect 33600 45543 33652 45552
rect 33600 45509 33609 45543
rect 33609 45509 33643 45543
rect 33643 45509 33652 45543
rect 33600 45500 33652 45509
rect 34060 45543 34112 45552
rect 34060 45509 34069 45543
rect 34069 45509 34103 45543
rect 34103 45509 34112 45543
rect 34060 45500 34112 45509
rect 34244 45500 34296 45552
rect 32588 45475 32640 45484
rect 32588 45441 32597 45475
rect 32597 45441 32631 45475
rect 32631 45441 32640 45475
rect 32588 45432 32640 45441
rect 33140 45432 33192 45484
rect 34336 45432 34388 45484
rect 36268 45432 36320 45484
rect 27988 45364 28040 45416
rect 22008 45228 22060 45280
rect 25504 45228 25556 45280
rect 32864 45364 32916 45416
rect 33692 45364 33744 45416
rect 34520 45364 34572 45416
rect 31760 45296 31812 45348
rect 32956 45296 33008 45348
rect 35808 45296 35860 45348
rect 36544 45475 36596 45484
rect 36544 45441 36553 45475
rect 36553 45441 36587 45475
rect 36587 45441 36596 45475
rect 39212 45500 39264 45552
rect 36544 45432 36596 45441
rect 37648 45475 37700 45484
rect 37648 45441 37657 45475
rect 37657 45441 37691 45475
rect 37691 45441 37700 45475
rect 37648 45432 37700 45441
rect 37924 45432 37976 45484
rect 39028 45475 39080 45484
rect 36452 45407 36504 45416
rect 36452 45373 36461 45407
rect 36461 45373 36495 45407
rect 36495 45373 36504 45407
rect 36452 45364 36504 45373
rect 37280 45364 37332 45416
rect 38016 45364 38068 45416
rect 39028 45441 39037 45475
rect 39037 45441 39071 45475
rect 39071 45441 39080 45475
rect 39028 45432 39080 45441
rect 37648 45296 37700 45348
rect 39764 45364 39816 45416
rect 43812 45568 43864 45620
rect 38936 45296 38988 45348
rect 39948 45296 40000 45348
rect 33416 45271 33468 45280
rect 33416 45237 33425 45271
rect 33425 45237 33459 45271
rect 33459 45237 33468 45271
rect 33416 45228 33468 45237
rect 34612 45228 34664 45280
rect 34796 45228 34848 45280
rect 35992 45271 36044 45280
rect 35992 45237 36001 45271
rect 36001 45237 36035 45271
rect 36035 45237 36044 45271
rect 35992 45228 36044 45237
rect 41972 45271 42024 45280
rect 41972 45237 41981 45271
rect 41981 45237 42015 45271
rect 42015 45237 42024 45271
rect 41972 45228 42024 45237
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 17960 45024 18012 45076
rect 20168 45024 20220 45076
rect 22560 45024 22612 45076
rect 24768 45024 24820 45076
rect 27160 45067 27212 45076
rect 27160 45033 27169 45067
rect 27169 45033 27203 45067
rect 27203 45033 27212 45067
rect 27160 45024 27212 45033
rect 23572 44999 23624 45008
rect 23572 44965 23581 44999
rect 23581 44965 23615 44999
rect 23615 44965 23624 44999
rect 23572 44956 23624 44965
rect 23664 44956 23716 45008
rect 19800 44863 19852 44872
rect 19800 44829 19809 44863
rect 19809 44829 19843 44863
rect 19843 44829 19852 44863
rect 19800 44820 19852 44829
rect 19984 44820 20036 44872
rect 20812 44888 20864 44940
rect 27988 45024 28040 45076
rect 28172 45024 28224 45076
rect 29552 45024 29604 45076
rect 32312 45024 32364 45076
rect 34152 45067 34204 45076
rect 34152 45033 34161 45067
rect 34161 45033 34195 45067
rect 34195 45033 34204 45067
rect 34152 45024 34204 45033
rect 35716 45024 35768 45076
rect 22008 44863 22060 44872
rect 22008 44829 22017 44863
rect 22017 44829 22051 44863
rect 22051 44829 22060 44863
rect 22008 44820 22060 44829
rect 24400 44820 24452 44872
rect 24584 44863 24636 44872
rect 24584 44829 24593 44863
rect 24593 44829 24627 44863
rect 24627 44829 24636 44863
rect 24584 44820 24636 44829
rect 24676 44863 24728 44872
rect 24676 44829 24685 44863
rect 24685 44829 24719 44863
rect 24719 44829 24728 44863
rect 24676 44820 24728 44829
rect 20168 44684 20220 44736
rect 20444 44684 20496 44736
rect 20812 44684 20864 44736
rect 22744 44727 22796 44736
rect 22744 44693 22753 44727
rect 22753 44693 22787 44727
rect 22787 44693 22796 44727
rect 22744 44684 22796 44693
rect 23388 44727 23440 44736
rect 23388 44693 23397 44727
rect 23397 44693 23431 44727
rect 23431 44693 23440 44727
rect 23388 44684 23440 44693
rect 24768 44752 24820 44804
rect 25320 44820 25372 44872
rect 25964 44820 26016 44872
rect 27344 44820 27396 44872
rect 29092 44956 29144 45008
rect 27988 44888 28040 44940
rect 33416 44956 33468 45008
rect 27712 44863 27764 44872
rect 27712 44829 27721 44863
rect 27721 44829 27755 44863
rect 27755 44829 27764 44863
rect 28080 44863 28132 44872
rect 27712 44820 27764 44829
rect 28080 44829 28088 44863
rect 28088 44829 28122 44863
rect 28122 44829 28132 44863
rect 28080 44820 28132 44829
rect 26424 44752 26476 44804
rect 27436 44752 27488 44804
rect 29920 44863 29972 44872
rect 29920 44829 29929 44863
rect 29929 44829 29963 44863
rect 29963 44829 29972 44863
rect 29920 44820 29972 44829
rect 30196 44863 30248 44872
rect 30196 44829 30205 44863
rect 30205 44829 30239 44863
rect 30239 44829 30248 44863
rect 30196 44820 30248 44829
rect 31300 44820 31352 44872
rect 32496 44888 32548 44940
rect 32680 44863 32732 44872
rect 32680 44829 32689 44863
rect 32689 44829 32723 44863
rect 32723 44829 32732 44863
rect 32680 44820 32732 44829
rect 33968 44888 34020 44940
rect 34336 44820 34388 44872
rect 28540 44752 28592 44804
rect 29368 44752 29420 44804
rect 24308 44684 24360 44736
rect 26608 44684 26660 44736
rect 35808 44820 35860 44872
rect 36452 44956 36504 45008
rect 36360 44931 36412 44940
rect 36360 44897 36369 44931
rect 36369 44897 36403 44931
rect 36403 44897 36412 44931
rect 36360 44888 36412 44897
rect 37832 45024 37884 45076
rect 39764 45024 39816 45076
rect 41236 45024 41288 45076
rect 44180 45024 44232 45076
rect 40224 44956 40276 45008
rect 37556 44931 37608 44940
rect 37556 44897 37565 44931
rect 37565 44897 37599 44931
rect 37599 44897 37608 44931
rect 37556 44888 37608 44897
rect 37648 44888 37700 44940
rect 41972 44888 42024 44940
rect 36544 44820 36596 44872
rect 37464 44863 37516 44872
rect 37464 44829 37473 44863
rect 37473 44829 37507 44863
rect 37507 44829 37516 44863
rect 37464 44820 37516 44829
rect 37924 44820 37976 44872
rect 35440 44752 35492 44804
rect 38108 44684 38160 44736
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 19984 44480 20036 44532
rect 20536 44480 20588 44532
rect 23204 44523 23256 44532
rect 23204 44489 23213 44523
rect 23213 44489 23247 44523
rect 23247 44489 23256 44523
rect 23204 44480 23256 44489
rect 25412 44523 25464 44532
rect 25412 44489 25421 44523
rect 25421 44489 25455 44523
rect 25455 44489 25464 44523
rect 25412 44480 25464 44489
rect 25504 44480 25556 44532
rect 22376 44412 22428 44464
rect 26148 44412 26200 44464
rect 20812 44387 20864 44396
rect 20812 44353 20821 44387
rect 20821 44353 20855 44387
rect 20855 44353 20864 44387
rect 20812 44344 20864 44353
rect 23388 44344 23440 44396
rect 23940 44387 23992 44396
rect 23940 44353 23949 44387
rect 23949 44353 23983 44387
rect 23983 44353 23992 44387
rect 23940 44344 23992 44353
rect 24860 44344 24912 44396
rect 25872 44344 25924 44396
rect 26424 44344 26476 44396
rect 25320 44276 25372 44328
rect 24492 44208 24544 44260
rect 26608 44387 26660 44396
rect 26608 44353 26617 44387
rect 26617 44353 26651 44387
rect 26651 44353 26660 44387
rect 28080 44412 28132 44464
rect 28172 44455 28224 44464
rect 28172 44421 28181 44455
rect 28181 44421 28215 44455
rect 28215 44421 28224 44455
rect 28172 44412 28224 44421
rect 26608 44344 26660 44353
rect 27712 44387 27764 44396
rect 27712 44353 27721 44387
rect 27721 44353 27755 44387
rect 27755 44353 27764 44387
rect 30380 44480 30432 44532
rect 30932 44480 30984 44532
rect 33324 44480 33376 44532
rect 36360 44480 36412 44532
rect 37556 44523 37608 44532
rect 37556 44489 37565 44523
rect 37565 44489 37599 44523
rect 37599 44489 37608 44523
rect 37556 44480 37608 44489
rect 37740 44480 37792 44532
rect 38108 44480 38160 44532
rect 39028 44480 39080 44532
rect 41236 44480 41288 44532
rect 30656 44412 30708 44464
rect 33140 44412 33192 44464
rect 35440 44412 35492 44464
rect 35992 44412 36044 44464
rect 27712 44344 27764 44353
rect 29644 44387 29696 44396
rect 27344 44276 27396 44328
rect 29644 44353 29653 44387
rect 29653 44353 29687 44387
rect 29687 44353 29696 44387
rect 29644 44344 29696 44353
rect 32956 44344 33008 44396
rect 34612 44387 34664 44396
rect 29092 44276 29144 44328
rect 30104 44276 30156 44328
rect 32220 44276 32272 44328
rect 33232 44276 33284 44328
rect 34612 44353 34621 44387
rect 34621 44353 34655 44387
rect 34655 44353 34664 44387
rect 34612 44344 34664 44353
rect 34796 44387 34848 44396
rect 34796 44353 34805 44387
rect 34805 44353 34839 44387
rect 34839 44353 34848 44387
rect 34796 44344 34848 44353
rect 36176 44344 36228 44396
rect 36912 44412 36964 44464
rect 40224 44455 40276 44464
rect 36544 44344 36596 44396
rect 38016 44387 38068 44396
rect 38016 44353 38025 44387
rect 38025 44353 38059 44387
rect 38059 44353 38068 44387
rect 40224 44421 40233 44455
rect 40233 44421 40267 44455
rect 40267 44421 40276 44455
rect 40224 44412 40276 44421
rect 38016 44344 38068 44353
rect 35348 44276 35400 44328
rect 37648 44276 37700 44328
rect 28080 44208 28132 44260
rect 35440 44140 35492 44192
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 22376 43979 22428 43988
rect 22376 43945 22385 43979
rect 22385 43945 22419 43979
rect 22419 43945 22428 43979
rect 22376 43936 22428 43945
rect 24216 43936 24268 43988
rect 28080 43979 28132 43988
rect 28080 43945 28089 43979
rect 28089 43945 28123 43979
rect 28123 43945 28132 43979
rect 28080 43936 28132 43945
rect 29184 43979 29236 43988
rect 29184 43945 29193 43979
rect 29193 43945 29227 43979
rect 29227 43945 29236 43979
rect 29184 43936 29236 43945
rect 29644 43936 29696 43988
rect 30196 43936 30248 43988
rect 31392 43979 31444 43988
rect 31392 43945 31401 43979
rect 31401 43945 31435 43979
rect 31435 43945 31444 43979
rect 31392 43936 31444 43945
rect 32588 43936 32640 43988
rect 33692 43979 33744 43988
rect 33692 43945 33701 43979
rect 33701 43945 33735 43979
rect 33735 43945 33744 43979
rect 33692 43936 33744 43945
rect 34796 43936 34848 43988
rect 35348 43979 35400 43988
rect 35348 43945 35357 43979
rect 35357 43945 35391 43979
rect 35391 43945 35400 43979
rect 35348 43936 35400 43945
rect 36360 43936 36412 43988
rect 36912 43979 36964 43988
rect 36912 43945 36921 43979
rect 36921 43945 36955 43979
rect 36955 43945 36964 43979
rect 36912 43936 36964 43945
rect 37648 43936 37700 43988
rect 39948 43936 40000 43988
rect 23940 43911 23992 43920
rect 23940 43877 23949 43911
rect 23949 43877 23983 43911
rect 23983 43877 23992 43911
rect 23940 43868 23992 43877
rect 24584 43800 24636 43852
rect 26700 43868 26752 43920
rect 25872 43843 25924 43852
rect 25872 43809 25881 43843
rect 25881 43809 25915 43843
rect 25915 43809 25924 43843
rect 25872 43800 25924 43809
rect 26608 43843 26660 43852
rect 26608 43809 26617 43843
rect 26617 43809 26651 43843
rect 26651 43809 26660 43843
rect 26608 43800 26660 43809
rect 27528 43843 27580 43852
rect 27528 43809 27537 43843
rect 27537 43809 27571 43843
rect 27571 43809 27580 43843
rect 27528 43800 27580 43809
rect 20720 43707 20772 43716
rect 20720 43673 20729 43707
rect 20729 43673 20763 43707
rect 20763 43673 20772 43707
rect 20720 43664 20772 43673
rect 24768 43732 24820 43784
rect 25504 43732 25556 43784
rect 27252 43732 27304 43784
rect 29368 43868 29420 43920
rect 34704 43868 34756 43920
rect 38016 43911 38068 43920
rect 38016 43877 38025 43911
rect 38025 43877 38059 43911
rect 38059 43877 38068 43911
rect 38016 43868 38068 43877
rect 29092 43800 29144 43852
rect 33232 43800 33284 43852
rect 36636 43800 36688 43852
rect 28540 43775 28592 43784
rect 28540 43741 28549 43775
rect 28549 43741 28583 43775
rect 28583 43741 28592 43775
rect 28540 43732 28592 43741
rect 29736 43732 29788 43784
rect 30288 43775 30340 43784
rect 30288 43741 30297 43775
rect 30297 43741 30331 43775
rect 30331 43741 30340 43775
rect 30288 43732 30340 43741
rect 31484 43732 31536 43784
rect 32496 43732 32548 43784
rect 33140 43732 33192 43784
rect 33968 43732 34020 43784
rect 35440 43775 35492 43784
rect 35440 43741 35449 43775
rect 35449 43741 35483 43775
rect 35483 43741 35492 43775
rect 35440 43732 35492 43741
rect 35992 43732 36044 43784
rect 25320 43664 25372 43716
rect 28172 43664 28224 43716
rect 32680 43664 32732 43716
rect 36544 43664 36596 43716
rect 36912 43664 36964 43716
rect 20444 43596 20496 43648
rect 22468 43596 22520 43648
rect 22836 43596 22888 43648
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 22836 43435 22888 43444
rect 22836 43401 22845 43435
rect 22845 43401 22879 43435
rect 22879 43401 22888 43435
rect 22836 43392 22888 43401
rect 24584 43435 24636 43444
rect 24584 43401 24593 43435
rect 24593 43401 24627 43435
rect 24627 43401 24636 43435
rect 24584 43392 24636 43401
rect 24952 43324 25004 43376
rect 25504 43324 25556 43376
rect 25044 43256 25096 43308
rect 20720 43188 20772 43240
rect 24124 43188 24176 43240
rect 24860 43188 24912 43240
rect 26700 43392 26752 43444
rect 27252 43435 27304 43444
rect 27252 43401 27261 43435
rect 27261 43401 27295 43435
rect 27295 43401 27304 43435
rect 27252 43392 27304 43401
rect 27712 43392 27764 43444
rect 28908 43392 28960 43444
rect 30288 43392 30340 43444
rect 30380 43392 30432 43444
rect 32680 43392 32732 43444
rect 35532 43392 35584 43444
rect 36544 43435 36596 43444
rect 36544 43401 36553 43435
rect 36553 43401 36587 43435
rect 36587 43401 36596 43435
rect 36544 43392 36596 43401
rect 37648 43392 37700 43444
rect 38016 43392 38068 43444
rect 38660 43392 38712 43444
rect 34520 43367 34572 43376
rect 34520 43333 34529 43367
rect 34529 43333 34563 43367
rect 34563 43333 34572 43367
rect 34520 43324 34572 43333
rect 39948 43324 40000 43376
rect 28080 43256 28132 43308
rect 29920 43256 29972 43308
rect 30472 43299 30524 43308
rect 30472 43265 30481 43299
rect 30481 43265 30515 43299
rect 30515 43265 30524 43299
rect 30472 43256 30524 43265
rect 31576 43299 31628 43308
rect 31576 43265 31585 43299
rect 31585 43265 31619 43299
rect 31619 43265 31628 43299
rect 31576 43256 31628 43265
rect 33784 43299 33836 43308
rect 33784 43265 33793 43299
rect 33793 43265 33827 43299
rect 33827 43265 33836 43299
rect 33784 43256 33836 43265
rect 34612 43256 34664 43308
rect 35532 43256 35584 43308
rect 27896 43188 27948 43240
rect 26240 43052 26292 43104
rect 27436 43095 27488 43104
rect 27436 43061 27445 43095
rect 27445 43061 27479 43095
rect 27479 43061 27488 43095
rect 27436 43052 27488 43061
rect 39672 43095 39724 43104
rect 39672 43061 39681 43095
rect 39681 43061 39715 43095
rect 39715 43061 39724 43095
rect 39672 43052 39724 43061
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 24768 42848 24820 42900
rect 24860 42848 24912 42900
rect 25596 42848 25648 42900
rect 26240 42848 26292 42900
rect 27712 42848 27764 42900
rect 29368 42848 29420 42900
rect 29736 42891 29788 42900
rect 29736 42857 29745 42891
rect 29745 42857 29779 42891
rect 29779 42857 29788 42891
rect 29736 42848 29788 42857
rect 30380 42891 30432 42900
rect 30380 42857 30389 42891
rect 30389 42857 30423 42891
rect 30423 42857 30432 42891
rect 30380 42848 30432 42857
rect 30472 42848 30524 42900
rect 32680 42848 32732 42900
rect 34612 42848 34664 42900
rect 37648 42848 37700 42900
rect 28908 42780 28960 42832
rect 23020 42755 23072 42764
rect 23020 42721 23029 42755
rect 23029 42721 23063 42755
rect 23063 42721 23072 42755
rect 23020 42712 23072 42721
rect 24216 42712 24268 42764
rect 25136 42712 25188 42764
rect 26700 42712 26752 42764
rect 29000 42712 29052 42764
rect 31300 42712 31352 42764
rect 34336 42712 34388 42764
rect 38752 42712 38804 42764
rect 39672 42712 39724 42764
rect 24952 42687 25004 42696
rect 24952 42653 24961 42687
rect 24961 42653 24995 42687
rect 24995 42653 25004 42687
rect 24952 42644 25004 42653
rect 38016 42576 38068 42628
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 24124 42347 24176 42356
rect 24124 42313 24133 42347
rect 24133 42313 24167 42347
rect 24167 42313 24176 42347
rect 24124 42304 24176 42313
rect 25136 42347 25188 42356
rect 25136 42313 25145 42347
rect 25145 42313 25179 42347
rect 25179 42313 25188 42347
rect 25136 42304 25188 42313
rect 25596 42347 25648 42356
rect 25596 42313 25605 42347
rect 25605 42313 25639 42347
rect 25639 42313 25648 42347
rect 25596 42304 25648 42313
rect 26148 42304 26200 42356
rect 29000 42304 29052 42356
rect 29368 42304 29420 42356
rect 29644 42304 29696 42356
rect 30012 42304 30064 42356
rect 33232 42304 33284 42356
rect 34704 42304 34756 42356
rect 37464 42304 37516 42356
rect 30380 42236 30432 42288
rect 30472 42279 30524 42288
rect 30472 42245 30481 42279
rect 30481 42245 30515 42279
rect 30515 42245 30524 42279
rect 30472 42236 30524 42245
rect 34336 42236 34388 42288
rect 27712 42007 27764 42016
rect 27712 41973 27721 42007
rect 27721 41973 27755 42007
rect 27755 41973 27764 42007
rect 27712 41964 27764 41973
rect 30472 41964 30524 42016
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 24216 41760 24268 41812
rect 26240 41803 26292 41812
rect 26240 41769 26249 41803
rect 26249 41769 26283 41803
rect 26283 41769 26292 41803
rect 26240 41760 26292 41769
rect 26700 41760 26752 41812
rect 29736 41803 29788 41812
rect 29736 41769 29745 41803
rect 29745 41769 29779 41803
rect 29779 41769 29788 41803
rect 29736 41760 29788 41769
rect 27712 41692 27764 41744
rect 29368 41692 29420 41744
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 29644 41216 29696 41268
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 22928 6783 22980 6792
rect 22928 6749 22937 6783
rect 22937 6749 22971 6783
rect 22971 6749 22980 6783
rect 22928 6740 22980 6749
rect 20536 6672 20588 6724
rect 27160 6672 27212 6724
rect 23204 6604 23256 6656
rect 24768 6604 24820 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 20536 6443 20588 6452
rect 20536 6409 20545 6443
rect 20545 6409 20579 6443
rect 20579 6409 20588 6443
rect 20536 6400 20588 6409
rect 27160 6443 27212 6452
rect 27160 6409 27169 6443
rect 27169 6409 27203 6443
rect 27203 6409 27212 6443
rect 27160 6400 27212 6409
rect 25044 6332 25096 6384
rect 21088 6264 21140 6316
rect 22928 6307 22980 6316
rect 22928 6273 22937 6307
rect 22937 6273 22971 6307
rect 22971 6273 22980 6307
rect 22928 6264 22980 6273
rect 24032 6196 24084 6248
rect 25872 6239 25924 6248
rect 25872 6205 25881 6239
rect 25881 6205 25915 6239
rect 25915 6205 25924 6239
rect 25872 6196 25924 6205
rect 26608 6196 26660 6248
rect 24768 6128 24820 6180
rect 24952 6171 25004 6180
rect 24952 6137 24961 6171
rect 24961 6137 24995 6171
rect 24995 6137 25004 6171
rect 24952 6128 25004 6137
rect 22560 6060 22612 6112
rect 23112 6060 23164 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 20536 5856 20588 5908
rect 24032 5899 24084 5908
rect 24032 5865 24041 5899
rect 24041 5865 24075 5899
rect 24075 5865 24084 5899
rect 24032 5856 24084 5865
rect 25044 5899 25096 5908
rect 25044 5865 25053 5899
rect 25053 5865 25087 5899
rect 25087 5865 25096 5899
rect 25044 5856 25096 5865
rect 24768 5788 24820 5840
rect 22928 5763 22980 5772
rect 22928 5729 22937 5763
rect 22937 5729 22971 5763
rect 22971 5729 22980 5763
rect 22928 5720 22980 5729
rect 20260 5652 20312 5704
rect 21088 5695 21140 5704
rect 21088 5661 21097 5695
rect 21097 5661 21131 5695
rect 21131 5661 21140 5695
rect 21088 5652 21140 5661
rect 26240 5720 26292 5772
rect 22560 5627 22612 5636
rect 22560 5593 22569 5627
rect 22569 5593 22603 5627
rect 22603 5593 22612 5627
rect 22560 5584 22612 5593
rect 21732 5516 21784 5568
rect 26240 5627 26292 5636
rect 26240 5593 26249 5627
rect 26249 5593 26283 5627
rect 26283 5593 26292 5627
rect 26240 5584 26292 5593
rect 26700 5584 26752 5636
rect 29000 5652 29052 5704
rect 29092 5584 29144 5636
rect 27344 5516 27396 5568
rect 28540 5516 28592 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 20812 5355 20864 5364
rect 20812 5321 20821 5355
rect 20821 5321 20855 5355
rect 20855 5321 20864 5355
rect 20812 5312 20864 5321
rect 21088 5312 21140 5364
rect 23112 5287 23164 5296
rect 23112 5253 23121 5287
rect 23121 5253 23155 5287
rect 23155 5253 23164 5287
rect 23112 5244 23164 5253
rect 24584 5287 24636 5296
rect 24584 5253 24593 5287
rect 24593 5253 24627 5287
rect 24627 5253 24636 5287
rect 24584 5244 24636 5253
rect 27344 5287 27396 5296
rect 27344 5253 27353 5287
rect 27353 5253 27387 5287
rect 27387 5253 27396 5287
rect 27344 5244 27396 5253
rect 28540 5287 28592 5296
rect 28540 5253 28549 5287
rect 28549 5253 28583 5287
rect 28583 5253 28592 5287
rect 28540 5244 28592 5253
rect 29092 5244 29144 5296
rect 20536 5176 20588 5228
rect 25872 5176 25924 5228
rect 26240 5176 26292 5228
rect 29828 5176 29880 5228
rect 25228 5108 25280 5160
rect 27344 5108 27396 5160
rect 28448 5151 28500 5160
rect 28448 5117 28457 5151
rect 28457 5117 28491 5151
rect 28491 5117 28500 5151
rect 28448 5108 28500 5117
rect 29184 5108 29236 5160
rect 27804 5083 27856 5092
rect 19432 5015 19484 5024
rect 19432 4981 19441 5015
rect 19441 4981 19475 5015
rect 19475 4981 19484 5015
rect 19432 4972 19484 4981
rect 20352 4972 20404 5024
rect 23480 4972 23532 5024
rect 27804 5049 27813 5083
rect 27813 5049 27847 5083
rect 27847 5049 27856 5083
rect 27804 5040 27856 5049
rect 29092 4972 29144 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 27344 4811 27396 4820
rect 27344 4777 27353 4811
rect 27353 4777 27387 4811
rect 27387 4777 27396 4811
rect 27344 4768 27396 4777
rect 22192 4743 22244 4752
rect 20260 4675 20312 4684
rect 20260 4641 20269 4675
rect 20269 4641 20303 4675
rect 20303 4641 20312 4675
rect 20260 4632 20312 4641
rect 22192 4709 22201 4743
rect 22201 4709 22235 4743
rect 22235 4709 22244 4743
rect 22192 4700 22244 4709
rect 23572 4675 23624 4684
rect 23572 4641 23581 4675
rect 23581 4641 23615 4675
rect 23615 4641 23624 4675
rect 23572 4632 23624 4641
rect 26056 4675 26108 4684
rect 26056 4641 26065 4675
rect 26065 4641 26099 4675
rect 26099 4641 26108 4675
rect 26056 4632 26108 4641
rect 28816 4675 28868 4684
rect 28816 4641 28825 4675
rect 28825 4641 28859 4675
rect 28859 4641 28868 4675
rect 28816 4632 28868 4641
rect 29000 4632 29052 4684
rect 16948 4607 17000 4616
rect 16948 4573 16957 4607
rect 16957 4573 16991 4607
rect 16991 4573 17000 4607
rect 16948 4564 17000 4573
rect 19984 4564 20036 4616
rect 27160 4564 27212 4616
rect 20352 4539 20404 4548
rect 20352 4505 20361 4539
rect 20361 4505 20395 4539
rect 20395 4505 20404 4539
rect 20352 4496 20404 4505
rect 21088 4496 21140 4548
rect 21732 4539 21784 4548
rect 21732 4505 21741 4539
rect 21741 4505 21775 4539
rect 21775 4505 21784 4539
rect 21732 4496 21784 4505
rect 21916 4496 21968 4548
rect 23204 4539 23256 4548
rect 23204 4505 23213 4539
rect 23213 4505 23247 4539
rect 23247 4505 23256 4539
rect 25688 4539 25740 4548
rect 23204 4496 23256 4505
rect 25688 4505 25697 4539
rect 25697 4505 25731 4539
rect 25731 4505 25740 4539
rect 25688 4496 25740 4505
rect 29000 4539 29052 4548
rect 29000 4505 29009 4539
rect 29009 4505 29043 4539
rect 29043 4505 29052 4539
rect 29000 4496 29052 4505
rect 26700 4471 26752 4480
rect 26700 4437 26709 4471
rect 26709 4437 26743 4471
rect 26743 4437 26752 4471
rect 26700 4428 26752 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 24584 4224 24636 4276
rect 25688 4224 25740 4276
rect 20812 4156 20864 4208
rect 24308 4199 24360 4208
rect 24308 4165 24317 4199
rect 24317 4165 24351 4199
rect 24351 4165 24360 4199
rect 24308 4156 24360 4165
rect 27712 4199 27764 4208
rect 27712 4165 27721 4199
rect 27721 4165 27755 4199
rect 27755 4165 27764 4199
rect 27712 4156 27764 4165
rect 23664 4088 23716 4140
rect 24860 4088 24912 4140
rect 29828 4131 29880 4140
rect 29828 4097 29837 4131
rect 29837 4097 29871 4131
rect 29871 4097 29880 4131
rect 29828 4088 29880 4097
rect 22468 4063 22520 4072
rect 22468 4029 22477 4063
rect 22477 4029 22511 4063
rect 22511 4029 22520 4063
rect 22468 4020 22520 4029
rect 24676 4063 24728 4072
rect 19156 3952 19208 4004
rect 24676 4029 24685 4063
rect 24685 4029 24719 4063
rect 24719 4029 24728 4063
rect 24676 4020 24728 4029
rect 27436 4063 27488 4072
rect 27436 4029 27445 4063
rect 27445 4029 27479 4063
rect 27479 4029 27488 4063
rect 27436 4020 27488 4029
rect 28908 4020 28960 4072
rect 29736 4020 29788 4072
rect 28448 3952 28500 4004
rect 15016 3927 15068 3936
rect 15016 3893 15025 3927
rect 15025 3893 15059 3927
rect 15059 3893 15068 3927
rect 15016 3884 15068 3893
rect 16120 3927 16172 3936
rect 16120 3893 16129 3927
rect 16129 3893 16163 3927
rect 16163 3893 16172 3927
rect 16120 3884 16172 3893
rect 18052 3884 18104 3936
rect 18880 3927 18932 3936
rect 18880 3893 18889 3927
rect 18889 3893 18923 3927
rect 18923 3893 18932 3927
rect 18880 3884 18932 3893
rect 21916 3884 21968 3936
rect 23664 3884 23716 3936
rect 24768 3884 24820 3936
rect 29092 3884 29144 3936
rect 29920 3884 29972 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 20812 3680 20864 3732
rect 25320 3680 25372 3732
rect 27712 3680 27764 3732
rect 28908 3723 28960 3732
rect 28908 3689 28917 3723
rect 28917 3689 28951 3723
rect 28951 3689 28960 3723
rect 28908 3680 28960 3689
rect 29736 3723 29788 3732
rect 29736 3689 29745 3723
rect 29745 3689 29779 3723
rect 29779 3689 29788 3723
rect 29736 3680 29788 3689
rect 17224 3612 17276 3664
rect 20260 3612 20312 3664
rect 24124 3612 24176 3664
rect 15844 3544 15896 3596
rect 18604 3544 18656 3596
rect 18880 3544 18932 3596
rect 21364 3544 21416 3596
rect 27988 3612 28040 3664
rect 29184 3612 29236 3664
rect 32956 3612 33008 3664
rect 36820 3612 36872 3664
rect 25504 3587 25556 3596
rect 25504 3553 25513 3587
rect 25513 3553 25547 3587
rect 25547 3553 25556 3587
rect 25504 3544 25556 3553
rect 28264 3544 28316 3596
rect 30196 3544 30248 3596
rect 34796 3544 34848 3596
rect 4160 3476 4212 3528
rect 5172 3519 5224 3528
rect 5172 3485 5181 3519
rect 5181 3485 5215 3519
rect 5215 3485 5224 3519
rect 5172 3476 5224 3485
rect 6000 3519 6052 3528
rect 6000 3485 6009 3519
rect 6009 3485 6043 3519
rect 6043 3485 6052 3519
rect 6000 3476 6052 3485
rect 6828 3519 6880 3528
rect 6828 3485 6837 3519
rect 6837 3485 6871 3519
rect 6871 3485 6880 3519
rect 6828 3476 6880 3485
rect 7656 3519 7708 3528
rect 7656 3485 7665 3519
rect 7665 3485 7699 3519
rect 7699 3485 7708 3519
rect 7656 3476 7708 3485
rect 8484 3519 8536 3528
rect 8484 3485 8493 3519
rect 8493 3485 8527 3519
rect 8527 3485 8536 3519
rect 8484 3476 8536 3485
rect 9312 3519 9364 3528
rect 9312 3485 9321 3519
rect 9321 3485 9355 3519
rect 9355 3485 9364 3519
rect 9312 3476 9364 3485
rect 10140 3519 10192 3528
rect 10140 3485 10149 3519
rect 10149 3485 10183 3519
rect 10183 3485 10192 3519
rect 10140 3476 10192 3485
rect 10968 3519 11020 3528
rect 10968 3485 10977 3519
rect 10977 3485 11011 3519
rect 11011 3485 11020 3519
rect 10968 3476 11020 3485
rect 11796 3476 11848 3528
rect 12532 3476 12584 3528
rect 13084 3476 13136 3528
rect 13636 3519 13688 3528
rect 13636 3485 13645 3519
rect 13645 3485 13679 3519
rect 13679 3485 13688 3519
rect 13636 3476 13688 3485
rect 16396 3476 16448 3528
rect 19248 3476 19300 3528
rect 20720 3476 20772 3528
rect 23664 3476 23716 3528
rect 26700 3476 26752 3528
rect 23020 3340 23072 3392
rect 25044 3340 25096 3392
rect 25320 3451 25372 3460
rect 25320 3417 25338 3451
rect 25338 3417 25372 3451
rect 25320 3408 25372 3417
rect 28356 3451 28408 3460
rect 28356 3417 28365 3451
rect 28365 3417 28399 3451
rect 28399 3417 28408 3451
rect 28356 3408 28408 3417
rect 30288 3476 30340 3528
rect 29828 3408 29880 3460
rect 31116 3476 31168 3528
rect 31852 3476 31904 3528
rect 32404 3476 32456 3528
rect 34336 3476 34388 3528
rect 35716 3476 35768 3528
rect 36268 3476 36320 3528
rect 37648 3476 37700 3528
rect 38200 3476 38252 3528
rect 39580 3476 39632 3528
rect 40408 3476 40460 3528
rect 40960 3476 41012 3528
rect 41512 3476 41564 3528
rect 42892 3519 42944 3528
rect 42892 3485 42901 3519
rect 42901 3485 42935 3519
rect 42935 3485 42944 3519
rect 42892 3476 42944 3485
rect 43168 3476 43220 3528
rect 44824 3476 44876 3528
rect 45652 3476 45704 3528
rect 46480 3519 46532 3528
rect 46480 3485 46489 3519
rect 46489 3485 46523 3519
rect 46523 3485 46532 3519
rect 46480 3476 46532 3485
rect 46756 3476 46808 3528
rect 47308 3476 47360 3528
rect 30932 3408 30984 3460
rect 28908 3340 28960 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 16672 3000 16724 3052
rect 20076 3136 20128 3188
rect 23020 3111 23072 3120
rect 23020 3077 23029 3111
rect 23029 3077 23063 3111
rect 23063 3077 23072 3111
rect 23020 3068 23072 3077
rect 24124 3111 24176 3120
rect 24124 3077 24133 3111
rect 24133 3077 24167 3111
rect 24167 3077 24176 3111
rect 24124 3068 24176 3077
rect 25044 3136 25096 3188
rect 18420 3000 18472 3052
rect 19248 3000 19300 3052
rect 20168 3000 20220 3052
rect 20628 3000 20680 3052
rect 5448 2932 5500 2984
rect 7932 2932 7984 2984
rect 9864 2932 9916 2984
rect 4896 2864 4948 2916
rect 6276 2864 6328 2916
rect 3148 2796 3200 2848
rect 3884 2796 3936 2848
rect 6552 2796 6604 2848
rect 8760 2864 8812 2916
rect 11244 2864 11296 2916
rect 13360 2864 13412 2916
rect 14464 2864 14516 2916
rect 17500 2864 17552 2916
rect 21640 2932 21692 2984
rect 18788 2864 18840 2916
rect 22008 2864 22060 2916
rect 9036 2796 9088 2848
rect 10692 2796 10744 2848
rect 12072 2796 12124 2848
rect 13912 2796 13964 2848
rect 15292 2796 15344 2848
rect 15384 2796 15436 2848
rect 17776 2796 17828 2848
rect 18972 2839 19024 2848
rect 18972 2805 18981 2839
rect 18981 2805 19015 2839
rect 19015 2805 19024 2839
rect 18972 2796 19024 2805
rect 20076 2796 20128 2848
rect 20536 2796 20588 2848
rect 20628 2796 20680 2848
rect 22376 2932 22428 2984
rect 23848 2932 23900 2984
rect 24400 2975 24452 2984
rect 24400 2941 24409 2975
rect 24409 2941 24443 2975
rect 24443 2941 24452 2975
rect 24400 2932 24452 2941
rect 28908 3111 28960 3120
rect 28908 3077 28917 3111
rect 28917 3077 28951 3111
rect 28951 3077 28960 3111
rect 28908 3068 28960 3077
rect 31024 3136 31076 3188
rect 30932 3000 30984 3052
rect 32680 3000 32732 3052
rect 25780 2975 25832 2984
rect 25780 2941 25789 2975
rect 25789 2941 25823 2975
rect 25823 2941 25832 2975
rect 25780 2932 25832 2941
rect 27252 2975 27304 2984
rect 23664 2796 23716 2848
rect 27252 2941 27261 2975
rect 27261 2941 27295 2975
rect 27295 2941 27304 2975
rect 27252 2932 27304 2941
rect 28540 2975 28592 2984
rect 26884 2864 26936 2916
rect 28540 2941 28549 2975
rect 28549 2941 28583 2975
rect 28583 2941 28592 2975
rect 28540 2932 28592 2941
rect 29368 2932 29420 2984
rect 31668 2932 31720 2984
rect 32128 2932 32180 2984
rect 34060 2932 34112 2984
rect 37096 2932 37148 2984
rect 38752 2932 38804 2984
rect 40684 2932 40736 2984
rect 42616 2932 42668 2984
rect 44548 2932 44600 2984
rect 28356 2864 28408 2916
rect 30840 2864 30892 2916
rect 31576 2864 31628 2916
rect 33508 2864 33560 2916
rect 35348 2864 35400 2916
rect 37924 2864 37976 2916
rect 29736 2796 29788 2848
rect 35992 2796 36044 2848
rect 39028 2796 39080 2848
rect 40132 2796 40184 2848
rect 42064 2796 42116 2848
rect 43444 2796 43496 2848
rect 43996 2796 44048 2848
rect 45376 2796 45428 2848
rect 45928 2796 45980 2848
rect 47032 2796 47084 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 15384 2592 15436 2644
rect 7104 2524 7156 2576
rect 9588 2524 9640 2576
rect 11520 2524 11572 2576
rect 14188 2524 14240 2576
rect 18328 2524 18380 2576
rect 3516 2456 3568 2508
rect 8208 2456 8260 2508
rect 10416 2456 10468 2508
rect 12808 2456 12860 2508
rect 14740 2456 14792 2508
rect 22284 2456 22336 2508
rect 22744 2499 22796 2508
rect 22744 2465 22753 2499
rect 22753 2465 22787 2499
rect 22787 2465 22796 2499
rect 22744 2456 22796 2465
rect 2596 2388 2648 2440
rect 4620 2388 4672 2440
rect 5724 2388 5776 2440
rect 12256 2388 12308 2440
rect 15568 2388 15620 2440
rect 16304 2431 16356 2440
rect 16304 2397 16313 2431
rect 16313 2397 16347 2431
rect 16347 2397 16356 2431
rect 16304 2388 16356 2397
rect 18420 2388 18472 2440
rect 18880 2431 18932 2440
rect 18880 2397 18889 2431
rect 18889 2397 18923 2431
rect 18923 2397 18932 2431
rect 18880 2388 18932 2397
rect 20168 2388 20220 2440
rect 7380 2320 7432 2372
rect 21916 2320 21968 2372
rect 22008 2252 22060 2304
rect 24308 2592 24360 2644
rect 27252 2592 27304 2644
rect 29736 2635 29788 2644
rect 29736 2601 29745 2635
rect 29745 2601 29779 2635
rect 29779 2601 29788 2635
rect 29736 2592 29788 2601
rect 30288 2592 30340 2644
rect 31024 2635 31076 2644
rect 31024 2601 31033 2635
rect 31033 2601 31067 2635
rect 31067 2601 31076 2635
rect 31024 2592 31076 2601
rect 31668 2592 31720 2644
rect 33232 2524 33284 2576
rect 35440 2524 35492 2576
rect 38476 2524 38528 2576
rect 42340 2524 42392 2576
rect 45100 2524 45152 2576
rect 24124 2456 24176 2508
rect 31300 2456 31352 2508
rect 34612 2456 34664 2508
rect 37372 2456 37424 2508
rect 39304 2456 39356 2508
rect 41236 2456 41288 2508
rect 43720 2456 43772 2508
rect 23664 2388 23716 2440
rect 30840 2388 30892 2440
rect 27160 2363 27212 2372
rect 27160 2329 27169 2363
rect 27169 2329 27203 2363
rect 27203 2329 27212 2363
rect 27160 2320 27212 2329
rect 30472 2320 30524 2372
rect 33784 2388 33836 2440
rect 36544 2388 36596 2440
rect 39856 2388 39908 2440
rect 41788 2388 41840 2440
rect 44272 2320 44324 2372
rect 46204 2388 46256 2440
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 18880 2048 18932 2100
rect 22376 2048 22428 2100
rect 16304 1912 16356 1964
rect 19984 1912 20036 1964
<< metal2 >>
rect 3974 49314 4030 50000
rect 2792 49286 4030 49314
rect 2792 45286 2820 49286
rect 3974 49200 4030 49286
rect 4342 49200 4398 50000
rect 4710 49200 4766 50000
rect 5078 49200 5134 50000
rect 5446 49200 5502 50000
rect 5814 49200 5870 50000
rect 6182 49314 6238 50000
rect 6012 49286 6238 49314
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 4724 47258 4752 49200
rect 4712 47252 4764 47258
rect 4712 47194 4764 47200
rect 5092 46481 5120 49200
rect 5828 47258 5856 49200
rect 6012 47258 6040 49286
rect 6182 49200 6238 49286
rect 6550 49200 6606 50000
rect 6918 49200 6974 50000
rect 7286 49314 7342 50000
rect 7116 49286 7342 49314
rect 5816 47252 5868 47258
rect 5816 47194 5868 47200
rect 6000 47252 6052 47258
rect 6000 47194 6052 47200
rect 6932 46578 6960 49200
rect 7116 47258 7144 49286
rect 7286 49200 7342 49286
rect 7654 49200 7710 50000
rect 8022 49314 8078 50000
rect 7760 49286 8078 49314
rect 7760 47258 7788 49286
rect 8022 49200 8078 49286
rect 8390 49200 8446 50000
rect 8758 49200 8814 50000
rect 9126 49200 9182 50000
rect 9494 49200 9550 50000
rect 9862 49200 9918 50000
rect 10230 49200 10286 50000
rect 10598 49200 10654 50000
rect 10966 49200 11022 50000
rect 11334 49314 11390 50000
rect 11164 49286 11390 49314
rect 8404 47258 8432 49200
rect 9140 47258 9168 49200
rect 7104 47252 7156 47258
rect 7104 47194 7156 47200
rect 7748 47252 7800 47258
rect 7748 47194 7800 47200
rect 8392 47252 8444 47258
rect 8392 47194 8444 47200
rect 9128 47252 9180 47258
rect 9128 47194 9180 47200
rect 9508 46617 9536 49200
rect 10244 47258 10272 49200
rect 10232 47252 10284 47258
rect 10232 47194 10284 47200
rect 9494 46608 9550 46617
rect 6920 46572 6972 46578
rect 9494 46543 9550 46552
rect 6920 46514 6972 46520
rect 5078 46472 5134 46481
rect 5078 46407 5134 46416
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 10612 45937 10640 49200
rect 11164 47258 11192 49286
rect 11334 49200 11390 49286
rect 11702 49200 11758 50000
rect 12070 49200 12126 50000
rect 12438 49200 12494 50000
rect 12806 49200 12862 50000
rect 13174 49200 13230 50000
rect 13542 49200 13598 50000
rect 13910 49200 13966 50000
rect 14278 49200 14334 50000
rect 14646 49200 14702 50000
rect 15014 49200 15070 50000
rect 15382 49200 15438 50000
rect 15750 49314 15806 50000
rect 15672 49286 15806 49314
rect 11152 47252 11204 47258
rect 11152 47194 11204 47200
rect 11716 45966 11744 49200
rect 12452 47258 12480 49200
rect 12440 47252 12492 47258
rect 12440 47194 12492 47200
rect 12820 46646 12848 49200
rect 13556 47258 13584 49200
rect 13544 47252 13596 47258
rect 13544 47194 13596 47200
rect 12808 46640 12860 46646
rect 12808 46582 12860 46588
rect 11704 45960 11756 45966
rect 10598 45928 10654 45937
rect 11704 45902 11756 45908
rect 10598 45863 10654 45872
rect 13924 45626 13952 49200
rect 14660 47258 14688 49200
rect 14648 47252 14700 47258
rect 14648 47194 14700 47200
rect 15028 46345 15056 49200
rect 15672 47258 15700 49286
rect 15750 49200 15806 49286
rect 16118 49200 16174 50000
rect 16486 49200 16542 50000
rect 16854 49200 16910 50000
rect 17222 49200 17278 50000
rect 17590 49200 17646 50000
rect 17958 49200 18014 50000
rect 18326 49200 18382 50000
rect 18694 49200 18750 50000
rect 19062 49200 19118 50000
rect 19430 49200 19486 50000
rect 19798 49200 19854 50000
rect 20166 49200 20222 50000
rect 20534 49200 20590 50000
rect 20902 49200 20958 50000
rect 21270 49200 21326 50000
rect 21638 49200 21694 50000
rect 22006 49200 22062 50000
rect 22374 49314 22430 50000
rect 22742 49314 22798 50000
rect 22112 49286 22430 49314
rect 15660 47252 15712 47258
rect 15660 47194 15712 47200
rect 16132 46714 16160 49200
rect 16868 47258 16896 49200
rect 16856 47252 16908 47258
rect 16856 47194 16908 47200
rect 16948 46912 17000 46918
rect 16948 46854 17000 46860
rect 16120 46708 16172 46714
rect 16120 46650 16172 46656
rect 15014 46336 15070 46345
rect 15014 46271 15070 46280
rect 16960 46170 16988 46854
rect 16948 46164 17000 46170
rect 16948 46106 17000 46112
rect 17236 45898 17264 49200
rect 17868 47048 17920 47054
rect 17868 46990 17920 46996
rect 17880 46714 17908 46990
rect 17868 46708 17920 46714
rect 17868 46650 17920 46656
rect 17972 46578 18000 49200
rect 17960 46572 18012 46578
rect 17960 46514 18012 46520
rect 18052 46572 18104 46578
rect 18052 46514 18104 46520
rect 18064 46170 18092 46514
rect 18340 46374 18368 49200
rect 18880 47456 18932 47462
rect 18880 47398 18932 47404
rect 18892 47258 18920 47398
rect 18880 47252 18932 47258
rect 18880 47194 18932 47200
rect 18328 46368 18380 46374
rect 18328 46310 18380 46316
rect 17868 46164 17920 46170
rect 17868 46106 17920 46112
rect 18052 46164 18104 46170
rect 18052 46106 18104 46112
rect 17224 45892 17276 45898
rect 17224 45834 17276 45840
rect 13912 45620 13964 45626
rect 13912 45562 13964 45568
rect 17880 45554 17908 46106
rect 19076 46102 19104 49200
rect 19444 47598 19472 49200
rect 19432 47592 19484 47598
rect 19432 47534 19484 47540
rect 19892 47524 19944 47530
rect 19892 47466 19944 47472
rect 19432 47184 19484 47190
rect 19432 47126 19484 47132
rect 19340 46980 19392 46986
rect 19340 46922 19392 46928
rect 19352 46646 19380 46922
rect 19340 46640 19392 46646
rect 19340 46582 19392 46588
rect 19444 46458 19472 47126
rect 19904 47002 19932 47466
rect 20180 47122 20208 49200
rect 20260 47592 20312 47598
rect 20260 47534 20312 47540
rect 20168 47116 20220 47122
rect 20168 47058 20220 47064
rect 19904 46974 20116 47002
rect 19904 46918 19932 46974
rect 19892 46912 19944 46918
rect 19892 46854 19944 46860
rect 19984 46912 20036 46918
rect 19984 46854 20036 46860
rect 19574 46812 19882 46821
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46747 19882 46756
rect 19892 46572 19944 46578
rect 19892 46514 19944 46520
rect 19352 46430 19472 46458
rect 19248 46368 19300 46374
rect 19248 46310 19300 46316
rect 19260 46102 19288 46310
rect 19064 46096 19116 46102
rect 19064 46038 19116 46044
rect 19248 46096 19300 46102
rect 19248 46038 19300 46044
rect 17880 45526 18000 45554
rect 2780 45280 2832 45286
rect 2780 45222 2832 45228
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 17972 45082 18000 45526
rect 19352 45354 19380 46430
rect 19432 46368 19484 46374
rect 19432 46310 19484 46316
rect 19444 45490 19472 46310
rect 19904 46102 19932 46514
rect 19892 46096 19944 46102
rect 19892 46038 19944 46044
rect 19996 46034 20024 46854
rect 19984 46028 20036 46034
rect 19984 45970 20036 45976
rect 19892 45960 19944 45966
rect 20088 45914 20116 46974
rect 20168 46980 20220 46986
rect 20168 46922 20220 46928
rect 20180 46374 20208 46922
rect 20272 46646 20300 47534
rect 20548 47190 20576 49200
rect 21284 47258 21312 49200
rect 21272 47252 21324 47258
rect 21272 47194 21324 47200
rect 20536 47184 20588 47190
rect 20536 47126 20588 47132
rect 20352 47048 20404 47054
rect 20352 46990 20404 46996
rect 20364 46714 20392 46990
rect 20444 46912 20496 46918
rect 20444 46854 20496 46860
rect 20352 46708 20404 46714
rect 20352 46650 20404 46656
rect 20260 46640 20312 46646
rect 20260 46582 20312 46588
rect 20260 46504 20312 46510
rect 20260 46446 20312 46452
rect 20168 46368 20220 46374
rect 20168 46310 20220 46316
rect 19944 45908 20116 45914
rect 19892 45902 20116 45908
rect 20168 45960 20220 45966
rect 20272 45948 20300 46446
rect 20364 46209 20392 46650
rect 20350 46200 20406 46209
rect 20350 46135 20406 46144
rect 20220 45920 20300 45948
rect 20168 45902 20220 45908
rect 19904 45886 20116 45902
rect 19574 45724 19882 45733
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45659 19882 45668
rect 19432 45484 19484 45490
rect 19432 45426 19484 45432
rect 19800 45416 19852 45422
rect 19800 45358 19852 45364
rect 19340 45348 19392 45354
rect 19340 45290 19392 45296
rect 17960 45076 18012 45082
rect 17960 45018 18012 45024
rect 19812 44878 19840 45358
rect 20180 45082 20208 45902
rect 20456 45898 20484 46854
rect 21652 46730 21680 49200
rect 22112 47598 22140 49286
rect 22374 49200 22430 49286
rect 22572 49286 22798 49314
rect 21916 47592 21968 47598
rect 21916 47534 21968 47540
rect 22100 47592 22152 47598
rect 22100 47534 22152 47540
rect 21560 46702 21680 46730
rect 21456 46572 21508 46578
rect 21456 46514 21508 46520
rect 20720 46504 20772 46510
rect 20720 46446 20772 46452
rect 20536 46164 20588 46170
rect 20536 46106 20588 46112
rect 20444 45892 20496 45898
rect 20444 45834 20496 45840
rect 20548 45422 20576 46106
rect 20732 45830 20760 46446
rect 21468 45966 21496 46514
rect 21560 46442 21588 46702
rect 21928 46510 21956 47534
rect 22192 47048 22244 47054
rect 22192 46990 22244 46996
rect 22468 47048 22520 47054
rect 22468 46990 22520 46996
rect 22204 46714 22232 46990
rect 22284 46912 22336 46918
rect 22284 46854 22336 46860
rect 22192 46708 22244 46714
rect 22192 46650 22244 46656
rect 21916 46504 21968 46510
rect 21916 46446 21968 46452
rect 21548 46436 21600 46442
rect 21548 46378 21600 46384
rect 21456 45960 21508 45966
rect 21456 45902 21508 45908
rect 22008 45960 22060 45966
rect 22008 45902 22060 45908
rect 21732 45892 21784 45898
rect 21916 45892 21968 45898
rect 21784 45852 21916 45880
rect 21732 45834 21784 45840
rect 21916 45834 21968 45840
rect 20720 45824 20772 45830
rect 20720 45766 20772 45772
rect 20996 45824 21048 45830
rect 20996 45766 21048 45772
rect 20812 45620 20864 45626
rect 20812 45562 20864 45568
rect 20536 45416 20588 45422
rect 20536 45358 20588 45364
rect 20168 45076 20220 45082
rect 20168 45018 20220 45024
rect 19800 44872 19852 44878
rect 19800 44814 19852 44820
rect 19984 44872 20036 44878
rect 19984 44814 20036 44820
rect 19574 44636 19882 44645
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44571 19882 44580
rect 19996 44538 20024 44814
rect 20180 44742 20208 45018
rect 20168 44736 20220 44742
rect 20168 44678 20220 44684
rect 20444 44736 20496 44742
rect 20444 44678 20496 44684
rect 19984 44532 20036 44538
rect 19984 44474 20036 44480
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 20456 43654 20484 44678
rect 20548 44538 20576 45358
rect 20824 44946 20852 45562
rect 21008 45558 21036 45766
rect 20996 45552 21048 45558
rect 20996 45494 21048 45500
rect 22020 45422 22048 45902
rect 22204 45801 22232 46650
rect 22296 46646 22324 46854
rect 22284 46640 22336 46646
rect 22284 46582 22336 46588
rect 22376 46504 22428 46510
rect 22282 46472 22338 46481
rect 22480 46481 22508 46990
rect 22376 46446 22428 46452
rect 22466 46472 22522 46481
rect 22282 46407 22284 46416
rect 22336 46407 22338 46416
rect 22284 46378 22336 46384
rect 22284 45960 22336 45966
rect 22282 45928 22284 45937
rect 22388 45948 22416 46446
rect 22466 46407 22522 46416
rect 22336 45928 22416 45948
rect 22338 45920 22416 45928
rect 22282 45863 22338 45872
rect 22190 45792 22246 45801
rect 22190 45727 22246 45736
rect 22480 45422 22508 46407
rect 22008 45416 22060 45422
rect 22008 45358 22060 45364
rect 22468 45416 22520 45422
rect 22468 45358 22520 45364
rect 22008 45280 22060 45286
rect 22008 45222 22060 45228
rect 20812 44940 20864 44946
rect 20812 44882 20864 44888
rect 22020 44878 22048 45222
rect 22008 44872 22060 44878
rect 22008 44814 22060 44820
rect 20812 44736 20864 44742
rect 20812 44678 20864 44684
rect 20536 44532 20588 44538
rect 20536 44474 20588 44480
rect 20824 44402 20852 44678
rect 22376 44464 22428 44470
rect 22376 44406 22428 44412
rect 20812 44396 20864 44402
rect 20812 44338 20864 44344
rect 22388 43994 22416 44406
rect 22376 43988 22428 43994
rect 22376 43930 22428 43936
rect 20720 43716 20772 43722
rect 20720 43658 20772 43664
rect 20444 43648 20496 43654
rect 20444 43590 20496 43596
rect 19574 43548 19882 43557
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43483 19882 43492
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 20456 16574 20484 43590
rect 20732 43246 20760 43658
rect 22480 43654 22508 45358
rect 22572 45354 22600 49286
rect 22742 49200 22798 49286
rect 23110 49200 23166 50000
rect 23478 49200 23534 50000
rect 23846 49200 23902 50000
rect 24214 49200 24270 50000
rect 24582 49200 24638 50000
rect 24950 49200 25006 50000
rect 25318 49200 25374 50000
rect 25686 49200 25742 50000
rect 26054 49200 26110 50000
rect 26422 49314 26478 50000
rect 26422 49286 26740 49314
rect 26422 49200 26478 49286
rect 23492 47462 23520 49200
rect 23480 47456 23532 47462
rect 23480 47398 23532 47404
rect 23112 47184 23164 47190
rect 23112 47126 23164 47132
rect 22744 47048 22796 47054
rect 22744 46990 22796 46996
rect 22650 46744 22706 46753
rect 22650 46679 22706 46688
rect 22664 46646 22692 46679
rect 22652 46640 22704 46646
rect 22652 46582 22704 46588
rect 22652 46096 22704 46102
rect 22652 46038 22704 46044
rect 22664 45966 22692 46038
rect 22652 45960 22704 45966
rect 22652 45902 22704 45908
rect 22664 45626 22692 45902
rect 22652 45620 22704 45626
rect 22652 45562 22704 45568
rect 22560 45348 22612 45354
rect 22560 45290 22612 45296
rect 22572 45082 22600 45290
rect 22560 45076 22612 45082
rect 22560 45018 22612 45024
rect 22756 44742 22784 46990
rect 23018 46744 23074 46753
rect 23018 46679 23074 46688
rect 22926 46608 22982 46617
rect 22926 46543 22982 46552
rect 22836 46504 22888 46510
rect 22836 46446 22888 46452
rect 22848 46170 22876 46446
rect 22940 46442 22968 46543
rect 22928 46436 22980 46442
rect 22928 46378 22980 46384
rect 22836 46164 22888 46170
rect 22836 46106 22888 46112
rect 22926 46064 22982 46073
rect 22926 45999 22982 46008
rect 22940 45966 22968 45999
rect 22928 45960 22980 45966
rect 22928 45902 22980 45908
rect 22744 44736 22796 44742
rect 22744 44678 22796 44684
rect 22468 43648 22520 43654
rect 22468 43590 22520 43596
rect 22836 43648 22888 43654
rect 22836 43590 22888 43596
rect 22848 43450 22876 43590
rect 22836 43444 22888 43450
rect 22836 43386 22888 43392
rect 20720 43240 20772 43246
rect 20720 43182 20772 43188
rect 23032 42770 23060 46679
rect 23124 46578 23152 47126
rect 23860 47122 23888 49200
rect 24124 47456 24176 47462
rect 24124 47398 24176 47404
rect 24032 47184 24084 47190
rect 24032 47126 24084 47132
rect 23848 47116 23900 47122
rect 23848 47058 23900 47064
rect 23204 46980 23256 46986
rect 23204 46922 23256 46928
rect 23388 46980 23440 46986
rect 23388 46922 23440 46928
rect 23112 46572 23164 46578
rect 23112 46514 23164 46520
rect 23216 46510 23244 46922
rect 23204 46504 23256 46510
rect 23204 46446 23256 46452
rect 23216 44538 23244 46446
rect 23400 46345 23428 46922
rect 23860 46646 23888 47058
rect 23848 46640 23900 46646
rect 23848 46582 23900 46588
rect 23664 46436 23716 46442
rect 23664 46378 23716 46384
rect 23386 46336 23442 46345
rect 23386 46271 23442 46280
rect 23294 46200 23350 46209
rect 23294 46135 23350 46144
rect 23308 45626 23336 46135
rect 23676 45830 23704 46378
rect 23756 45960 23808 45966
rect 23756 45902 23808 45908
rect 23664 45824 23716 45830
rect 23664 45766 23716 45772
rect 23296 45620 23348 45626
rect 23296 45562 23348 45568
rect 23480 45484 23532 45490
rect 23676 45472 23704 45766
rect 23532 45444 23704 45472
rect 23480 45426 23532 45432
rect 23584 45014 23612 45444
rect 23664 45348 23716 45354
rect 23768 45336 23796 45902
rect 24044 45830 24072 47126
rect 24136 47054 24164 47398
rect 24124 47048 24176 47054
rect 24124 46990 24176 46996
rect 24228 46918 24256 49200
rect 24216 46912 24268 46918
rect 24216 46854 24268 46860
rect 24124 46572 24176 46578
rect 24124 46514 24176 46520
rect 24136 45898 24164 46514
rect 24124 45892 24176 45898
rect 24124 45834 24176 45840
rect 24032 45824 24084 45830
rect 24032 45766 24084 45772
rect 24044 45490 24072 45766
rect 24228 45558 24256 46854
rect 24400 46572 24452 46578
rect 24400 46514 24452 46520
rect 24308 46504 24360 46510
rect 24308 46446 24360 46452
rect 24320 46345 24348 46446
rect 24306 46336 24362 46345
rect 24306 46271 24362 46280
rect 24216 45552 24268 45558
rect 24216 45494 24268 45500
rect 24032 45484 24084 45490
rect 24032 45426 24084 45432
rect 23716 45308 23796 45336
rect 23664 45290 23716 45296
rect 23676 45014 23704 45290
rect 23572 45008 23624 45014
rect 23572 44950 23624 44956
rect 23664 45008 23716 45014
rect 23664 44950 23716 44956
rect 23388 44736 23440 44742
rect 23388 44678 23440 44684
rect 23204 44532 23256 44538
rect 23204 44474 23256 44480
rect 23400 44402 23428 44678
rect 23388 44396 23440 44402
rect 23388 44338 23440 44344
rect 23940 44396 23992 44402
rect 23940 44338 23992 44344
rect 23952 43926 23980 44338
rect 24228 43994 24256 45494
rect 24320 44742 24348 46271
rect 24412 45830 24440 46514
rect 24400 45824 24452 45830
rect 24400 45766 24452 45772
rect 24412 44878 24440 45766
rect 24596 45472 24624 49200
rect 24676 46980 24728 46986
rect 24676 46922 24728 46928
rect 24504 45444 24624 45472
rect 24400 44872 24452 44878
rect 24400 44814 24452 44820
rect 24308 44736 24360 44742
rect 24308 44678 24360 44684
rect 24504 44266 24532 45444
rect 24688 44878 24716 46922
rect 24768 46572 24820 46578
rect 24768 46514 24820 46520
rect 24780 46481 24808 46514
rect 24766 46472 24822 46481
rect 24766 46407 24822 46416
rect 24860 45892 24912 45898
rect 24860 45834 24912 45840
rect 24872 45665 24900 45834
rect 24858 45656 24914 45665
rect 24858 45591 24860 45600
rect 24912 45591 24914 45600
rect 24860 45562 24912 45568
rect 24768 45552 24820 45558
rect 24768 45494 24820 45500
rect 24780 45082 24808 45494
rect 24768 45076 24820 45082
rect 24768 45018 24820 45024
rect 24584 44872 24636 44878
rect 24584 44814 24636 44820
rect 24676 44872 24728 44878
rect 24676 44814 24728 44820
rect 24492 44260 24544 44266
rect 24492 44202 24544 44208
rect 24216 43988 24268 43994
rect 24216 43930 24268 43936
rect 23940 43920 23992 43926
rect 23940 43862 23992 43868
rect 24124 43240 24176 43246
rect 24124 43182 24176 43188
rect 23020 42764 23072 42770
rect 23020 42706 23072 42712
rect 24136 42362 24164 43182
rect 24228 42770 24256 43930
rect 24596 43858 24624 44814
rect 24768 44804 24820 44810
rect 24768 44746 24820 44752
rect 24584 43852 24636 43858
rect 24584 43794 24636 43800
rect 24596 43450 24624 43794
rect 24780 43790 24808 44746
rect 24872 44402 24900 45562
rect 24860 44396 24912 44402
rect 24860 44338 24912 44344
rect 24768 43784 24820 43790
rect 24768 43726 24820 43732
rect 24584 43444 24636 43450
rect 24584 43386 24636 43392
rect 24780 42906 24808 43726
rect 24872 43246 24900 44338
rect 24964 43874 24992 49200
rect 25228 47048 25280 47054
rect 25228 46990 25280 46996
rect 25240 46578 25268 46990
rect 25228 46572 25280 46578
rect 25228 46514 25280 46520
rect 25240 46102 25268 46514
rect 25332 46442 25360 49200
rect 25504 47116 25556 47122
rect 25504 47058 25556 47064
rect 25516 46578 25544 47058
rect 25596 46980 25648 46986
rect 25596 46922 25648 46928
rect 25504 46572 25556 46578
rect 25504 46514 25556 46520
rect 25320 46436 25372 46442
rect 25320 46378 25372 46384
rect 25228 46096 25280 46102
rect 25228 46038 25280 46044
rect 25412 45484 25464 45490
rect 25412 45426 25464 45432
rect 25320 45348 25372 45354
rect 25320 45290 25372 45296
rect 25332 44878 25360 45290
rect 25320 44872 25372 44878
rect 25320 44814 25372 44820
rect 25332 44334 25360 44814
rect 25424 44538 25452 45426
rect 25516 45286 25544 46514
rect 25608 45558 25636 46922
rect 25700 46170 25728 49200
rect 26068 47580 26096 49200
rect 26068 47552 26280 47580
rect 26252 47258 26280 47552
rect 26240 47252 26292 47258
rect 26240 47194 26292 47200
rect 25964 47184 26016 47190
rect 25964 47126 26016 47132
rect 25872 47048 25924 47054
rect 25872 46990 25924 46996
rect 25884 46714 25912 46990
rect 25976 46918 26004 47126
rect 26148 47116 26200 47122
rect 26148 47058 26200 47064
rect 25964 46912 26016 46918
rect 25964 46854 26016 46860
rect 25976 46730 26004 46854
rect 25976 46714 26096 46730
rect 25872 46708 25924 46714
rect 25976 46708 26108 46714
rect 25976 46702 26056 46708
rect 25872 46650 25924 46656
rect 26056 46650 26108 46656
rect 26160 46578 26188 47058
rect 26424 47048 26476 47054
rect 26424 46990 26476 46996
rect 26240 46912 26292 46918
rect 26240 46854 26292 46860
rect 25964 46572 26016 46578
rect 25964 46514 26016 46520
rect 26148 46572 26200 46578
rect 26148 46514 26200 46520
rect 25780 46368 25832 46374
rect 25780 46310 25832 46316
rect 25688 46164 25740 46170
rect 25688 46106 25740 46112
rect 25792 45966 25820 46310
rect 25780 45960 25832 45966
rect 25780 45902 25832 45908
rect 25976 45626 26004 46514
rect 26252 46186 26280 46854
rect 26436 46374 26464 46990
rect 26712 46714 26740 49286
rect 26790 49200 26846 50000
rect 27158 49200 27214 50000
rect 27526 49200 27582 50000
rect 27894 49200 27950 50000
rect 28262 49200 28318 50000
rect 28630 49314 28686 50000
rect 28368 49286 28686 49314
rect 26804 47598 26832 49200
rect 26792 47592 26844 47598
rect 26792 47534 26844 47540
rect 26700 46708 26752 46714
rect 26700 46650 26752 46656
rect 26608 46504 26660 46510
rect 26608 46446 26660 46452
rect 26424 46368 26476 46374
rect 26424 46310 26476 46316
rect 26068 46158 26280 46186
rect 26068 45665 26096 46158
rect 26148 46096 26200 46102
rect 26148 46038 26200 46044
rect 26054 45656 26110 45665
rect 25964 45620 26016 45626
rect 26054 45591 26056 45600
rect 25964 45562 26016 45568
rect 26108 45591 26110 45600
rect 26056 45562 26108 45568
rect 25596 45552 25648 45558
rect 25596 45494 25648 45500
rect 25872 45552 25924 45558
rect 25872 45494 25924 45500
rect 25504 45280 25556 45286
rect 25504 45222 25556 45228
rect 25412 44532 25464 44538
rect 25412 44474 25464 44480
rect 25504 44532 25556 44538
rect 25504 44474 25556 44480
rect 25320 44328 25372 44334
rect 25320 44270 25372 44276
rect 24964 43846 25084 43874
rect 24952 43376 25004 43382
rect 24952 43318 25004 43324
rect 24860 43240 24912 43246
rect 24860 43182 24912 43188
rect 24872 42906 24900 43182
rect 24768 42900 24820 42906
rect 24768 42842 24820 42848
rect 24860 42900 24912 42906
rect 24860 42842 24912 42848
rect 24216 42764 24268 42770
rect 24216 42706 24268 42712
rect 24124 42356 24176 42362
rect 24124 42298 24176 42304
rect 24228 41818 24256 42706
rect 24964 42702 24992 43318
rect 25056 43314 25084 43846
rect 25332 43722 25360 44270
rect 25516 43790 25544 44474
rect 25884 44402 25912 45494
rect 25976 44878 26004 45562
rect 26068 45531 26096 45562
rect 25964 44872 26016 44878
rect 25964 44814 26016 44820
rect 26160 44470 26188 46038
rect 26620 46034 26648 46446
rect 26608 46028 26660 46034
rect 26608 45970 26660 45976
rect 26712 45966 26740 46650
rect 26792 46368 26844 46374
rect 26792 46310 26844 46316
rect 26516 45960 26568 45966
rect 26516 45902 26568 45908
rect 26700 45960 26752 45966
rect 26700 45902 26752 45908
rect 26332 45892 26384 45898
rect 26332 45834 26384 45840
rect 26344 45626 26372 45834
rect 26528 45626 26556 45902
rect 26332 45620 26384 45626
rect 26332 45562 26384 45568
rect 26516 45620 26568 45626
rect 26516 45562 26568 45568
rect 26424 44804 26476 44810
rect 26424 44746 26476 44752
rect 26148 44464 26200 44470
rect 26148 44406 26200 44412
rect 25872 44396 25924 44402
rect 25872 44338 25924 44344
rect 25884 43858 25912 44338
rect 25872 43852 25924 43858
rect 25872 43794 25924 43800
rect 25504 43784 25556 43790
rect 25504 43726 25556 43732
rect 25320 43716 25372 43722
rect 25320 43658 25372 43664
rect 25516 43382 25544 43726
rect 25504 43376 25556 43382
rect 25504 43318 25556 43324
rect 25044 43308 25096 43314
rect 25044 43250 25096 43256
rect 25596 42900 25648 42906
rect 25596 42842 25648 42848
rect 25136 42764 25188 42770
rect 25136 42706 25188 42712
rect 24952 42696 25004 42702
rect 24952 42638 25004 42644
rect 25148 42362 25176 42706
rect 25608 42362 25636 42842
rect 26160 42362 26188 44406
rect 26436 44402 26464 44746
rect 26608 44736 26660 44742
rect 26608 44678 26660 44684
rect 26620 44402 26648 44678
rect 26424 44396 26476 44402
rect 26424 44338 26476 44344
rect 26608 44396 26660 44402
rect 26608 44338 26660 44344
rect 26620 43858 26648 44338
rect 26712 43926 26740 45902
rect 26804 45830 26832 46310
rect 26792 45824 26844 45830
rect 26792 45766 26844 45772
rect 27172 45082 27200 49200
rect 27540 46560 27568 49200
rect 27712 46912 27764 46918
rect 27712 46854 27764 46860
rect 27724 46578 27752 46854
rect 27448 46532 27568 46560
rect 27712 46572 27764 46578
rect 27344 46504 27396 46510
rect 27344 46446 27396 46452
rect 27356 46170 27384 46446
rect 27344 46164 27396 46170
rect 27344 46106 27396 46112
rect 27448 46102 27476 46532
rect 27712 46514 27764 46520
rect 27804 46572 27856 46578
rect 27804 46514 27856 46520
rect 27528 46436 27580 46442
rect 27528 46378 27580 46384
rect 27436 46096 27488 46102
rect 27436 46038 27488 46044
rect 27160 45076 27212 45082
rect 27160 45018 27212 45024
rect 27344 44872 27396 44878
rect 27344 44814 27396 44820
rect 27356 44334 27384 44814
rect 27436 44804 27488 44810
rect 27436 44746 27488 44752
rect 27344 44328 27396 44334
rect 27344 44270 27396 44276
rect 26700 43920 26752 43926
rect 26700 43862 26752 43868
rect 26608 43852 26660 43858
rect 26608 43794 26660 43800
rect 26712 43450 26740 43862
rect 27252 43784 27304 43790
rect 27252 43726 27304 43732
rect 27264 43450 27292 43726
rect 26700 43444 26752 43450
rect 26700 43386 26752 43392
rect 27252 43444 27304 43450
rect 27252 43386 27304 43392
rect 26240 43104 26292 43110
rect 26240 43046 26292 43052
rect 26252 42906 26280 43046
rect 26240 42900 26292 42906
rect 26240 42842 26292 42848
rect 25136 42356 25188 42362
rect 25136 42298 25188 42304
rect 25596 42356 25648 42362
rect 25596 42298 25648 42304
rect 26148 42356 26200 42362
rect 26148 42298 26200 42304
rect 26252 41818 26280 42842
rect 26712 42770 26740 43386
rect 27448 43110 27476 44746
rect 27540 43858 27568 46378
rect 27710 46200 27766 46209
rect 27710 46135 27766 46144
rect 27620 46096 27672 46102
rect 27620 46038 27672 46044
rect 27632 45966 27660 46038
rect 27724 46034 27752 46135
rect 27712 46028 27764 46034
rect 27712 45970 27764 45976
rect 27620 45960 27672 45966
rect 27620 45902 27672 45908
rect 27712 45892 27764 45898
rect 27816 45880 27844 46514
rect 27764 45852 27844 45880
rect 27712 45834 27764 45840
rect 27712 44872 27764 44878
rect 27712 44814 27764 44820
rect 27724 44402 27752 44814
rect 27712 44396 27764 44402
rect 27712 44338 27764 44344
rect 27528 43852 27580 43858
rect 27528 43794 27580 43800
rect 27724 43450 27752 44338
rect 27712 43444 27764 43450
rect 27712 43386 27764 43392
rect 27436 43104 27488 43110
rect 27436 43046 27488 43052
rect 27724 42906 27752 43386
rect 27908 43246 27936 49200
rect 28172 47048 28224 47054
rect 28172 46990 28224 46996
rect 27988 46368 28040 46374
rect 27988 46310 28040 46316
rect 28000 45422 28028 46310
rect 28080 46028 28132 46034
rect 28080 45970 28132 45976
rect 27988 45416 28040 45422
rect 27988 45358 28040 45364
rect 27988 45076 28040 45082
rect 27988 45018 28040 45024
rect 28000 44946 28028 45018
rect 27988 44940 28040 44946
rect 27988 44882 28040 44888
rect 28092 44878 28120 45970
rect 28184 45558 28212 46990
rect 28276 45665 28304 49200
rect 28368 47190 28396 49286
rect 28630 49200 28686 49286
rect 28998 49200 29054 50000
rect 29366 49314 29422 50000
rect 29196 49286 29422 49314
rect 29012 47666 29040 49200
rect 29000 47660 29052 47666
rect 29000 47602 29052 47608
rect 28816 47592 28868 47598
rect 28816 47534 28868 47540
rect 28828 47190 28856 47534
rect 28356 47184 28408 47190
rect 28356 47126 28408 47132
rect 28724 47184 28776 47190
rect 28724 47126 28776 47132
rect 28816 47184 28868 47190
rect 28816 47126 28868 47132
rect 28448 47048 28500 47054
rect 28448 46990 28500 46996
rect 28356 46708 28408 46714
rect 28356 46650 28408 46656
rect 28368 45898 28396 46650
rect 28460 45966 28488 46990
rect 28540 46912 28592 46918
rect 28540 46854 28592 46860
rect 28552 46714 28580 46854
rect 28540 46708 28592 46714
rect 28540 46650 28592 46656
rect 28736 46102 28764 47126
rect 29092 47116 29144 47122
rect 29092 47058 29144 47064
rect 29000 46572 29052 46578
rect 29000 46514 29052 46520
rect 28814 46336 28870 46345
rect 28814 46271 28870 46280
rect 28828 46170 28856 46271
rect 28906 46200 28962 46209
rect 28816 46164 28868 46170
rect 28906 46135 28962 46144
rect 28816 46106 28868 46112
rect 28724 46096 28776 46102
rect 28724 46038 28776 46044
rect 28448 45960 28500 45966
rect 28448 45902 28500 45908
rect 28724 45960 28776 45966
rect 28920 45948 28948 46135
rect 29012 46073 29040 46514
rect 28998 46064 29054 46073
rect 28998 45999 29054 46008
rect 29104 46000 29132 47058
rect 29092 45994 29144 46000
rect 28920 45920 28994 45948
rect 29092 45936 29144 45942
rect 28724 45902 28776 45908
rect 28966 45914 28994 45920
rect 28356 45892 28408 45898
rect 28356 45834 28408 45840
rect 28262 45656 28318 45665
rect 28262 45591 28318 45600
rect 28172 45552 28224 45558
rect 28172 45494 28224 45500
rect 28460 45490 28488 45902
rect 28736 45626 28764 45902
rect 28966 45898 29040 45914
rect 28966 45892 29052 45898
rect 28966 45886 29000 45892
rect 29000 45834 29052 45840
rect 28908 45824 28960 45830
rect 28908 45766 28960 45772
rect 28920 45665 28948 45766
rect 28906 45656 28962 45665
rect 28724 45620 28776 45626
rect 28906 45591 28962 45600
rect 28724 45562 28776 45568
rect 28448 45484 28500 45490
rect 28448 45426 28500 45432
rect 28172 45076 28224 45082
rect 28172 45018 28224 45024
rect 28080 44872 28132 44878
rect 28080 44814 28132 44820
rect 28092 44470 28120 44814
rect 28184 44470 28212 45018
rect 29104 45014 29132 45936
rect 29092 45008 29144 45014
rect 29092 44950 29144 44956
rect 28540 44804 28592 44810
rect 28540 44746 28592 44752
rect 28080 44464 28132 44470
rect 28080 44406 28132 44412
rect 28172 44464 28224 44470
rect 28172 44406 28224 44412
rect 28080 44260 28132 44266
rect 28080 44202 28132 44208
rect 28092 43994 28120 44202
rect 28080 43988 28132 43994
rect 28080 43930 28132 43936
rect 28092 43314 28120 43930
rect 28184 43722 28212 44406
rect 28552 43790 28580 44746
rect 29104 44334 29132 44950
rect 29092 44328 29144 44334
rect 29092 44270 29144 44276
rect 29104 43858 29132 44270
rect 29196 43994 29224 49286
rect 29366 49200 29422 49286
rect 29734 49200 29790 50000
rect 30102 49200 30158 50000
rect 30470 49314 30526 50000
rect 30470 49286 30696 49314
rect 30470 49200 30526 49286
rect 29748 47122 29776 49200
rect 29920 47184 29972 47190
rect 29920 47126 29972 47132
rect 29736 47116 29788 47122
rect 29736 47058 29788 47064
rect 29368 47048 29420 47054
rect 29368 46990 29420 46996
rect 29274 46744 29330 46753
rect 29274 46679 29276 46688
rect 29328 46679 29330 46688
rect 29276 46650 29328 46656
rect 29276 46572 29328 46578
rect 29276 46514 29328 46520
rect 29288 46374 29316 46514
rect 29380 46442 29408 46990
rect 29368 46436 29420 46442
rect 29368 46378 29420 46384
rect 29276 46368 29328 46374
rect 29276 46310 29328 46316
rect 29380 44810 29408 46378
rect 29748 46034 29776 47058
rect 29932 46510 29960 47126
rect 29920 46504 29972 46510
rect 29920 46446 29972 46452
rect 30012 46504 30064 46510
rect 30012 46446 30064 46452
rect 29736 46028 29788 46034
rect 29736 45970 29788 45976
rect 29552 45824 29604 45830
rect 29552 45766 29604 45772
rect 29564 45082 29592 45766
rect 29552 45076 29604 45082
rect 29552 45018 29604 45024
rect 29368 44804 29420 44810
rect 29368 44746 29420 44752
rect 29184 43988 29236 43994
rect 29184 43930 29236 43936
rect 29380 43926 29408 44746
rect 29644 44396 29696 44402
rect 29644 44338 29696 44344
rect 29656 43994 29684 44338
rect 29644 43988 29696 43994
rect 29644 43930 29696 43936
rect 29368 43920 29420 43926
rect 29368 43862 29420 43868
rect 29092 43852 29144 43858
rect 29092 43794 29144 43800
rect 28540 43784 28592 43790
rect 28540 43726 28592 43732
rect 28172 43716 28224 43722
rect 28172 43658 28224 43664
rect 28908 43444 28960 43450
rect 28908 43386 28960 43392
rect 28080 43308 28132 43314
rect 28080 43250 28132 43256
rect 27896 43240 27948 43246
rect 27896 43182 27948 43188
rect 27712 42900 27764 42906
rect 27712 42842 27764 42848
rect 28920 42838 28948 43386
rect 29380 42906 29408 43862
rect 29748 43790 29776 45970
rect 29932 45490 29960 46446
rect 30024 46073 30052 46446
rect 30010 46064 30066 46073
rect 30010 45999 30066 46008
rect 30012 45824 30064 45830
rect 30012 45766 30064 45772
rect 30024 45558 30052 45766
rect 30012 45552 30064 45558
rect 30012 45494 30064 45500
rect 29920 45484 29972 45490
rect 29920 45426 29972 45432
rect 29932 44878 29960 45426
rect 29920 44872 29972 44878
rect 29920 44814 29972 44820
rect 29736 43784 29788 43790
rect 29736 43726 29788 43732
rect 29748 42906 29776 43726
rect 29932 43314 29960 44814
rect 29920 43308 29972 43314
rect 29920 43250 29972 43256
rect 29368 42900 29420 42906
rect 29368 42842 29420 42848
rect 29736 42900 29788 42906
rect 29736 42842 29788 42848
rect 28908 42832 28960 42838
rect 28908 42774 28960 42780
rect 26700 42764 26752 42770
rect 26700 42706 26752 42712
rect 29000 42764 29052 42770
rect 29000 42706 29052 42712
rect 26712 41818 26740 42706
rect 29012 42362 29040 42706
rect 29380 42362 29408 42842
rect 29000 42356 29052 42362
rect 29000 42298 29052 42304
rect 29368 42356 29420 42362
rect 29368 42298 29420 42304
rect 29644 42356 29696 42362
rect 29644 42298 29696 42304
rect 27712 42016 27764 42022
rect 27712 41958 27764 41964
rect 24216 41812 24268 41818
rect 24216 41754 24268 41760
rect 26240 41812 26292 41818
rect 26240 41754 26292 41760
rect 26700 41812 26752 41818
rect 26700 41754 26752 41760
rect 27724 41750 27752 41958
rect 29380 41750 29408 42298
rect 27712 41744 27764 41750
rect 27712 41686 27764 41692
rect 29368 41744 29420 41750
rect 29368 41686 29420 41692
rect 29656 41274 29684 42298
rect 29748 41818 29776 42842
rect 30024 42362 30052 45494
rect 30116 44418 30144 49200
rect 30196 47456 30248 47462
rect 30196 47398 30248 47404
rect 30208 46714 30236 47398
rect 30564 47048 30616 47054
rect 30564 46990 30616 46996
rect 30288 46912 30340 46918
rect 30288 46854 30340 46860
rect 30380 46912 30432 46918
rect 30380 46854 30432 46860
rect 30196 46708 30248 46714
rect 30196 46650 30248 46656
rect 30300 46186 30328 46854
rect 30208 46158 30328 46186
rect 30208 44878 30236 46158
rect 30392 45966 30420 46854
rect 30576 46578 30604 46990
rect 30564 46572 30616 46578
rect 30564 46514 30616 46520
rect 30668 46442 30696 49286
rect 30838 49200 30894 50000
rect 31206 49314 31262 50000
rect 31206 49286 31432 49314
rect 31206 49200 31262 49286
rect 30852 47410 30880 49200
rect 30852 47382 30972 47410
rect 30840 47252 30892 47258
rect 30840 47194 30892 47200
rect 30748 46980 30800 46986
rect 30748 46922 30800 46928
rect 30760 46617 30788 46922
rect 30746 46608 30802 46617
rect 30746 46543 30802 46552
rect 30748 46504 30800 46510
rect 30748 46446 30800 46452
rect 30656 46436 30708 46442
rect 30656 46378 30708 46384
rect 30654 46064 30710 46073
rect 30654 45999 30710 46008
rect 30380 45960 30432 45966
rect 30380 45902 30432 45908
rect 30288 45892 30340 45898
rect 30288 45834 30340 45840
rect 30300 45490 30328 45834
rect 30288 45484 30340 45490
rect 30288 45426 30340 45432
rect 30196 44872 30248 44878
rect 30196 44814 30248 44820
rect 30380 44532 30432 44538
rect 30380 44474 30432 44480
rect 30116 44390 30236 44418
rect 30104 44328 30156 44334
rect 30104 44270 30156 44276
rect 30012 42356 30064 42362
rect 30012 42298 30064 42304
rect 29736 41812 29788 41818
rect 29736 41754 29788 41760
rect 29644 41268 29696 41274
rect 29644 41210 29696 41216
rect 20456 16546 20576 16574
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 20548 6730 20576 16546
rect 30116 12434 30144 44270
rect 30208 43994 30236 44390
rect 30196 43988 30248 43994
rect 30196 43930 30248 43936
rect 30288 43784 30340 43790
rect 30288 43726 30340 43732
rect 30300 43450 30328 43726
rect 30392 43450 30420 44474
rect 30668 44470 30696 45999
rect 30760 45966 30788 46446
rect 30852 46170 30880 47194
rect 30840 46164 30892 46170
rect 30840 46106 30892 46112
rect 30838 46064 30894 46073
rect 30838 45999 30894 46008
rect 30748 45960 30800 45966
rect 30748 45902 30800 45908
rect 30852 45898 30880 45999
rect 30840 45892 30892 45898
rect 30840 45834 30892 45840
rect 30944 45626 30972 47382
rect 31024 47048 31076 47054
rect 31024 46990 31076 46996
rect 31036 46714 31064 46990
rect 31024 46708 31076 46714
rect 31024 46650 31076 46656
rect 31036 46374 31064 46650
rect 31300 46504 31352 46510
rect 31300 46446 31352 46452
rect 31024 46368 31076 46374
rect 31024 46310 31076 46316
rect 31024 46096 31076 46102
rect 31024 46038 31076 46044
rect 31036 45830 31064 46038
rect 31312 45898 31340 46446
rect 31300 45892 31352 45898
rect 31300 45834 31352 45840
rect 31024 45824 31076 45830
rect 31024 45766 31076 45772
rect 30932 45620 30984 45626
rect 30932 45562 30984 45568
rect 30944 44538 30972 45562
rect 31312 45558 31340 45834
rect 31300 45552 31352 45558
rect 31300 45494 31352 45500
rect 31300 44872 31352 44878
rect 31300 44814 31352 44820
rect 30932 44532 30984 44538
rect 30932 44474 30984 44480
rect 30656 44464 30708 44470
rect 30656 44406 30708 44412
rect 30288 43444 30340 43450
rect 30288 43386 30340 43392
rect 30380 43444 30432 43450
rect 30380 43386 30432 43392
rect 30392 42906 30420 43386
rect 30472 43308 30524 43314
rect 30472 43250 30524 43256
rect 30484 42906 30512 43250
rect 30380 42900 30432 42906
rect 30380 42842 30432 42848
rect 30472 42900 30524 42906
rect 30472 42842 30524 42848
rect 30392 42294 30420 42842
rect 30484 42294 30512 42842
rect 31312 42770 31340 44814
rect 31404 43994 31432 49286
rect 31574 49200 31630 50000
rect 31942 49200 31998 50000
rect 32310 49200 32366 50000
rect 32678 49200 32734 50000
rect 33046 49200 33102 50000
rect 33414 49200 33470 50000
rect 33782 49200 33838 50000
rect 34150 49200 34206 50000
rect 34518 49200 34574 50000
rect 34886 49200 34942 50000
rect 35254 49314 35310 50000
rect 35254 49286 35480 49314
rect 35254 49200 35310 49286
rect 31484 45824 31536 45830
rect 31484 45766 31536 45772
rect 31392 43988 31444 43994
rect 31392 43930 31444 43936
rect 31496 43790 31524 45766
rect 31484 43784 31536 43790
rect 31484 43726 31536 43732
rect 31588 43314 31616 49200
rect 31668 46572 31720 46578
rect 31668 46514 31720 46520
rect 31760 46572 31812 46578
rect 31760 46514 31812 46520
rect 31680 46481 31708 46514
rect 31666 46472 31722 46481
rect 31666 46407 31722 46416
rect 31680 45898 31708 46407
rect 31668 45892 31720 45898
rect 31668 45834 31720 45840
rect 31772 45354 31800 46514
rect 31956 46102 31984 49200
rect 32324 46646 32352 49200
rect 32692 47258 32720 49200
rect 32956 47660 33008 47666
rect 32956 47602 33008 47608
rect 32680 47252 32732 47258
rect 32680 47194 32732 47200
rect 32404 46980 32456 46986
rect 32404 46922 32456 46928
rect 32220 46640 32272 46646
rect 32220 46582 32272 46588
rect 32312 46640 32364 46646
rect 32312 46582 32364 46588
rect 31944 46096 31996 46102
rect 31944 46038 31996 46044
rect 32036 45960 32088 45966
rect 32036 45902 32088 45908
rect 31852 45892 31904 45898
rect 31852 45834 31904 45840
rect 31864 45490 31892 45834
rect 32048 45490 32076 45902
rect 31852 45484 31904 45490
rect 31852 45426 31904 45432
rect 32036 45484 32088 45490
rect 32036 45426 32088 45432
rect 31760 45348 31812 45354
rect 31760 45290 31812 45296
rect 32232 44334 32260 46582
rect 32312 46504 32364 46510
rect 32416 46492 32444 46922
rect 32588 46912 32640 46918
rect 32588 46854 32640 46860
rect 32772 46912 32824 46918
rect 32824 46872 32904 46900
rect 32772 46854 32824 46860
rect 32600 46594 32628 46854
rect 32508 46578 32628 46594
rect 32496 46572 32628 46578
rect 32548 46566 32628 46572
rect 32496 46514 32548 46520
rect 32364 46464 32444 46492
rect 32312 46446 32364 46452
rect 32324 45626 32352 46446
rect 32508 46170 32536 46514
rect 32876 46510 32904 46872
rect 32864 46504 32916 46510
rect 32864 46446 32916 46452
rect 32772 46436 32824 46442
rect 32772 46378 32824 46384
rect 32496 46164 32548 46170
rect 32496 46106 32548 46112
rect 32784 46102 32812 46378
rect 32876 46345 32904 46446
rect 32968 46374 32996 47602
rect 33060 47002 33088 49200
rect 33324 47592 33376 47598
rect 33324 47534 33376 47540
rect 33060 46986 33272 47002
rect 33060 46980 33284 46986
rect 33060 46974 33232 46980
rect 33232 46922 33284 46928
rect 33336 46918 33364 47534
rect 33324 46912 33376 46918
rect 33324 46854 33376 46860
rect 33428 46617 33456 49200
rect 33600 47048 33652 47054
rect 33600 46990 33652 46996
rect 33612 46918 33640 46990
rect 33600 46912 33652 46918
rect 33600 46854 33652 46860
rect 33414 46608 33470 46617
rect 33414 46543 33470 46552
rect 33140 46504 33192 46510
rect 33138 46472 33140 46481
rect 33192 46472 33194 46481
rect 33138 46407 33194 46416
rect 32956 46368 33008 46374
rect 32862 46336 32918 46345
rect 32956 46310 33008 46316
rect 32862 46271 32918 46280
rect 33612 46170 33640 46854
rect 33600 46164 33652 46170
rect 33600 46106 33652 46112
rect 32772 46096 32824 46102
rect 32772 46038 32824 46044
rect 33140 45960 33192 45966
rect 33140 45902 33192 45908
rect 32588 45824 32640 45830
rect 32588 45766 32640 45772
rect 32864 45824 32916 45830
rect 32864 45766 32916 45772
rect 32312 45620 32364 45626
rect 32312 45562 32364 45568
rect 32600 45490 32628 45766
rect 32312 45484 32364 45490
rect 32312 45426 32364 45432
rect 32588 45484 32640 45490
rect 32588 45426 32640 45432
rect 32324 45082 32352 45426
rect 32312 45076 32364 45082
rect 32312 45018 32364 45024
rect 32496 44940 32548 44946
rect 32496 44882 32548 44888
rect 32220 44328 32272 44334
rect 32220 44270 32272 44276
rect 32508 43790 32536 44882
rect 32600 43994 32628 45426
rect 32876 45422 32904 45766
rect 32956 45620 33008 45626
rect 32956 45562 33008 45568
rect 32864 45416 32916 45422
rect 32864 45358 32916 45364
rect 32968 45354 32996 45562
rect 33152 45490 33180 45902
rect 33324 45892 33376 45898
rect 33324 45834 33376 45840
rect 33336 45558 33364 45834
rect 33600 45824 33652 45830
rect 33600 45766 33652 45772
rect 33612 45558 33640 45766
rect 33324 45552 33376 45558
rect 33324 45494 33376 45500
rect 33600 45552 33652 45558
rect 33600 45494 33652 45500
rect 33140 45484 33192 45490
rect 33140 45426 33192 45432
rect 32956 45348 33008 45354
rect 32956 45290 33008 45296
rect 32680 44872 32732 44878
rect 32680 44814 32732 44820
rect 32588 43988 32640 43994
rect 32588 43930 32640 43936
rect 32496 43784 32548 43790
rect 32496 43726 32548 43732
rect 32692 43722 32720 44814
rect 32968 44402 32996 45290
rect 33152 44470 33180 45426
rect 33336 44538 33364 45494
rect 33692 45416 33744 45422
rect 33692 45358 33744 45364
rect 33416 45280 33468 45286
rect 33416 45222 33468 45228
rect 33428 45014 33456 45222
rect 33416 45008 33468 45014
rect 33416 44950 33468 44956
rect 33324 44532 33376 44538
rect 33324 44474 33376 44480
rect 33140 44464 33192 44470
rect 33140 44406 33192 44412
rect 32956 44396 33008 44402
rect 32956 44338 33008 44344
rect 33152 43790 33180 44406
rect 33232 44328 33284 44334
rect 33232 44270 33284 44276
rect 33244 43858 33272 44270
rect 33704 43994 33732 45358
rect 33692 43988 33744 43994
rect 33692 43930 33744 43936
rect 33232 43852 33284 43858
rect 33232 43794 33284 43800
rect 33140 43784 33192 43790
rect 33140 43726 33192 43732
rect 32680 43716 32732 43722
rect 32680 43658 32732 43664
rect 32692 43450 32720 43658
rect 32680 43444 32732 43450
rect 32680 43386 32732 43392
rect 31576 43308 31628 43314
rect 31576 43250 31628 43256
rect 32692 42906 32720 43386
rect 32680 42900 32732 42906
rect 32680 42842 32732 42848
rect 31300 42764 31352 42770
rect 31300 42706 31352 42712
rect 33244 42362 33272 43794
rect 33796 43314 33824 49200
rect 34164 47530 34192 49200
rect 34152 47524 34204 47530
rect 34152 47466 34204 47472
rect 33980 47110 34284 47138
rect 33980 47002 34008 47110
rect 33888 46974 34008 47002
rect 34060 46980 34112 46986
rect 33888 46918 33916 46974
rect 34060 46922 34112 46928
rect 33876 46912 33928 46918
rect 33876 46854 33928 46860
rect 33968 46708 34020 46714
rect 33968 46650 34020 46656
rect 33980 46510 34008 46650
rect 33968 46504 34020 46510
rect 33968 46446 34020 46452
rect 33968 45960 34020 45966
rect 33968 45902 34020 45908
rect 33980 44946 34008 45902
rect 34072 45558 34100 46922
rect 34152 46640 34204 46646
rect 34152 46582 34204 46588
rect 34060 45552 34112 45558
rect 34060 45494 34112 45500
rect 34164 45082 34192 46582
rect 34256 46578 34284 47110
rect 34428 46912 34480 46918
rect 34428 46854 34480 46860
rect 34440 46714 34468 46854
rect 34428 46708 34480 46714
rect 34428 46650 34480 46656
rect 34244 46572 34296 46578
rect 34244 46514 34296 46520
rect 34256 45558 34284 46514
rect 34532 46374 34560 49200
rect 34900 47546 34928 49200
rect 34808 47518 34928 47546
rect 34612 47184 34664 47190
rect 34612 47126 34664 47132
rect 34704 47184 34756 47190
rect 34704 47126 34756 47132
rect 34428 46368 34480 46374
rect 34428 46310 34480 46316
rect 34520 46368 34572 46374
rect 34520 46310 34572 46316
rect 34336 46164 34388 46170
rect 34336 46106 34388 46112
rect 34348 45966 34376 46106
rect 34336 45960 34388 45966
rect 34336 45902 34388 45908
rect 34244 45552 34296 45558
rect 34244 45494 34296 45500
rect 34348 45490 34376 45902
rect 34440 45898 34468 46310
rect 34624 45966 34652 47126
rect 34716 46918 34744 47126
rect 34704 46912 34756 46918
rect 34704 46854 34756 46860
rect 34612 45960 34664 45966
rect 34612 45902 34664 45908
rect 34428 45892 34480 45898
rect 34428 45834 34480 45840
rect 34336 45484 34388 45490
rect 34336 45426 34388 45432
rect 34152 45076 34204 45082
rect 34152 45018 34204 45024
rect 33968 44940 34020 44946
rect 33968 44882 34020 44888
rect 33980 43790 34008 44882
rect 34348 44878 34376 45426
rect 34520 45416 34572 45422
rect 34520 45358 34572 45364
rect 34716 45370 34744 46854
rect 34808 46753 34836 47518
rect 35348 47456 35400 47462
rect 35348 47398 35400 47404
rect 34934 47356 35242 47365
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47291 35242 47300
rect 35360 47138 35388 47398
rect 35176 47110 35388 47138
rect 35176 47054 35204 47110
rect 35164 47048 35216 47054
rect 35164 46990 35216 46996
rect 35256 47048 35308 47054
rect 35256 46990 35308 46996
rect 34794 46744 34850 46753
rect 35268 46714 35296 46990
rect 35452 46986 35480 49286
rect 35622 49200 35678 50000
rect 35990 49200 36046 50000
rect 36358 49200 36414 50000
rect 36726 49314 36782 50000
rect 36726 49286 37044 49314
rect 36726 49200 36782 49286
rect 35440 46980 35492 46986
rect 35440 46922 35492 46928
rect 34794 46679 34850 46688
rect 35256 46708 35308 46714
rect 35256 46650 35308 46656
rect 34934 46268 35242 46277
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46203 35242 46212
rect 34980 45960 35032 45966
rect 34978 45928 34980 45937
rect 35032 45928 35034 45937
rect 34978 45863 35034 45872
rect 34336 44872 34388 44878
rect 34336 44814 34388 44820
rect 33968 43784 34020 43790
rect 33968 43726 34020 43732
rect 33784 43308 33836 43314
rect 33784 43250 33836 43256
rect 34348 42770 34376 44814
rect 34532 43382 34560 45358
rect 34716 45342 34836 45370
rect 34612 45280 34664 45286
rect 34612 45222 34664 45228
rect 34624 44402 34652 45222
rect 34612 44396 34664 44402
rect 34612 44338 34664 44344
rect 34716 43926 34744 45342
rect 34808 45286 34836 45342
rect 34796 45280 34848 45286
rect 34796 45222 34848 45228
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 35452 44810 35480 46922
rect 35532 46912 35584 46918
rect 35636 46889 35664 49200
rect 35532 46854 35584 46860
rect 35622 46880 35678 46889
rect 35544 45966 35572 46854
rect 35622 46815 35678 46824
rect 36004 46714 36032 49200
rect 36372 47274 36400 49200
rect 36372 47246 36676 47274
rect 36544 47116 36596 47122
rect 36544 47058 36596 47064
rect 36084 46980 36136 46986
rect 36084 46922 36136 46928
rect 35992 46708 36044 46714
rect 35992 46650 36044 46656
rect 35716 46504 35768 46510
rect 35716 46446 35768 46452
rect 35532 45960 35584 45966
rect 35532 45902 35584 45908
rect 35728 45948 35756 46446
rect 36096 45966 36124 46922
rect 36556 46918 36584 47058
rect 36648 46918 36676 47246
rect 36544 46912 36596 46918
rect 36544 46854 36596 46860
rect 36636 46912 36688 46918
rect 36636 46854 36688 46860
rect 36556 46578 36584 46854
rect 36360 46572 36412 46578
rect 36360 46514 36412 46520
rect 36544 46572 36596 46578
rect 36544 46514 36596 46520
rect 36176 46436 36228 46442
rect 36176 46378 36228 46384
rect 35900 45960 35952 45966
rect 35728 45920 35900 45948
rect 35728 45082 35756 45920
rect 35900 45902 35952 45908
rect 36084 45960 36136 45966
rect 36084 45902 36136 45908
rect 35808 45348 35860 45354
rect 35808 45290 35860 45296
rect 35716 45076 35768 45082
rect 35716 45018 35768 45024
rect 35820 44878 35848 45290
rect 35992 45280 36044 45286
rect 35992 45222 36044 45228
rect 35808 44872 35860 44878
rect 35808 44814 35860 44820
rect 35440 44804 35492 44810
rect 35440 44746 35492 44752
rect 35452 44554 35480 44746
rect 35452 44526 35572 44554
rect 35440 44464 35492 44470
rect 35440 44406 35492 44412
rect 34796 44396 34848 44402
rect 34796 44338 34848 44344
rect 34808 43994 34836 44338
rect 35348 44328 35400 44334
rect 35348 44270 35400 44276
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 35360 43994 35388 44270
rect 35452 44198 35480 44406
rect 35440 44192 35492 44198
rect 35440 44134 35492 44140
rect 34796 43988 34848 43994
rect 34796 43930 34848 43936
rect 35348 43988 35400 43994
rect 35348 43930 35400 43936
rect 34704 43920 34756 43926
rect 34704 43862 34756 43868
rect 34520 43376 34572 43382
rect 34520 43318 34572 43324
rect 34612 43308 34664 43314
rect 34612 43250 34664 43256
rect 34624 42906 34652 43250
rect 34612 42900 34664 42906
rect 34612 42842 34664 42848
rect 34336 42764 34388 42770
rect 34336 42706 34388 42712
rect 33232 42356 33284 42362
rect 33232 42298 33284 42304
rect 34348 42294 34376 42706
rect 34716 42362 34744 43862
rect 35452 43790 35480 44134
rect 35440 43784 35492 43790
rect 35440 43726 35492 43732
rect 35544 43450 35572 44526
rect 36004 44470 36032 45222
rect 35992 44464 36044 44470
rect 35992 44406 36044 44412
rect 36004 43790 36032 44406
rect 36188 44402 36216 46378
rect 36372 45966 36400 46514
rect 36360 45960 36412 45966
rect 36360 45902 36412 45908
rect 36268 45892 36320 45898
rect 36268 45834 36320 45840
rect 36280 45490 36308 45834
rect 36268 45484 36320 45490
rect 36268 45426 36320 45432
rect 36544 45484 36596 45490
rect 36544 45426 36596 45432
rect 36452 45416 36504 45422
rect 36452 45358 36504 45364
rect 36464 45014 36492 45358
rect 36452 45008 36504 45014
rect 36452 44950 36504 44956
rect 36360 44940 36412 44946
rect 36360 44882 36412 44888
rect 36372 44538 36400 44882
rect 36556 44878 36584 45426
rect 36544 44872 36596 44878
rect 36544 44814 36596 44820
rect 36360 44532 36412 44538
rect 36360 44474 36412 44480
rect 36176 44396 36228 44402
rect 36176 44338 36228 44344
rect 36372 43994 36400 44474
rect 36556 44402 36584 44814
rect 36544 44396 36596 44402
rect 36544 44338 36596 44344
rect 36360 43988 36412 43994
rect 36360 43930 36412 43936
rect 36648 43858 36676 46854
rect 36728 46504 36780 46510
rect 36728 46446 36780 46452
rect 36740 46170 36768 46446
rect 36728 46164 36780 46170
rect 36728 46106 36780 46112
rect 37016 46102 37044 49286
rect 37094 49200 37150 50000
rect 37462 49314 37518 50000
rect 37292 49286 37518 49314
rect 37108 47190 37136 49200
rect 37096 47184 37148 47190
rect 37096 47126 37148 47132
rect 37292 47054 37320 49286
rect 37462 49200 37518 49286
rect 37830 49200 37886 50000
rect 38198 49200 38254 50000
rect 38566 49200 38622 50000
rect 38934 49314 38990 50000
rect 38934 49286 39252 49314
rect 38934 49200 38990 49286
rect 37740 47524 37792 47530
rect 37740 47466 37792 47472
rect 37752 47054 37780 47466
rect 37280 47048 37332 47054
rect 37280 46990 37332 46996
rect 37740 47048 37792 47054
rect 37740 46990 37792 46996
rect 37004 46096 37056 46102
rect 37004 46038 37056 46044
rect 37096 45824 37148 45830
rect 37096 45766 37148 45772
rect 37108 45626 37136 45766
rect 37096 45620 37148 45626
rect 37096 45562 37148 45568
rect 37292 45422 37320 46990
rect 37648 46980 37700 46986
rect 37648 46922 37700 46928
rect 37556 46368 37608 46374
rect 37556 46310 37608 46316
rect 37568 45801 37596 46310
rect 37554 45792 37610 45801
rect 37554 45727 37610 45736
rect 37660 45490 37688 46922
rect 37648 45484 37700 45490
rect 37648 45426 37700 45432
rect 37280 45416 37332 45422
rect 37280 45358 37332 45364
rect 37660 45354 37688 45426
rect 37648 45348 37700 45354
rect 37648 45290 37700 45296
rect 37660 44946 37688 45290
rect 37556 44940 37608 44946
rect 37556 44882 37608 44888
rect 37648 44940 37700 44946
rect 37648 44882 37700 44888
rect 37464 44872 37516 44878
rect 37464 44814 37516 44820
rect 36912 44464 36964 44470
rect 36912 44406 36964 44412
rect 36924 43994 36952 44406
rect 36912 43988 36964 43994
rect 36912 43930 36964 43936
rect 36636 43852 36688 43858
rect 36636 43794 36688 43800
rect 35992 43784 36044 43790
rect 35992 43726 36044 43732
rect 36924 43722 36952 43930
rect 36544 43716 36596 43722
rect 36544 43658 36596 43664
rect 36912 43716 36964 43722
rect 36912 43658 36964 43664
rect 36556 43450 36584 43658
rect 35532 43444 35584 43450
rect 35532 43386 35584 43392
rect 36544 43444 36596 43450
rect 36544 43386 36596 43392
rect 35544 43314 35572 43386
rect 35532 43308 35584 43314
rect 35532 43250 35584 43256
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 37476 42362 37504 44814
rect 37568 44538 37596 44882
rect 37556 44532 37608 44538
rect 37556 44474 37608 44480
rect 37660 44334 37688 44882
rect 37752 44538 37780 46990
rect 37844 45082 37872 49200
rect 38108 46572 38160 46578
rect 38108 46514 38160 46520
rect 37924 46164 37976 46170
rect 37924 46106 37976 46112
rect 37936 46034 37964 46106
rect 38014 46064 38070 46073
rect 37924 46028 37976 46034
rect 38014 45999 38070 46008
rect 37924 45970 37976 45976
rect 37936 45626 37964 45970
rect 38028 45898 38056 45999
rect 38016 45892 38068 45898
rect 38016 45834 38068 45840
rect 37924 45620 37976 45626
rect 37924 45562 37976 45568
rect 37924 45484 37976 45490
rect 37924 45426 37976 45432
rect 37832 45076 37884 45082
rect 37832 45018 37884 45024
rect 37936 44878 37964 45426
rect 38016 45416 38068 45422
rect 38016 45358 38068 45364
rect 37924 44872 37976 44878
rect 37924 44814 37976 44820
rect 37740 44532 37792 44538
rect 37740 44474 37792 44480
rect 38028 44402 38056 45358
rect 38120 44742 38148 46514
rect 38212 45626 38240 49200
rect 38580 47054 38608 49200
rect 38752 47524 38804 47530
rect 38752 47466 38804 47472
rect 38844 47524 38896 47530
rect 38844 47466 38896 47472
rect 38568 47048 38620 47054
rect 38568 46990 38620 46996
rect 38764 46986 38792 47466
rect 38752 46980 38804 46986
rect 38752 46922 38804 46928
rect 38568 46912 38620 46918
rect 38620 46860 38700 46866
rect 38568 46854 38700 46860
rect 38580 46838 38700 46854
rect 38672 46578 38700 46838
rect 38856 46578 38884 47466
rect 39120 47048 39172 47054
rect 39120 46990 39172 46996
rect 38936 46912 38988 46918
rect 38936 46854 38988 46860
rect 38660 46572 38712 46578
rect 38660 46514 38712 46520
rect 38844 46572 38896 46578
rect 38844 46514 38896 46520
rect 38382 46472 38438 46481
rect 38382 46407 38438 46416
rect 38292 46164 38344 46170
rect 38292 46106 38344 46112
rect 38304 46034 38332 46106
rect 38292 46028 38344 46034
rect 38292 45970 38344 45976
rect 38396 45966 38424 46407
rect 38384 45960 38436 45966
rect 38384 45902 38436 45908
rect 38200 45620 38252 45626
rect 38200 45562 38252 45568
rect 38108 44736 38160 44742
rect 38108 44678 38160 44684
rect 38120 44538 38148 44678
rect 38108 44532 38160 44538
rect 38108 44474 38160 44480
rect 38016 44396 38068 44402
rect 38016 44338 38068 44344
rect 37648 44328 37700 44334
rect 37648 44270 37700 44276
rect 37660 43994 37688 44270
rect 37648 43988 37700 43994
rect 37648 43930 37700 43936
rect 37660 43450 37688 43930
rect 38028 43926 38056 44338
rect 38016 43920 38068 43926
rect 38016 43862 38068 43868
rect 38028 43450 38056 43862
rect 38672 43450 38700 46514
rect 38856 45966 38884 46514
rect 38948 46510 38976 46854
rect 39132 46617 39160 46990
rect 39118 46608 39174 46617
rect 39118 46543 39174 46552
rect 39224 46510 39252 49286
rect 39302 49200 39358 50000
rect 39670 49314 39726 50000
rect 39670 49286 39804 49314
rect 39670 49200 39726 49286
rect 38936 46504 38988 46510
rect 38936 46446 38988 46452
rect 39212 46504 39264 46510
rect 39212 46446 39264 46452
rect 38844 45960 38896 45966
rect 38764 45920 38844 45948
rect 38764 45830 38792 45920
rect 38844 45902 38896 45908
rect 38752 45824 38804 45830
rect 38752 45766 38804 45772
rect 37648 43444 37700 43450
rect 37648 43386 37700 43392
rect 38016 43444 38068 43450
rect 38016 43386 38068 43392
rect 38660 43444 38712 43450
rect 38660 43386 38712 43392
rect 37660 42906 37688 43386
rect 37648 42900 37700 42906
rect 37648 42842 37700 42848
rect 38028 42634 38056 43386
rect 38764 42770 38792 45766
rect 38948 45354 38976 46446
rect 39316 46170 39344 49200
rect 39776 47462 39804 49286
rect 40038 49200 40094 50000
rect 40406 49314 40462 50000
rect 40406 49286 40724 49314
rect 40406 49200 40462 49286
rect 39764 47456 39816 47462
rect 39764 47398 39816 47404
rect 39396 46708 39448 46714
rect 39396 46650 39448 46656
rect 39304 46164 39356 46170
rect 39304 46106 39356 46112
rect 39212 45960 39264 45966
rect 39212 45902 39264 45908
rect 39224 45558 39252 45902
rect 39408 45898 39436 46650
rect 39396 45892 39448 45898
rect 39396 45834 39448 45840
rect 39212 45552 39264 45558
rect 39212 45494 39264 45500
rect 39028 45484 39080 45490
rect 39028 45426 39080 45432
rect 38936 45348 38988 45354
rect 38936 45290 38988 45296
rect 39040 44538 39068 45426
rect 39776 45422 39804 47398
rect 40052 46578 40080 49200
rect 40696 47258 40724 49286
rect 40774 49200 40830 50000
rect 41142 49314 41198 50000
rect 41142 49286 41368 49314
rect 41142 49200 41198 49286
rect 40788 47530 40816 49200
rect 40776 47524 40828 47530
rect 40776 47466 40828 47472
rect 40684 47252 40736 47258
rect 40684 47194 40736 47200
rect 40224 47116 40276 47122
rect 40224 47058 40276 47064
rect 40132 47048 40184 47054
rect 40132 46990 40184 46996
rect 40144 46753 40172 46990
rect 40130 46744 40186 46753
rect 40130 46679 40186 46688
rect 40040 46572 40092 46578
rect 40040 46514 40092 46520
rect 39764 45416 39816 45422
rect 39764 45358 39816 45364
rect 39776 45082 39804 45358
rect 39948 45348 40000 45354
rect 39948 45290 40000 45296
rect 39764 45076 39816 45082
rect 39764 45018 39816 45024
rect 39028 44532 39080 44538
rect 39028 44474 39080 44480
rect 39960 43994 39988 45290
rect 40236 45014 40264 47058
rect 40684 47048 40736 47054
rect 40684 46990 40736 46996
rect 40696 46889 40724 46990
rect 40682 46880 40738 46889
rect 40682 46815 40738 46824
rect 40788 46102 40816 47466
rect 41340 46170 41368 49286
rect 41510 49200 41566 50000
rect 41878 49200 41934 50000
rect 42246 49200 42302 50000
rect 42614 49314 42670 50000
rect 42614 49286 42748 49314
rect 42614 49200 42670 49286
rect 41524 46170 41552 49200
rect 41892 46714 41920 49200
rect 41880 46708 41932 46714
rect 41880 46650 41932 46656
rect 42260 46578 42288 49200
rect 42720 47240 42748 49286
rect 42982 49200 43038 50000
rect 43350 49200 43406 50000
rect 43718 49200 43774 50000
rect 44086 49314 44142 50000
rect 43824 49286 44142 49314
rect 42800 47252 42852 47258
rect 42720 47212 42800 47240
rect 42800 47194 42852 47200
rect 42248 46572 42300 46578
rect 42248 46514 42300 46520
rect 41328 46164 41380 46170
rect 41328 46106 41380 46112
rect 41512 46164 41564 46170
rect 41512 46106 41564 46112
rect 40776 46096 40828 46102
rect 40776 46038 40828 46044
rect 42996 45937 43024 49200
rect 43364 47258 43392 49200
rect 43352 47252 43404 47258
rect 43352 47194 43404 47200
rect 43732 46578 43760 49200
rect 43720 46572 43772 46578
rect 43720 46514 43772 46520
rect 43824 46170 43852 49286
rect 44086 49200 44142 49286
rect 44454 49200 44510 50000
rect 44822 49200 44878 50000
rect 45190 49314 45246 50000
rect 44928 49286 45246 49314
rect 44468 46578 44496 49200
rect 44836 47258 44864 49200
rect 44824 47252 44876 47258
rect 44824 47194 44876 47200
rect 44456 46572 44508 46578
rect 44456 46514 44508 46520
rect 43812 46164 43864 46170
rect 43812 46106 43864 46112
rect 42982 45928 43038 45937
rect 42982 45863 43038 45872
rect 43824 45626 43852 46106
rect 43812 45620 43864 45626
rect 43812 45562 43864 45568
rect 44928 45554 44956 49286
rect 45190 49200 45246 49286
rect 45558 49314 45614 50000
rect 45558 49286 45876 49314
rect 45558 49200 45614 49286
rect 45848 47258 45876 49286
rect 45926 49200 45982 50000
rect 45940 47258 45968 49200
rect 45836 47252 45888 47258
rect 45836 47194 45888 47200
rect 45928 47252 45980 47258
rect 45928 47194 45980 47200
rect 44192 45526 44956 45554
rect 41972 45280 42024 45286
rect 41972 45222 42024 45228
rect 41236 45076 41288 45082
rect 41236 45018 41288 45024
rect 40224 45008 40276 45014
rect 40224 44950 40276 44956
rect 40236 44470 40264 44950
rect 41248 44538 41276 45018
rect 41984 44946 42012 45222
rect 44192 45082 44220 45526
rect 44180 45076 44232 45082
rect 44180 45018 44232 45024
rect 41972 44940 42024 44946
rect 41972 44882 42024 44888
rect 41236 44532 41288 44538
rect 41236 44474 41288 44480
rect 40224 44464 40276 44470
rect 40224 44406 40276 44412
rect 39948 43988 40000 43994
rect 39948 43930 40000 43936
rect 39960 43382 39988 43930
rect 39948 43376 40000 43382
rect 39948 43318 40000 43324
rect 39672 43104 39724 43110
rect 39672 43046 39724 43052
rect 39684 42770 39712 43046
rect 38752 42764 38804 42770
rect 38752 42706 38804 42712
rect 39672 42764 39724 42770
rect 39672 42706 39724 42712
rect 38016 42628 38068 42634
rect 38016 42570 38068 42576
rect 34704 42356 34756 42362
rect 34704 42298 34756 42304
rect 37464 42356 37516 42362
rect 37464 42298 37516 42304
rect 30380 42288 30432 42294
rect 30380 42230 30432 42236
rect 30472 42288 30524 42294
rect 30472 42230 30524 42236
rect 34336 42288 34388 42294
rect 34336 42230 34388 42236
rect 30484 42022 30512 42230
rect 30472 42016 30524 42022
rect 30472 41958 30524 41964
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 29656 12406 30144 12434
rect 22928 6792 22980 6798
rect 22928 6734 22980 6740
rect 20536 6724 20588 6730
rect 20536 6666 20588 6672
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 20548 6458 20576 6666
rect 20536 6452 20588 6458
rect 20536 6394 20588 6400
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 20548 5914 20576 6394
rect 22940 6322 22968 6734
rect 27160 6724 27212 6730
rect 27160 6666 27212 6672
rect 23204 6656 23256 6662
rect 23204 6598 23256 6604
rect 24768 6656 24820 6662
rect 24768 6598 24820 6604
rect 21088 6316 21140 6322
rect 21088 6258 21140 6264
rect 22928 6316 22980 6322
rect 22928 6258 22980 6264
rect 20536 5908 20588 5914
rect 20536 5850 20588 5856
rect 20260 5704 20312 5710
rect 20260 5646 20312 5652
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19432 5024 19484 5030
rect 19432 4966 19484 4972
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 16948 4616 17000 4622
rect 16948 4558 17000 4564
rect 15016 3936 15068 3942
rect 15016 3878 15068 3884
rect 16120 3936 16172 3942
rect 16120 3878 16172 3884
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4160 3528 4212 3534
rect 4160 3470 4212 3476
rect 5172 3528 5224 3534
rect 5172 3470 5224 3476
rect 6000 3528 6052 3534
rect 6000 3470 6052 3476
rect 6828 3528 6880 3534
rect 6828 3470 6880 3476
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 8484 3528 8536 3534
rect 8484 3470 8536 3476
rect 9312 3528 9364 3534
rect 9312 3470 9364 3476
rect 10140 3528 10192 3534
rect 10140 3470 10192 3476
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 11796 3528 11848 3534
rect 11796 3470 11848 3476
rect 12532 3528 12584 3534
rect 12532 3470 12584 3476
rect 13084 3528 13136 3534
rect 13084 3470 13136 3476
rect 13636 3528 13688 3534
rect 13636 3470 13688 3476
rect 4172 2938 4200 3470
rect 4080 2910 4200 2938
rect 4896 2916 4948 2922
rect 3148 2848 3200 2854
rect 3148 2790 3200 2796
rect 3884 2848 3936 2854
rect 3884 2790 3936 2796
rect 2596 2440 2648 2446
rect 2596 2382 2648 2388
rect 2608 800 2636 2382
rect 3160 800 3188 2790
rect 3516 2508 3568 2514
rect 3516 2450 3568 2456
rect 3528 800 3556 2450
rect 3896 800 3924 2790
rect 4080 2564 4108 2910
rect 4896 2858 4948 2864
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4080 2536 4292 2564
rect 4264 800 4292 2536
rect 4620 2440 4672 2446
rect 4620 2382 4672 2388
rect 4632 800 4660 2382
rect 4908 800 4936 2858
rect 5184 800 5212 3470
rect 5448 2984 5500 2990
rect 5448 2926 5500 2932
rect 5460 800 5488 2926
rect 5724 2440 5776 2446
rect 5724 2382 5776 2388
rect 5736 800 5764 2382
rect 6012 800 6040 3470
rect 6276 2916 6328 2922
rect 6276 2858 6328 2864
rect 6288 800 6316 2858
rect 6552 2848 6604 2854
rect 6552 2790 6604 2796
rect 6564 800 6592 2790
rect 6840 800 6868 3470
rect 7104 2576 7156 2582
rect 7104 2518 7156 2524
rect 7116 800 7144 2518
rect 7380 2372 7432 2378
rect 7380 2314 7432 2320
rect 7392 800 7420 2314
rect 7668 800 7696 3470
rect 7932 2984 7984 2990
rect 7932 2926 7984 2932
rect 7944 800 7972 2926
rect 8208 2508 8260 2514
rect 8208 2450 8260 2456
rect 8220 800 8248 2450
rect 8496 800 8524 3470
rect 8760 2916 8812 2922
rect 8760 2858 8812 2864
rect 8772 800 8800 2858
rect 9036 2848 9088 2854
rect 9036 2790 9088 2796
rect 9048 800 9076 2790
rect 9324 800 9352 3470
rect 9864 2984 9916 2990
rect 9864 2926 9916 2932
rect 9588 2576 9640 2582
rect 9588 2518 9640 2524
rect 9600 800 9628 2518
rect 9876 800 9904 2926
rect 10152 800 10180 3470
rect 10692 2848 10744 2854
rect 10692 2790 10744 2796
rect 10416 2508 10468 2514
rect 10416 2450 10468 2456
rect 10428 800 10456 2450
rect 10704 800 10732 2790
rect 10980 800 11008 3470
rect 11244 2916 11296 2922
rect 11244 2858 11296 2864
rect 11256 800 11284 2858
rect 11520 2576 11572 2582
rect 11520 2518 11572 2524
rect 11532 800 11560 2518
rect 11808 800 11836 3470
rect 12072 2848 12124 2854
rect 12072 2790 12124 2796
rect 12084 800 12112 2790
rect 12256 2440 12308 2446
rect 12256 2382 12308 2388
rect 12268 800 12296 2382
rect 12544 800 12572 3470
rect 12808 2508 12860 2514
rect 12808 2450 12860 2456
rect 12820 800 12848 2450
rect 13096 800 13124 3470
rect 13360 2916 13412 2922
rect 13360 2858 13412 2864
rect 13372 800 13400 2858
rect 13648 800 13676 3470
rect 14464 2916 14516 2922
rect 14464 2858 14516 2864
rect 13912 2848 13964 2854
rect 13912 2790 13964 2796
rect 13924 800 13952 2790
rect 14188 2576 14240 2582
rect 14188 2518 14240 2524
rect 14200 800 14228 2518
rect 14476 800 14504 2858
rect 14740 2508 14792 2514
rect 14740 2450 14792 2456
rect 14752 800 14780 2450
rect 15028 800 15056 3878
rect 15844 3596 15896 3602
rect 15844 3538 15896 3544
rect 15292 2848 15344 2854
rect 15292 2790 15344 2796
rect 15384 2848 15436 2854
rect 15384 2790 15436 2796
rect 15304 800 15332 2790
rect 15396 2650 15424 2790
rect 15384 2644 15436 2650
rect 15384 2586 15436 2592
rect 15568 2440 15620 2446
rect 15568 2382 15620 2388
rect 15580 800 15608 2382
rect 15856 800 15884 3538
rect 16132 800 16160 3878
rect 16396 3528 16448 3534
rect 16396 3470 16448 3476
rect 16304 2440 16356 2446
rect 16304 2382 16356 2388
rect 16316 1970 16344 2382
rect 16304 1964 16356 1970
rect 16304 1906 16356 1912
rect 16408 800 16436 3470
rect 16672 3052 16724 3058
rect 16672 2994 16724 3000
rect 16684 800 16712 2994
rect 16960 800 16988 4558
rect 19156 4004 19208 4010
rect 19156 3946 19208 3952
rect 18052 3936 18104 3942
rect 18052 3878 18104 3884
rect 18880 3936 18932 3942
rect 18880 3878 18932 3884
rect 17224 3664 17276 3670
rect 17224 3606 17276 3612
rect 17236 800 17264 3606
rect 17500 2916 17552 2922
rect 17500 2858 17552 2864
rect 17512 800 17540 2858
rect 17776 2848 17828 2854
rect 17776 2790 17828 2796
rect 17788 800 17816 2790
rect 18064 800 18092 3878
rect 18892 3602 18920 3878
rect 18604 3596 18656 3602
rect 18604 3538 18656 3544
rect 18880 3596 18932 3602
rect 18880 3538 18932 3544
rect 18420 3052 18472 3058
rect 18420 2994 18472 3000
rect 18328 2576 18380 2582
rect 18328 2518 18380 2524
rect 18340 800 18368 2518
rect 18432 2446 18460 2994
rect 18420 2440 18472 2446
rect 18420 2382 18472 2388
rect 18616 800 18644 3538
rect 18788 2916 18840 2922
rect 18788 2858 18840 2864
rect 18800 1578 18828 2858
rect 18972 2848 19024 2854
rect 18970 2816 18972 2825
rect 19024 2816 19026 2825
rect 18970 2751 19026 2760
rect 18880 2440 18932 2446
rect 18880 2382 18932 2388
rect 18892 2106 18920 2382
rect 18880 2100 18932 2106
rect 18880 2042 18932 2048
rect 18800 1550 18920 1578
rect 18892 800 18920 1550
rect 19168 800 19196 3946
rect 19248 3528 19300 3534
rect 19248 3470 19300 3476
rect 19260 3058 19288 3470
rect 19248 3052 19300 3058
rect 19248 2994 19300 3000
rect 19444 800 19472 4966
rect 20272 4690 20300 5646
rect 20548 5234 20576 5850
rect 21100 5710 21128 6258
rect 22560 6112 22612 6118
rect 22560 6054 22612 6060
rect 23112 6112 23164 6118
rect 23112 6054 23164 6060
rect 21088 5704 21140 5710
rect 21088 5646 21140 5652
rect 21100 5370 21128 5646
rect 22572 5642 22600 6054
rect 22928 5772 22980 5778
rect 22928 5714 22980 5720
rect 22560 5636 22612 5642
rect 22560 5578 22612 5584
rect 21732 5568 21784 5574
rect 21732 5510 21784 5516
rect 20812 5364 20864 5370
rect 20812 5306 20864 5312
rect 21088 5364 21140 5370
rect 21088 5306 21140 5312
rect 20536 5228 20588 5234
rect 20536 5170 20588 5176
rect 20352 5024 20404 5030
rect 20352 4966 20404 4972
rect 20260 4684 20312 4690
rect 20260 4626 20312 4632
rect 19984 4616 20036 4622
rect 19984 4558 20036 4564
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19996 2088 20024 4558
rect 20364 4554 20392 4966
rect 20352 4548 20404 4554
rect 20352 4490 20404 4496
rect 20824 4214 20852 5306
rect 21744 4554 21772 5510
rect 22192 4752 22244 4758
rect 22192 4694 22244 4700
rect 21088 4548 21140 4554
rect 21088 4490 21140 4496
rect 21732 4548 21784 4554
rect 21732 4490 21784 4496
rect 21916 4548 21968 4554
rect 21916 4490 21968 4496
rect 20812 4208 20864 4214
rect 20812 4150 20864 4156
rect 20824 3890 20852 4150
rect 20732 3862 20852 3890
rect 20260 3664 20312 3670
rect 20260 3606 20312 3612
rect 20076 3188 20128 3194
rect 20076 3130 20128 3136
rect 20088 2854 20116 3130
rect 20168 3052 20220 3058
rect 20168 2994 20220 3000
rect 20076 2848 20128 2854
rect 20076 2790 20128 2796
rect 20180 2446 20208 2994
rect 20168 2440 20220 2446
rect 20168 2382 20220 2388
rect 19720 2060 20024 2088
rect 19720 800 19748 2060
rect 19984 1964 20036 1970
rect 19984 1906 20036 1912
rect 19996 800 20024 1906
rect 20272 800 20300 3606
rect 20732 3534 20760 3862
rect 20812 3732 20864 3738
rect 20812 3674 20864 3680
rect 20720 3528 20772 3534
rect 20720 3470 20772 3476
rect 20628 3052 20680 3058
rect 20628 2994 20680 3000
rect 20640 2854 20668 2994
rect 20536 2848 20588 2854
rect 20536 2790 20588 2796
rect 20628 2848 20680 2854
rect 20628 2790 20680 2796
rect 20548 800 20576 2790
rect 20824 800 20852 3674
rect 21100 800 21128 4490
rect 21928 3942 21956 4490
rect 21916 3936 21968 3942
rect 21916 3878 21968 3884
rect 21364 3596 21416 3602
rect 21364 3538 21416 3544
rect 21376 800 21404 3538
rect 21640 2984 21692 2990
rect 21640 2926 21692 2932
rect 21652 800 21680 2926
rect 22008 2916 22060 2922
rect 22008 2858 22060 2864
rect 21916 2372 21968 2378
rect 21916 2314 21968 2320
rect 21928 800 21956 2314
rect 22020 2310 22048 2858
rect 22008 2304 22060 2310
rect 22008 2246 22060 2252
rect 22204 800 22232 4694
rect 22468 4072 22520 4078
rect 22468 4014 22520 4020
rect 22376 2984 22428 2990
rect 22376 2926 22428 2932
rect 22282 2816 22338 2825
rect 22282 2751 22338 2760
rect 22296 2514 22324 2751
rect 22284 2508 22336 2514
rect 22284 2450 22336 2456
rect 22388 2106 22416 2926
rect 22376 2100 22428 2106
rect 22376 2042 22428 2048
rect 22480 800 22508 4014
rect 22940 2774 22968 5714
rect 23124 5302 23152 6054
rect 23112 5296 23164 5302
rect 23112 5238 23164 5244
rect 23216 4554 23244 6598
rect 24032 6248 24084 6254
rect 24032 6190 24084 6196
rect 24044 5914 24072 6190
rect 24780 6186 24808 6598
rect 27172 6458 27200 6666
rect 27160 6452 27212 6458
rect 27160 6394 27212 6400
rect 25044 6384 25096 6390
rect 25044 6326 25096 6332
rect 24768 6180 24820 6186
rect 24768 6122 24820 6128
rect 24952 6180 25004 6186
rect 24952 6122 25004 6128
rect 24032 5908 24084 5914
rect 24032 5850 24084 5856
rect 24780 5846 24808 6122
rect 24768 5840 24820 5846
rect 24768 5782 24820 5788
rect 24584 5296 24636 5302
rect 24584 5238 24636 5244
rect 23480 5024 23532 5030
rect 23480 4966 23532 4972
rect 23204 4548 23256 4554
rect 23204 4490 23256 4496
rect 23020 3392 23072 3398
rect 23020 3334 23072 3340
rect 23032 3126 23060 3334
rect 23020 3120 23072 3126
rect 23020 3062 23072 3068
rect 23492 2774 23520 4966
rect 23572 4684 23624 4690
rect 23572 4626 23624 4632
rect 22940 2746 23060 2774
rect 22744 2508 22796 2514
rect 22744 2450 22796 2456
rect 22756 800 22784 2450
rect 23032 800 23060 2746
rect 23308 2746 23520 2774
rect 23308 800 23336 2746
rect 23584 800 23612 4626
rect 24596 4282 24624 5238
rect 24584 4276 24636 4282
rect 24584 4218 24636 4224
rect 24308 4208 24360 4214
rect 24308 4150 24360 4156
rect 24780 4162 24808 5782
rect 23664 4140 23716 4146
rect 23664 4082 23716 4088
rect 23676 3942 23704 4082
rect 23664 3936 23716 3942
rect 23664 3878 23716 3884
rect 23676 3534 23704 3878
rect 24124 3664 24176 3670
rect 24124 3606 24176 3612
rect 23664 3528 23716 3534
rect 23664 3470 23716 3476
rect 23676 2854 23704 3470
rect 24136 3126 24164 3606
rect 24124 3120 24176 3126
rect 24124 3062 24176 3068
rect 23848 2984 23900 2990
rect 23848 2926 23900 2932
rect 23664 2848 23716 2854
rect 23664 2790 23716 2796
rect 23676 2446 23704 2790
rect 23664 2440 23716 2446
rect 23664 2382 23716 2388
rect 23860 800 23888 2926
rect 24320 2650 24348 4150
rect 24780 4146 24900 4162
rect 24780 4140 24912 4146
rect 24780 4134 24860 4140
rect 24676 4072 24728 4078
rect 24676 4014 24728 4020
rect 24400 2984 24452 2990
rect 24400 2926 24452 2932
rect 24308 2644 24360 2650
rect 24308 2586 24360 2592
rect 24124 2508 24176 2514
rect 24124 2450 24176 2456
rect 24136 800 24164 2450
rect 24412 800 24440 2926
rect 24688 800 24716 4014
rect 24780 3942 24808 4134
rect 24860 4082 24912 4088
rect 24768 3936 24820 3942
rect 24768 3878 24820 3884
rect 24964 800 24992 6122
rect 25056 5914 25084 6326
rect 25872 6248 25924 6254
rect 25872 6190 25924 6196
rect 26608 6248 26660 6254
rect 26608 6190 26660 6196
rect 25044 5908 25096 5914
rect 25044 5850 25096 5856
rect 25884 5234 25912 6190
rect 26252 5778 26372 5794
rect 26240 5772 26372 5778
rect 26292 5766 26372 5772
rect 26240 5714 26292 5720
rect 26240 5636 26292 5642
rect 26240 5578 26292 5584
rect 26252 5234 26280 5578
rect 25872 5228 25924 5234
rect 25872 5170 25924 5176
rect 26240 5228 26292 5234
rect 26240 5170 26292 5176
rect 25228 5160 25280 5166
rect 25228 5102 25280 5108
rect 25044 3392 25096 3398
rect 25044 3334 25096 3340
rect 25056 3194 25084 3334
rect 25044 3188 25096 3194
rect 25044 3130 25096 3136
rect 25240 800 25268 5102
rect 26056 4684 26108 4690
rect 26056 4626 26108 4632
rect 25688 4548 25740 4554
rect 25688 4490 25740 4496
rect 25700 4282 25728 4490
rect 25688 4276 25740 4282
rect 25688 4218 25740 4224
rect 25320 3732 25372 3738
rect 25320 3674 25372 3680
rect 25332 3466 25360 3674
rect 25504 3596 25556 3602
rect 25504 3538 25556 3544
rect 25320 3460 25372 3466
rect 25320 3402 25372 3408
rect 25516 800 25544 3538
rect 25780 2984 25832 2990
rect 25780 2926 25832 2932
rect 25792 800 25820 2926
rect 26068 800 26096 4626
rect 26344 800 26372 5766
rect 26620 800 26648 6190
rect 26700 5636 26752 5642
rect 26700 5578 26752 5584
rect 26712 4486 26740 5578
rect 27172 4622 27200 6394
rect 29000 5704 29052 5710
rect 29000 5646 29052 5652
rect 27344 5568 27396 5574
rect 27344 5510 27396 5516
rect 28540 5568 28592 5574
rect 28540 5510 28592 5516
rect 27356 5302 27384 5510
rect 28552 5302 28580 5510
rect 27344 5296 27396 5302
rect 27344 5238 27396 5244
rect 28540 5296 28592 5302
rect 28540 5238 28592 5244
rect 27344 5160 27396 5166
rect 27344 5102 27396 5108
rect 28448 5160 28500 5166
rect 28448 5102 28500 5108
rect 27356 4826 27384 5102
rect 27804 5092 27856 5098
rect 27804 5034 27856 5040
rect 27344 4820 27396 4826
rect 27344 4762 27396 4768
rect 27160 4616 27212 4622
rect 27160 4558 27212 4564
rect 26700 4480 26752 4486
rect 26700 4422 26752 4428
rect 26712 3534 26740 4422
rect 27712 4208 27764 4214
rect 27712 4150 27764 4156
rect 27436 4072 27488 4078
rect 27436 4014 27488 4020
rect 26700 3528 26752 3534
rect 26700 3470 26752 3476
rect 27252 2984 27304 2990
rect 27252 2926 27304 2932
rect 26884 2916 26936 2922
rect 26884 2858 26936 2864
rect 26896 800 26924 2858
rect 27264 2650 27292 2926
rect 27252 2644 27304 2650
rect 27252 2586 27304 2592
rect 27160 2372 27212 2378
rect 27160 2314 27212 2320
rect 27172 800 27200 2314
rect 27448 800 27476 4014
rect 27724 3738 27752 4150
rect 27712 3732 27764 3738
rect 27712 3674 27764 3680
rect 27816 2530 27844 5034
rect 28460 4010 28488 5102
rect 29012 4690 29040 5646
rect 29092 5636 29144 5642
rect 29092 5578 29144 5584
rect 29104 5302 29132 5578
rect 29092 5296 29144 5302
rect 29092 5238 29144 5244
rect 29184 5160 29236 5166
rect 29184 5102 29236 5108
rect 29092 5024 29144 5030
rect 29092 4966 29144 4972
rect 28816 4684 28868 4690
rect 28816 4626 28868 4632
rect 29000 4684 29052 4690
rect 29000 4626 29052 4632
rect 28448 4004 28500 4010
rect 28448 3946 28500 3952
rect 27988 3664 28040 3670
rect 27988 3606 28040 3612
rect 27724 2502 27844 2530
rect 27724 800 27752 2502
rect 28000 800 28028 3606
rect 28264 3596 28316 3602
rect 28264 3538 28316 3544
rect 28276 800 28304 3538
rect 28356 3460 28408 3466
rect 28356 3402 28408 3408
rect 28368 2922 28396 3402
rect 28540 2984 28592 2990
rect 28540 2926 28592 2932
rect 28356 2916 28408 2922
rect 28356 2858 28408 2864
rect 28552 800 28580 2926
rect 28828 800 28856 4626
rect 29000 4548 29052 4554
rect 29104 4536 29132 4966
rect 29052 4508 29132 4536
rect 29000 4490 29052 4496
rect 28908 4072 28960 4078
rect 28908 4014 28960 4020
rect 28920 3738 28948 4014
rect 29092 3936 29144 3942
rect 29092 3878 29144 3884
rect 28908 3732 28960 3738
rect 28908 3674 28960 3680
rect 28908 3392 28960 3398
rect 28908 3334 28960 3340
rect 28920 3126 28948 3334
rect 28908 3120 28960 3126
rect 28908 3062 28960 3068
rect 29104 800 29132 3878
rect 29196 3670 29224 5102
rect 29184 3664 29236 3670
rect 29184 3606 29236 3612
rect 29368 2984 29420 2990
rect 29368 2926 29420 2932
rect 29380 800 29408 2926
rect 29656 800 29684 12406
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 29828 5228 29880 5234
rect 29828 5170 29880 5176
rect 29840 4146 29868 5170
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 29828 4140 29880 4146
rect 29828 4082 29880 4088
rect 29736 4072 29788 4078
rect 29736 4014 29788 4020
rect 29748 3738 29776 4014
rect 29736 3732 29788 3738
rect 29736 3674 29788 3680
rect 29840 3466 29868 4082
rect 29920 3936 29972 3942
rect 29920 3878 29972 3884
rect 29828 3460 29880 3466
rect 29828 3402 29880 3408
rect 29736 2848 29788 2854
rect 29736 2790 29788 2796
rect 29748 2650 29776 2790
rect 29736 2644 29788 2650
rect 29736 2586 29788 2592
rect 29932 800 29960 3878
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 32956 3664 33008 3670
rect 32956 3606 33008 3612
rect 36820 3664 36872 3670
rect 36820 3606 36872 3612
rect 30196 3596 30248 3602
rect 30196 3538 30248 3544
rect 30208 800 30236 3538
rect 30288 3528 30340 3534
rect 30288 3470 30340 3476
rect 31116 3528 31168 3534
rect 31116 3470 31168 3476
rect 31852 3528 31904 3534
rect 31852 3470 31904 3476
rect 32404 3528 32456 3534
rect 32404 3470 32456 3476
rect 30300 2650 30328 3470
rect 30932 3460 30984 3466
rect 30932 3402 30984 3408
rect 30944 3058 30972 3402
rect 31024 3188 31076 3194
rect 31024 3130 31076 3136
rect 30932 3052 30984 3058
rect 30932 2994 30984 3000
rect 30840 2916 30892 2922
rect 30760 2876 30840 2904
rect 30288 2644 30340 2650
rect 30288 2586 30340 2592
rect 30472 2372 30524 2378
rect 30472 2314 30524 2320
rect 30484 800 30512 2314
rect 30760 800 30788 2876
rect 30840 2858 30892 2864
rect 30944 2774 30972 2994
rect 30852 2746 30972 2774
rect 30852 2446 30880 2746
rect 31036 2650 31064 3130
rect 31024 2644 31076 2650
rect 31024 2586 31076 2592
rect 30840 2440 30892 2446
rect 30840 2382 30892 2388
rect 31128 1850 31156 3470
rect 31668 2984 31720 2990
rect 31668 2926 31720 2932
rect 31576 2916 31628 2922
rect 31576 2858 31628 2864
rect 31300 2508 31352 2514
rect 31300 2450 31352 2456
rect 31036 1822 31156 1850
rect 31036 800 31064 1822
rect 31312 800 31340 2450
rect 31588 800 31616 2858
rect 31680 2650 31708 2926
rect 31668 2644 31720 2650
rect 31668 2586 31720 2592
rect 31864 800 31892 3470
rect 32128 2984 32180 2990
rect 32128 2926 32180 2932
rect 32140 800 32168 2926
rect 32416 800 32444 3470
rect 32680 3052 32732 3058
rect 32680 2994 32732 3000
rect 32692 800 32720 2994
rect 32968 800 32996 3606
rect 34796 3596 34848 3602
rect 34796 3538 34848 3544
rect 34336 3528 34388 3534
rect 34336 3470 34388 3476
rect 34060 2984 34112 2990
rect 34060 2926 34112 2932
rect 33508 2916 33560 2922
rect 33508 2858 33560 2864
rect 33232 2576 33284 2582
rect 33232 2518 33284 2524
rect 33244 800 33272 2518
rect 33520 800 33548 2858
rect 33784 2440 33836 2446
rect 33784 2382 33836 2388
rect 33796 800 33824 2382
rect 34072 800 34100 2926
rect 34348 800 34376 3470
rect 34612 2508 34664 2514
rect 34612 2450 34664 2456
rect 34624 800 34652 2450
rect 34808 1850 34836 3538
rect 35716 3528 35768 3534
rect 35716 3470 35768 3476
rect 36268 3528 36320 3534
rect 36268 3470 36320 3476
rect 35348 2916 35400 2922
rect 35348 2858 35400 2864
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 34808 1822 34928 1850
rect 34900 800 34928 1822
rect 35360 1442 35388 2858
rect 35440 2576 35492 2582
rect 35440 2518 35492 2524
rect 35176 1414 35388 1442
rect 35176 800 35204 1414
rect 35452 800 35480 2518
rect 35728 800 35756 3470
rect 35992 2848 36044 2854
rect 35992 2790 36044 2796
rect 36004 800 36032 2790
rect 36280 800 36308 3470
rect 36544 2440 36596 2446
rect 36544 2382 36596 2388
rect 36556 800 36584 2382
rect 36832 800 36860 3606
rect 37648 3528 37700 3534
rect 37648 3470 37700 3476
rect 38200 3528 38252 3534
rect 38200 3470 38252 3476
rect 39580 3528 39632 3534
rect 39580 3470 39632 3476
rect 40408 3528 40460 3534
rect 40408 3470 40460 3476
rect 40960 3528 41012 3534
rect 40960 3470 41012 3476
rect 41512 3528 41564 3534
rect 41512 3470 41564 3476
rect 42892 3528 42944 3534
rect 42892 3470 42944 3476
rect 43168 3528 43220 3534
rect 43168 3470 43220 3476
rect 44824 3528 44876 3534
rect 44824 3470 44876 3476
rect 45652 3528 45704 3534
rect 45652 3470 45704 3476
rect 46480 3528 46532 3534
rect 46480 3470 46532 3476
rect 46756 3528 46808 3534
rect 46756 3470 46808 3476
rect 47308 3528 47360 3534
rect 47308 3470 47360 3476
rect 37096 2984 37148 2990
rect 37096 2926 37148 2932
rect 37108 800 37136 2926
rect 37372 2508 37424 2514
rect 37372 2450 37424 2456
rect 37384 800 37412 2450
rect 37660 800 37688 3470
rect 37924 2916 37976 2922
rect 37924 2858 37976 2864
rect 37936 800 37964 2858
rect 38212 800 38240 3470
rect 38752 2984 38804 2990
rect 38752 2926 38804 2932
rect 38476 2576 38528 2582
rect 38476 2518 38528 2524
rect 38488 800 38516 2518
rect 38764 800 38792 2926
rect 39028 2848 39080 2854
rect 39028 2790 39080 2796
rect 39040 800 39068 2790
rect 39304 2508 39356 2514
rect 39304 2450 39356 2456
rect 39316 800 39344 2450
rect 39592 800 39620 3470
rect 40132 2848 40184 2854
rect 40132 2790 40184 2796
rect 39856 2440 39908 2446
rect 39856 2382 39908 2388
rect 39868 800 39896 2382
rect 40144 800 40172 2790
rect 40420 800 40448 3470
rect 40684 2984 40736 2990
rect 40684 2926 40736 2932
rect 40696 800 40724 2926
rect 40972 800 41000 3470
rect 41236 2508 41288 2514
rect 41236 2450 41288 2456
rect 41248 800 41276 2450
rect 41524 800 41552 3470
rect 42616 2984 42668 2990
rect 42616 2926 42668 2932
rect 42064 2848 42116 2854
rect 42064 2790 42116 2796
rect 41788 2440 41840 2446
rect 41788 2382 41840 2388
rect 41800 800 41828 2382
rect 42076 800 42104 2790
rect 42340 2576 42392 2582
rect 42340 2518 42392 2524
rect 42352 800 42380 2518
rect 42628 800 42656 2926
rect 42904 800 42932 3470
rect 43180 800 43208 3470
rect 44548 2984 44600 2990
rect 44548 2926 44600 2932
rect 43444 2848 43496 2854
rect 43444 2790 43496 2796
rect 43996 2848 44048 2854
rect 43996 2790 44048 2796
rect 43456 800 43484 2790
rect 43720 2508 43772 2514
rect 43720 2450 43772 2456
rect 43732 800 43760 2450
rect 44008 800 44036 2790
rect 44272 2372 44324 2378
rect 44272 2314 44324 2320
rect 44284 800 44312 2314
rect 44560 800 44588 2926
rect 44836 800 44864 3470
rect 45376 2848 45428 2854
rect 45376 2790 45428 2796
rect 45100 2576 45152 2582
rect 45100 2518 45152 2524
rect 45112 800 45140 2518
rect 45388 800 45416 2790
rect 45664 800 45692 3470
rect 45928 2848 45980 2854
rect 45928 2790 45980 2796
rect 45940 800 45968 2790
rect 46204 2440 46256 2446
rect 46204 2382 46256 2388
rect 46216 800 46244 2382
rect 46492 800 46520 3470
rect 46768 800 46796 3470
rect 47032 2848 47084 2854
rect 47032 2790 47084 2796
rect 47044 800 47072 2790
rect 47320 800 47348 3470
rect 2410 0 2466 800
rect 2502 0 2558 800
rect 2594 0 2650 800
rect 2686 0 2742 800
rect 2778 0 2834 800
rect 2870 0 2926 800
rect 2962 0 3018 800
rect 3054 0 3110 800
rect 3146 0 3202 800
rect 3238 0 3294 800
rect 3330 0 3386 800
rect 3422 0 3478 800
rect 3514 0 3570 800
rect 3606 0 3662 800
rect 3698 0 3754 800
rect 3790 0 3846 800
rect 3882 0 3938 800
rect 3974 0 4030 800
rect 4066 0 4122 800
rect 4158 0 4214 800
rect 4250 0 4306 800
rect 4342 0 4398 800
rect 4434 0 4490 800
rect 4526 0 4582 800
rect 4618 0 4674 800
rect 4710 0 4766 800
rect 4802 0 4858 800
rect 4894 0 4950 800
rect 4986 0 5042 800
rect 5078 0 5134 800
rect 5170 0 5226 800
rect 5262 0 5318 800
rect 5354 0 5410 800
rect 5446 0 5502 800
rect 5538 0 5594 800
rect 5630 0 5686 800
rect 5722 0 5778 800
rect 5814 0 5870 800
rect 5906 0 5962 800
rect 5998 0 6054 800
rect 6090 0 6146 800
rect 6182 0 6238 800
rect 6274 0 6330 800
rect 6366 0 6422 800
rect 6458 0 6514 800
rect 6550 0 6606 800
rect 6642 0 6698 800
rect 6734 0 6790 800
rect 6826 0 6882 800
rect 6918 0 6974 800
rect 7010 0 7066 800
rect 7102 0 7158 800
rect 7194 0 7250 800
rect 7286 0 7342 800
rect 7378 0 7434 800
rect 7470 0 7526 800
rect 7562 0 7618 800
rect 7654 0 7710 800
rect 7746 0 7802 800
rect 7838 0 7894 800
rect 7930 0 7986 800
rect 8022 0 8078 800
rect 8114 0 8170 800
rect 8206 0 8262 800
rect 8298 0 8354 800
rect 8390 0 8446 800
rect 8482 0 8538 800
rect 8574 0 8630 800
rect 8666 0 8722 800
rect 8758 0 8814 800
rect 8850 0 8906 800
rect 8942 0 8998 800
rect 9034 0 9090 800
rect 9126 0 9182 800
rect 9218 0 9274 800
rect 9310 0 9366 800
rect 9402 0 9458 800
rect 9494 0 9550 800
rect 9586 0 9642 800
rect 9678 0 9734 800
rect 9770 0 9826 800
rect 9862 0 9918 800
rect 9954 0 10010 800
rect 10046 0 10102 800
rect 10138 0 10194 800
rect 10230 0 10286 800
rect 10322 0 10378 800
rect 10414 0 10470 800
rect 10506 0 10562 800
rect 10598 0 10654 800
rect 10690 0 10746 800
rect 10782 0 10838 800
rect 10874 0 10930 800
rect 10966 0 11022 800
rect 11058 0 11114 800
rect 11150 0 11206 800
rect 11242 0 11298 800
rect 11334 0 11390 800
rect 11426 0 11482 800
rect 11518 0 11574 800
rect 11610 0 11666 800
rect 11702 0 11758 800
rect 11794 0 11850 800
rect 11886 0 11942 800
rect 11978 0 12034 800
rect 12070 0 12126 800
rect 12162 0 12218 800
rect 12254 0 12310 800
rect 12346 0 12402 800
rect 12438 0 12494 800
rect 12530 0 12586 800
rect 12622 0 12678 800
rect 12714 0 12770 800
rect 12806 0 12862 800
rect 12898 0 12954 800
rect 12990 0 13046 800
rect 13082 0 13138 800
rect 13174 0 13230 800
rect 13266 0 13322 800
rect 13358 0 13414 800
rect 13450 0 13506 800
rect 13542 0 13598 800
rect 13634 0 13690 800
rect 13726 0 13782 800
rect 13818 0 13874 800
rect 13910 0 13966 800
rect 14002 0 14058 800
rect 14094 0 14150 800
rect 14186 0 14242 800
rect 14278 0 14334 800
rect 14370 0 14426 800
rect 14462 0 14518 800
rect 14554 0 14610 800
rect 14646 0 14702 800
rect 14738 0 14794 800
rect 14830 0 14886 800
rect 14922 0 14978 800
rect 15014 0 15070 800
rect 15106 0 15162 800
rect 15198 0 15254 800
rect 15290 0 15346 800
rect 15382 0 15438 800
rect 15474 0 15530 800
rect 15566 0 15622 800
rect 15658 0 15714 800
rect 15750 0 15806 800
rect 15842 0 15898 800
rect 15934 0 15990 800
rect 16026 0 16082 800
rect 16118 0 16174 800
rect 16210 0 16266 800
rect 16302 0 16358 800
rect 16394 0 16450 800
rect 16486 0 16542 800
rect 16578 0 16634 800
rect 16670 0 16726 800
rect 16762 0 16818 800
rect 16854 0 16910 800
rect 16946 0 17002 800
rect 17038 0 17094 800
rect 17130 0 17186 800
rect 17222 0 17278 800
rect 17314 0 17370 800
rect 17406 0 17462 800
rect 17498 0 17554 800
rect 17590 0 17646 800
rect 17682 0 17738 800
rect 17774 0 17830 800
rect 17866 0 17922 800
rect 17958 0 18014 800
rect 18050 0 18106 800
rect 18142 0 18198 800
rect 18234 0 18290 800
rect 18326 0 18382 800
rect 18418 0 18474 800
rect 18510 0 18566 800
rect 18602 0 18658 800
rect 18694 0 18750 800
rect 18786 0 18842 800
rect 18878 0 18934 800
rect 18970 0 19026 800
rect 19062 0 19118 800
rect 19154 0 19210 800
rect 19246 0 19302 800
rect 19338 0 19394 800
rect 19430 0 19486 800
rect 19522 0 19578 800
rect 19614 0 19670 800
rect 19706 0 19762 800
rect 19798 0 19854 800
rect 19890 0 19946 800
rect 19982 0 20038 800
rect 20074 0 20130 800
rect 20166 0 20222 800
rect 20258 0 20314 800
rect 20350 0 20406 800
rect 20442 0 20498 800
rect 20534 0 20590 800
rect 20626 0 20682 800
rect 20718 0 20774 800
rect 20810 0 20866 800
rect 20902 0 20958 800
rect 20994 0 21050 800
rect 21086 0 21142 800
rect 21178 0 21234 800
rect 21270 0 21326 800
rect 21362 0 21418 800
rect 21454 0 21510 800
rect 21546 0 21602 800
rect 21638 0 21694 800
rect 21730 0 21786 800
rect 21822 0 21878 800
rect 21914 0 21970 800
rect 22006 0 22062 800
rect 22098 0 22154 800
rect 22190 0 22246 800
rect 22282 0 22338 800
rect 22374 0 22430 800
rect 22466 0 22522 800
rect 22558 0 22614 800
rect 22650 0 22706 800
rect 22742 0 22798 800
rect 22834 0 22890 800
rect 22926 0 22982 800
rect 23018 0 23074 800
rect 23110 0 23166 800
rect 23202 0 23258 800
rect 23294 0 23350 800
rect 23386 0 23442 800
rect 23478 0 23534 800
rect 23570 0 23626 800
rect 23662 0 23718 800
rect 23754 0 23810 800
rect 23846 0 23902 800
rect 23938 0 23994 800
rect 24030 0 24086 800
rect 24122 0 24178 800
rect 24214 0 24270 800
rect 24306 0 24362 800
rect 24398 0 24454 800
rect 24490 0 24546 800
rect 24582 0 24638 800
rect 24674 0 24730 800
rect 24766 0 24822 800
rect 24858 0 24914 800
rect 24950 0 25006 800
rect 25042 0 25098 800
rect 25134 0 25190 800
rect 25226 0 25282 800
rect 25318 0 25374 800
rect 25410 0 25466 800
rect 25502 0 25558 800
rect 25594 0 25650 800
rect 25686 0 25742 800
rect 25778 0 25834 800
rect 25870 0 25926 800
rect 25962 0 26018 800
rect 26054 0 26110 800
rect 26146 0 26202 800
rect 26238 0 26294 800
rect 26330 0 26386 800
rect 26422 0 26478 800
rect 26514 0 26570 800
rect 26606 0 26662 800
rect 26698 0 26754 800
rect 26790 0 26846 800
rect 26882 0 26938 800
rect 26974 0 27030 800
rect 27066 0 27122 800
rect 27158 0 27214 800
rect 27250 0 27306 800
rect 27342 0 27398 800
rect 27434 0 27490 800
rect 27526 0 27582 800
rect 27618 0 27674 800
rect 27710 0 27766 800
rect 27802 0 27858 800
rect 27894 0 27950 800
rect 27986 0 28042 800
rect 28078 0 28134 800
rect 28170 0 28226 800
rect 28262 0 28318 800
rect 28354 0 28410 800
rect 28446 0 28502 800
rect 28538 0 28594 800
rect 28630 0 28686 800
rect 28722 0 28778 800
rect 28814 0 28870 800
rect 28906 0 28962 800
rect 28998 0 29054 800
rect 29090 0 29146 800
rect 29182 0 29238 800
rect 29274 0 29330 800
rect 29366 0 29422 800
rect 29458 0 29514 800
rect 29550 0 29606 800
rect 29642 0 29698 800
rect 29734 0 29790 800
rect 29826 0 29882 800
rect 29918 0 29974 800
rect 30010 0 30066 800
rect 30102 0 30158 800
rect 30194 0 30250 800
rect 30286 0 30342 800
rect 30378 0 30434 800
rect 30470 0 30526 800
rect 30562 0 30618 800
rect 30654 0 30710 800
rect 30746 0 30802 800
rect 30838 0 30894 800
rect 30930 0 30986 800
rect 31022 0 31078 800
rect 31114 0 31170 800
rect 31206 0 31262 800
rect 31298 0 31354 800
rect 31390 0 31446 800
rect 31482 0 31538 800
rect 31574 0 31630 800
rect 31666 0 31722 800
rect 31758 0 31814 800
rect 31850 0 31906 800
rect 31942 0 31998 800
rect 32034 0 32090 800
rect 32126 0 32182 800
rect 32218 0 32274 800
rect 32310 0 32366 800
rect 32402 0 32458 800
rect 32494 0 32550 800
rect 32586 0 32642 800
rect 32678 0 32734 800
rect 32770 0 32826 800
rect 32862 0 32918 800
rect 32954 0 33010 800
rect 33046 0 33102 800
rect 33138 0 33194 800
rect 33230 0 33286 800
rect 33322 0 33378 800
rect 33414 0 33470 800
rect 33506 0 33562 800
rect 33598 0 33654 800
rect 33690 0 33746 800
rect 33782 0 33838 800
rect 33874 0 33930 800
rect 33966 0 34022 800
rect 34058 0 34114 800
rect 34150 0 34206 800
rect 34242 0 34298 800
rect 34334 0 34390 800
rect 34426 0 34482 800
rect 34518 0 34574 800
rect 34610 0 34666 800
rect 34702 0 34758 800
rect 34794 0 34850 800
rect 34886 0 34942 800
rect 34978 0 35034 800
rect 35070 0 35126 800
rect 35162 0 35218 800
rect 35254 0 35310 800
rect 35346 0 35402 800
rect 35438 0 35494 800
rect 35530 0 35586 800
rect 35622 0 35678 800
rect 35714 0 35770 800
rect 35806 0 35862 800
rect 35898 0 35954 800
rect 35990 0 36046 800
rect 36082 0 36138 800
rect 36174 0 36230 800
rect 36266 0 36322 800
rect 36358 0 36414 800
rect 36450 0 36506 800
rect 36542 0 36598 800
rect 36634 0 36690 800
rect 36726 0 36782 800
rect 36818 0 36874 800
rect 36910 0 36966 800
rect 37002 0 37058 800
rect 37094 0 37150 800
rect 37186 0 37242 800
rect 37278 0 37334 800
rect 37370 0 37426 800
rect 37462 0 37518 800
rect 37554 0 37610 800
rect 37646 0 37702 800
rect 37738 0 37794 800
rect 37830 0 37886 800
rect 37922 0 37978 800
rect 38014 0 38070 800
rect 38106 0 38162 800
rect 38198 0 38254 800
rect 38290 0 38346 800
rect 38382 0 38438 800
rect 38474 0 38530 800
rect 38566 0 38622 800
rect 38658 0 38714 800
rect 38750 0 38806 800
rect 38842 0 38898 800
rect 38934 0 38990 800
rect 39026 0 39082 800
rect 39118 0 39174 800
rect 39210 0 39266 800
rect 39302 0 39358 800
rect 39394 0 39450 800
rect 39486 0 39542 800
rect 39578 0 39634 800
rect 39670 0 39726 800
rect 39762 0 39818 800
rect 39854 0 39910 800
rect 39946 0 40002 800
rect 40038 0 40094 800
rect 40130 0 40186 800
rect 40222 0 40278 800
rect 40314 0 40370 800
rect 40406 0 40462 800
rect 40498 0 40554 800
rect 40590 0 40646 800
rect 40682 0 40738 800
rect 40774 0 40830 800
rect 40866 0 40922 800
rect 40958 0 41014 800
rect 41050 0 41106 800
rect 41142 0 41198 800
rect 41234 0 41290 800
rect 41326 0 41382 800
rect 41418 0 41474 800
rect 41510 0 41566 800
rect 41602 0 41658 800
rect 41694 0 41750 800
rect 41786 0 41842 800
rect 41878 0 41934 800
rect 41970 0 42026 800
rect 42062 0 42118 800
rect 42154 0 42210 800
rect 42246 0 42302 800
rect 42338 0 42394 800
rect 42430 0 42486 800
rect 42522 0 42578 800
rect 42614 0 42670 800
rect 42706 0 42762 800
rect 42798 0 42854 800
rect 42890 0 42946 800
rect 42982 0 43038 800
rect 43074 0 43130 800
rect 43166 0 43222 800
rect 43258 0 43314 800
rect 43350 0 43406 800
rect 43442 0 43498 800
rect 43534 0 43590 800
rect 43626 0 43682 800
rect 43718 0 43774 800
rect 43810 0 43866 800
rect 43902 0 43958 800
rect 43994 0 44050 800
rect 44086 0 44142 800
rect 44178 0 44234 800
rect 44270 0 44326 800
rect 44362 0 44418 800
rect 44454 0 44510 800
rect 44546 0 44602 800
rect 44638 0 44694 800
rect 44730 0 44786 800
rect 44822 0 44878 800
rect 44914 0 44970 800
rect 45006 0 45062 800
rect 45098 0 45154 800
rect 45190 0 45246 800
rect 45282 0 45338 800
rect 45374 0 45430 800
rect 45466 0 45522 800
rect 45558 0 45614 800
rect 45650 0 45706 800
rect 45742 0 45798 800
rect 45834 0 45890 800
rect 45926 0 45982 800
rect 46018 0 46074 800
rect 46110 0 46166 800
rect 46202 0 46258 800
rect 46294 0 46350 800
rect 46386 0 46442 800
rect 46478 0 46534 800
rect 46570 0 46626 800
rect 46662 0 46718 800
rect 46754 0 46810 800
rect 46846 0 46902 800
rect 46938 0 46994 800
rect 47030 0 47086 800
rect 47122 0 47178 800
rect 47214 0 47270 800
rect 47306 0 47362 800
rect 47398 0 47454 800
<< via2 >>
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 9494 46552 9550 46608
rect 5078 46416 5134 46472
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 10598 45872 10654 45928
rect 15014 46280 15070 46336
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 20350 46144 20406 46200
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 22282 46436 22338 46472
rect 22282 46416 22284 46436
rect 22284 46416 22336 46436
rect 22336 46416 22338 46436
rect 22466 46416 22522 46472
rect 22282 45908 22284 45928
rect 22284 45908 22336 45928
rect 22336 45908 22338 45928
rect 22282 45872 22338 45908
rect 22190 45736 22246 45792
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 22650 46688 22706 46744
rect 23018 46688 23074 46744
rect 22926 46552 22982 46608
rect 22926 46008 22982 46064
rect 23386 46280 23442 46336
rect 23294 46144 23350 46200
rect 24306 46280 24362 46336
rect 24766 46416 24822 46472
rect 24858 45620 24914 45656
rect 24858 45600 24860 45620
rect 24860 45600 24912 45620
rect 24912 45600 24914 45620
rect 26054 45620 26110 45656
rect 26054 45600 26056 45620
rect 26056 45600 26108 45620
rect 26108 45600 26110 45620
rect 27710 46144 27766 46200
rect 28814 46280 28870 46336
rect 28906 46144 28962 46200
rect 28998 46008 29054 46064
rect 28262 45600 28318 45656
rect 28906 45600 28962 45656
rect 29274 46708 29330 46744
rect 29274 46688 29276 46708
rect 29276 46688 29328 46708
rect 29328 46688 29330 46708
rect 30010 46008 30066 46064
rect 30746 46552 30802 46608
rect 30654 46008 30710 46064
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 30838 46008 30894 46064
rect 31666 46416 31722 46472
rect 33414 46552 33470 46608
rect 33138 46452 33140 46472
rect 33140 46452 33192 46472
rect 33192 46452 33194 46472
rect 33138 46416 33194 46452
rect 32862 46280 32918 46336
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34794 46688 34850 46744
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34978 45908 34980 45928
rect 34980 45908 35032 45928
rect 35032 45908 35034 45928
rect 34978 45872 35034 45908
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 35622 46824 35678 46880
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 37554 45736 37610 45792
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 38014 46008 38070 46064
rect 38382 46416 38438 46472
rect 39118 46552 39174 46608
rect 40130 46688 40186 46744
rect 40682 46824 40738 46880
rect 42982 45872 43038 45928
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 18970 2796 18972 2816
rect 18972 2796 19024 2816
rect 19024 2796 19026 2816
rect 18970 2760 19026 2796
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 22282 2760 22338 2816
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
<< metal3 >>
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 34930 47360 35246 47361
rect 34930 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35246 47360
rect 34930 47295 35246 47296
rect 35617 46882 35683 46885
rect 40677 46882 40743 46885
rect 35617 46880 40743 46882
rect 35617 46824 35622 46880
rect 35678 46824 40682 46880
rect 40738 46824 40743 46880
rect 35617 46822 40743 46824
rect 35617 46819 35683 46822
rect 40677 46819 40743 46822
rect 19570 46816 19886 46817
rect 19570 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19886 46816
rect 19570 46751 19886 46752
rect 22645 46746 22711 46749
rect 23013 46746 23079 46749
rect 29269 46746 29335 46749
rect 22050 46744 29335 46746
rect 22050 46688 22650 46744
rect 22706 46688 23018 46744
rect 23074 46688 29274 46744
rect 29330 46688 29335 46744
rect 22050 46686 29335 46688
rect 9489 46610 9555 46613
rect 22050 46610 22110 46686
rect 22645 46683 22711 46686
rect 23013 46683 23079 46686
rect 29269 46683 29335 46686
rect 34789 46746 34855 46749
rect 40125 46746 40191 46749
rect 34789 46744 40191 46746
rect 34789 46688 34794 46744
rect 34850 46688 40130 46744
rect 40186 46688 40191 46744
rect 34789 46686 40191 46688
rect 34789 46683 34855 46686
rect 40125 46683 40191 46686
rect 9489 46608 22110 46610
rect 9489 46552 9494 46608
rect 9550 46552 22110 46608
rect 9489 46550 22110 46552
rect 22921 46610 22987 46613
rect 30741 46610 30807 46613
rect 22921 46608 30807 46610
rect 22921 46552 22926 46608
rect 22982 46552 30746 46608
rect 30802 46552 30807 46608
rect 22921 46550 30807 46552
rect 9489 46547 9555 46550
rect 22921 46547 22987 46550
rect 30741 46547 30807 46550
rect 33409 46610 33475 46613
rect 39113 46610 39179 46613
rect 33409 46608 39179 46610
rect 33409 46552 33414 46608
rect 33470 46552 39118 46608
rect 39174 46552 39179 46608
rect 33409 46550 39179 46552
rect 33409 46547 33475 46550
rect 39113 46547 39179 46550
rect 5073 46474 5139 46477
rect 22277 46474 22343 46477
rect 5073 46472 22343 46474
rect 5073 46416 5078 46472
rect 5134 46416 22282 46472
rect 22338 46416 22343 46472
rect 5073 46414 22343 46416
rect 5073 46411 5139 46414
rect 22277 46411 22343 46414
rect 22461 46474 22527 46477
rect 24761 46474 24827 46477
rect 22461 46472 24827 46474
rect 22461 46416 22466 46472
rect 22522 46416 24766 46472
rect 24822 46416 24827 46472
rect 22461 46414 24827 46416
rect 22461 46411 22527 46414
rect 24761 46411 24827 46414
rect 31661 46474 31727 46477
rect 33133 46474 33199 46477
rect 38377 46474 38443 46477
rect 31661 46472 33199 46474
rect 31661 46416 31666 46472
rect 31722 46416 33138 46472
rect 33194 46416 33199 46472
rect 31661 46414 33199 46416
rect 31661 46411 31727 46414
rect 33133 46411 33199 46414
rect 33366 46472 38443 46474
rect 33366 46416 38382 46472
rect 38438 46416 38443 46472
rect 33366 46414 38443 46416
rect 15009 46338 15075 46341
rect 23381 46338 23447 46341
rect 15009 46336 23447 46338
rect 15009 46280 15014 46336
rect 15070 46280 23386 46336
rect 23442 46280 23447 46336
rect 15009 46278 23447 46280
rect 15009 46275 15075 46278
rect 23381 46275 23447 46278
rect 24301 46338 24367 46341
rect 28809 46338 28875 46341
rect 24301 46336 28875 46338
rect 24301 46280 24306 46336
rect 24362 46280 28814 46336
rect 28870 46280 28875 46336
rect 24301 46278 28875 46280
rect 24301 46275 24367 46278
rect 28809 46275 28875 46278
rect 32857 46338 32923 46341
rect 33366 46338 33426 46414
rect 38377 46411 38443 46414
rect 32857 46336 33426 46338
rect 32857 46280 32862 46336
rect 32918 46280 33426 46336
rect 32857 46278 33426 46280
rect 32857 46275 32923 46278
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 34930 46272 35246 46273
rect 34930 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35246 46272
rect 34930 46207 35246 46208
rect 20345 46202 20411 46205
rect 23289 46202 23355 46205
rect 20345 46200 23355 46202
rect 20345 46144 20350 46200
rect 20406 46144 23294 46200
rect 23350 46144 23355 46200
rect 20345 46142 23355 46144
rect 20345 46139 20411 46142
rect 23289 46139 23355 46142
rect 27705 46202 27771 46205
rect 28901 46202 28967 46205
rect 27705 46200 28967 46202
rect 27705 46144 27710 46200
rect 27766 46144 28906 46200
rect 28962 46144 28967 46200
rect 27705 46142 28967 46144
rect 27705 46139 27771 46142
rect 28901 46139 28967 46142
rect 22921 46066 22987 46069
rect 28993 46066 29059 46069
rect 30005 46066 30071 46069
rect 30649 46066 30715 46069
rect 22921 46064 30715 46066
rect 22921 46008 22926 46064
rect 22982 46008 28998 46064
rect 29054 46008 30010 46064
rect 30066 46008 30654 46064
rect 30710 46008 30715 46064
rect 22921 46006 30715 46008
rect 22921 46003 22987 46006
rect 28993 46003 29059 46006
rect 30005 46003 30071 46006
rect 30649 46003 30715 46006
rect 30833 46066 30899 46069
rect 38009 46066 38075 46069
rect 30833 46064 38075 46066
rect 30833 46008 30838 46064
rect 30894 46008 38014 46064
rect 38070 46008 38075 46064
rect 30833 46006 38075 46008
rect 30833 46003 30899 46006
rect 38009 46003 38075 46006
rect 10593 45930 10659 45933
rect 22277 45930 22343 45933
rect 10593 45928 22343 45930
rect 10593 45872 10598 45928
rect 10654 45872 22282 45928
rect 22338 45872 22343 45928
rect 10593 45870 22343 45872
rect 10593 45867 10659 45870
rect 22277 45867 22343 45870
rect 34973 45930 35039 45933
rect 42977 45930 43043 45933
rect 34973 45928 43043 45930
rect 34973 45872 34978 45928
rect 35034 45872 42982 45928
rect 43038 45872 43043 45928
rect 34973 45870 43043 45872
rect 34973 45867 35039 45870
rect 42977 45867 43043 45870
rect 22185 45794 22251 45797
rect 37549 45794 37615 45797
rect 22185 45792 37615 45794
rect 22185 45736 22190 45792
rect 22246 45736 37554 45792
rect 37610 45736 37615 45792
rect 22185 45734 37615 45736
rect 22185 45731 22251 45734
rect 37549 45731 37615 45734
rect 19570 45728 19886 45729
rect 19570 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19886 45728
rect 19570 45663 19886 45664
rect 24853 45658 24919 45661
rect 26049 45658 26115 45661
rect 24853 45656 26115 45658
rect 24853 45600 24858 45656
rect 24914 45600 26054 45656
rect 26110 45600 26115 45656
rect 24853 45598 26115 45600
rect 24853 45595 24919 45598
rect 26049 45595 26115 45598
rect 28257 45658 28323 45661
rect 28901 45658 28967 45661
rect 28257 45656 28967 45658
rect 28257 45600 28262 45656
rect 28318 45600 28906 45656
rect 28962 45600 28967 45656
rect 28257 45598 28967 45600
rect 28257 45595 28323 45598
rect 28901 45595 28967 45598
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 34930 45119 35246 45120
rect 19570 44640 19886 44641
rect 19570 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19886 44640
rect 19570 44575 19886 44576
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 34930 44031 35246 44032
rect 19570 43552 19886 43553
rect 19570 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19886 43552
rect 19570 43487 19886 43488
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 34930 42943 35246 42944
rect 19570 42464 19886 42465
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 34930 40767 35246 40768
rect 19570 40288 19886 40289
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 18965 2818 19031 2821
rect 22277 2818 22343 2821
rect 18965 2816 22343 2818
rect 18965 2760 18970 2816
rect 19026 2760 22282 2816
rect 22338 2760 22343 2816
rect 18965 2758 22343 2760
rect 18965 2755 19031 2758
rect 22277 2755 22343 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
<< via3 >>
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 47360 4528 47376
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 46816 19888 47376
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 47360 35248 47376
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__157__A dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 18676 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__158__A
timestamp 1666199351
transform -1 0 19780 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__159__A
timestamp 1666199351
transform -1 0 27324 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__170__A
timestamp 1666199351
transform 1 0 25760 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__181__A
timestamp 1666199351
transform 1 0 20424 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__192__A
timestamp 1666199351
transform 1 0 19412 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__193__A_N
timestamp 1666199351
transform 1 0 31372 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__193__B
timestamp 1666199351
transform 1 0 30360 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__194__A1
timestamp 1666199351
transform -1 0 32476 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__194__A2
timestamp 1666199351
transform -1 0 36708 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__194__A3
timestamp 1666199351
transform -1 0 29900 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__195__A
timestamp 1666199351
transform 1 0 29624 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__196__A
timestamp 1666199351
transform -1 0 22172 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__197__A1
timestamp 1666199351
transform 1 0 29900 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__197__A2
timestamp 1666199351
transform -1 0 31004 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__198__A
timestamp 1666199351
transform 1 0 30268 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__199__A
timestamp 1666199351
transform 1 0 25392 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__200__A_N
timestamp 1666199351
transform 1 0 28428 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__200__C
timestamp 1666199351
transform 1 0 28796 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__201__A1
timestamp 1666199351
transform 1 0 28980 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__201__B1_N
timestamp 1666199351
transform 1 0 28520 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__202__B1
timestamp 1666199351
transform 1 0 27784 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__203__A
timestamp 1666199351
transform 1 0 24012 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__203__B_N
timestamp 1666199351
transform 1 0 26496 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__204__A
timestamp 1666199351
transform 1 0 29072 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__206__A
timestamp 1666199351
transform 1 0 22356 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__207__A
timestamp 1666199351
transform 1 0 25024 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__209__A1
timestamp 1666199351
transform -1 0 28704 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__211__B1
timestamp 1666199351
transform -1 0 24196 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__213__A_N
timestamp 1666199351
transform 1 0 41676 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__213__B
timestamp 1666199351
transform 1 0 40020 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__214__A1
timestamp 1666199351
transform -1 0 41308 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__214__A2
timestamp 1666199351
transform 1 0 38548 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__214__A3
timestamp 1666199351
transform 1 0 41860 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__215__A
timestamp 1666199351
transform 1 0 42596 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__216__A
timestamp 1666199351
transform -1 0 32476 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__217__A1
timestamp 1666199351
transform 1 0 39560 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__217__A2
timestamp 1666199351
transform 1 0 39008 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__218__A
timestamp 1666199351
transform 1 0 40572 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__219__A
timestamp 1666199351
transform 1 0 32844 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__220__A_N
timestamp 1666199351
transform 1 0 37444 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__220__C
timestamp 1666199351
transform 1 0 37904 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__221__A1
timestamp 1666199351
transform 1 0 39008 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__221__B1_N
timestamp 1666199351
transform 1 0 38456 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__222__B1
timestamp 1666199351
transform -1 0 36616 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__223__A
timestamp 1666199351
transform -1 0 34592 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__223__B_N
timestamp 1666199351
transform -1 0 36156 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__224__A
timestamp 1666199351
transform 1 0 36800 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__226__A
timestamp 1666199351
transform 1 0 34224 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__227__A
timestamp 1666199351
transform -1 0 32660 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__229__A1
timestamp 1666199351
transform -1 0 43332 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__231__B1
timestamp 1666199351
transform -1 0 33120 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__235__B1
timestamp 1666199351
transform -1 0 23092 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__236__A
timestamp 1666199351
transform 1 0 33028 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__237__A1_N
timestamp 1666199351
transform 1 0 29348 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__237__A2_N
timestamp 1666199351
transform -1 0 23092 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__237__B2
timestamp 1666199351
transform -1 0 27048 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__238__A1
timestamp 1666199351
transform -1 0 26312 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__238__A2
timestamp 1666199351
transform -1 0 25484 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__239__A1
timestamp 1666199351
transform -1 0 24104 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__239__A2
timestamp 1666199351
transform -1 0 25760 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__239__A3
timestamp 1666199351
transform 1 0 23920 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__240__A
timestamp 1666199351
transform 1 0 35420 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__241__A1_N
timestamp 1666199351
transform 1 0 39008 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__241__A2_N
timestamp 1666199351
transform -1 0 37536 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__241__B2
timestamp 1666199351
transform 1 0 40204 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__242__A1
timestamp 1666199351
transform 1 0 40112 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__242__A2
timestamp 1666199351
transform -1 0 35880 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__243__A1
timestamp 1666199351
transform -1 0 42136 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__243__A2
timestamp 1666199351
transform 1 0 38456 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__243__A3
timestamp 1666199351
transform -1 0 33672 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__244__A
timestamp 1666199351
transform 1 0 17480 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__246__A
timestamp 1666199351
transform 1 0 18768 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__251__A1
timestamp 1666199351
transform -1 0 31004 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__251__A2
timestamp 1666199351
transform 1 0 31464 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__251__B1
timestamp 1666199351
transform -1 0 30452 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__252__A1
timestamp 1666199351
transform 1 0 29716 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__252__A2
timestamp 1666199351
transform 1 0 30452 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__253__A1
timestamp 1666199351
transform 1 0 34868 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__256__A1
timestamp 1666199351
transform -1 0 42780 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__256__A2
timestamp 1666199351
transform 1 0 43700 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__256__B1
timestamp 1666199351
transform -1 0 44712 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__257__A1
timestamp 1666199351
transform -1 0 36708 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__257__A2
timestamp 1666199351
transform 1 0 40756 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__258__A1
timestamp 1666199351
transform 1 0 40664 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__259__A
timestamp 1666199351
transform -1 0 17020 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__261__A
timestamp 1666199351
transform 1 0 21160 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__264__A1
timestamp 1666199351
transform 1 0 27692 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__264__A2
timestamp 1666199351
transform 1 0 27048 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__264__B1
timestamp 1666199351
transform -1 0 27324 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__265__A
timestamp 1666199351
transform -1 0 28796 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__265__B
timestamp 1666199351
transform -1 0 28152 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__266__A
timestamp 1666199351
transform 1 0 26036 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__268__B1
timestamp 1666199351
transform 1 0 25944 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__269__A1
timestamp 1666199351
transform 1 0 26496 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__270__A1
timestamp 1666199351
transform 1 0 41308 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__270__A2
timestamp 1666199351
transform -1 0 40204 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__270__B1
timestamp 1666199351
transform -1 0 36432 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__271__A
timestamp 1666199351
transform -1 0 36064 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__271__B
timestamp 1666199351
transform 1 0 35328 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__272__A
timestamp 1666199351
transform -1 0 33948 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__274__B1
timestamp 1666199351
transform -1 0 35144 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__275__A1
timestamp 1666199351
transform 1 0 34868 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__276__A
timestamp 1666199351
transform -1 0 20424 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__278__A
timestamp 1666199351
transform 1 0 21804 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__284__A
timestamp 1666199351
transform -1 0 20792 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__285__A1
timestamp 1666199351
transform -1 0 23460 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__285__A2
timestamp 1666199351
transform 1 0 29624 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__285__B1
timestamp 1666199351
transform -1 0 26312 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__286__A1
timestamp 1666199351
transform 1 0 30912 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__286__A2
timestamp 1666199351
transform 1 0 31924 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__291__A1
timestamp 1666199351
transform 1 0 39652 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__291__A2
timestamp 1666199351
transform 1 0 40572 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__291__B1
timestamp 1666199351
transform -1 0 39284 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__292__A1
timestamp 1666199351
transform -1 0 37260 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__292__A2
timestamp 1666199351
transform -1 0 38180 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__295__A1
timestamp 1666199351
transform 1 0 23368 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__295__C1
timestamp 1666199351
transform 1 0 22816 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 1380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 2208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19
timestamp 1666199351
transform 1 0 2852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40
timestamp 1666199351
transform 1 0 4784 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47
timestamp 1666199351
transform 1 0 5428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1666199351
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57
timestamp 1666199351
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68
timestamp 1666199351
transform 1 0 7360 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75
timestamp 1666199351
transform 1 0 8004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1666199351
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85
timestamp 1666199351
transform 1 0 8924 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_96
timestamp 1666199351
transform 1 0 9936 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_103
timestamp 1666199351
transform 1 0 10580 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1666199351
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_113
timestamp 1666199351
transform 1 0 11500 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_124
timestamp 1666199351
transform 1 0 12512 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_131
timestamp 1666199351
transform 1 0 13156 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1666199351
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_141
timestamp 1666199351
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_152
timestamp 1666199351
transform 1 0 15088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_159
timestamp 1666199351
transform 1 0 15732 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1666199351
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_169
timestamp 1666199351
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_180
timestamp 1666199351
transform 1 0 17664 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_187
timestamp 1666199351
transform 1 0 18308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1666199351
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1666199351
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_202
timestamp 1666199351
transform 1 0 19688 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_209
timestamp 1666199351
transform 1 0 20332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1666199351
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_225
timestamp 1666199351
transform 1 0 21804 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_240
timestamp 1666199351
transform 1 0 23184 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_246 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 23736 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1666199351
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1666199351
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_264
timestamp 1666199351
transform 1 0 25392 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_275
timestamp 1666199351
transform 1 0 26404 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_279
timestamp 1666199351
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1666199351
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_292
timestamp 1666199351
transform 1 0 27968 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_299
timestamp 1666199351
transform 1 0 28612 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_306
timestamp 1666199351
transform 1 0 29256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1666199351
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_314
timestamp 1666199351
transform 1 0 29992 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_321
timestamp 1666199351
transform 1 0 30636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_328
timestamp 1666199351
transform 1 0 31280 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1666199351
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_342
timestamp 1666199351
transform 1 0 32568 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_349
timestamp 1666199351
transform 1 0 33212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_356
timestamp 1666199351
transform 1 0 33856 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1666199351
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_370
timestamp 1666199351
transform 1 0 35144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_377
timestamp 1666199351
transform 1 0 35788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_384
timestamp 1666199351
transform 1 0 36432 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1666199351
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_398
timestamp 1666199351
transform 1 0 37720 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_405
timestamp 1666199351
transform 1 0 38364 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_412
timestamp 1666199351
transform 1 0 39008 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_421
timestamp 1666199351
transform 1 0 39836 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_426
timestamp 1666199351
transform 1 0 40296 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_433
timestamp 1666199351
transform 1 0 40940 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_440
timestamp 1666199351
transform 1 0 41584 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_449
timestamp 1666199351
transform 1 0 42412 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_454
timestamp 1666199351
transform 1 0 42872 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_461
timestamp 1666199351
transform 1 0 43516 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_468
timestamp 1666199351
transform 1 0 44160 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_477
timestamp 1666199351
transform 1 0 44988 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_482
timestamp 1666199351
transform 1 0 45448 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_489
timestamp 1666199351
transform 1 0 46092 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_496
timestamp 1666199351
transform 1 0 46736 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_505
timestamp 1666199351
transform 1 0 47564 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_510
timestamp 1666199351
transform 1 0 48024 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_15
timestamp 1666199351
transform 1 0 2484 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_19
timestamp 1666199351
transform 1 0 2852 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_26
timestamp 1666199351
transform 1 0 3496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_33
timestamp 1666199351
transform 1 0 4140 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_40
timestamp 1666199351
transform 1 0 4784 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_47
timestamp 1666199351
transform 1 0 5428 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1666199351
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_57
timestamp 1666199351
transform 1 0 6348 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_68
timestamp 1666199351
transform 1 0 7360 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_75
timestamp 1666199351
transform 1 0 8004 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_82
timestamp 1666199351
transform 1 0 8648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_89
timestamp 1666199351
transform 1 0 9292 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_96
timestamp 1666199351
transform 1 0 9936 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_103
timestamp 1666199351
transform 1 0 10580 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1666199351
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_113
timestamp 1666199351
transform 1 0 11500 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_124
timestamp 1666199351
transform 1 0 12512 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_131
timestamp 1666199351
transform 1 0 13156 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_138
timestamp 1666199351
transform 1 0 13800 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_145
timestamp 1666199351
transform 1 0 14444 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_152
timestamp 1666199351
transform 1 0 15088 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_159
timestamp 1666199351
transform 1 0 15732 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1666199351
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1666199351
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_174
timestamp 1666199351
transform 1 0 17112 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_181
timestamp 1666199351
transform 1 0 17756 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_188
timestamp 1666199351
transform 1 0 18400 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_195
timestamp 1666199351
transform 1 0 19044 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_202
timestamp 1666199351
transform 1 0 19688 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_209
timestamp 1666199351
transform 1 0 20332 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1666199351
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_225
timestamp 1666199351
transform 1 0 21804 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_232
timestamp 1666199351
transform 1 0 22448 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_245
timestamp 1666199351
transform 1 0 23644 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_258
timestamp 1666199351
transform 1 0 24840 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1666199351
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1666199351
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_281
timestamp 1666199351
transform 1 0 26956 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_292
timestamp 1666199351
transform 1 0 27968 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_305
timestamp 1666199351
transform 1 0 29164 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_318
timestamp 1666199351
transform 1 0 30360 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_325
timestamp 1666199351
transform 1 0 31004 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_332
timestamp 1666199351
transform 1 0 31648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp 1666199351
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_342
timestamp 1666199351
transform 1 0 32568 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_349
timestamp 1666199351
transform 1 0 33212 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_356
timestamp 1666199351
transform 1 0 33856 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_363
timestamp 1666199351
transform 1 0 34500 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_370
timestamp 1666199351
transform 1 0 35144 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_377
timestamp 1666199351
transform 1 0 35788 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_384
timestamp 1666199351
transform 1 0 36432 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_393
timestamp 1666199351
transform 1 0 37260 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_398
timestamp 1666199351
transform 1 0 37720 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_405
timestamp 1666199351
transform 1 0 38364 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_412
timestamp 1666199351
transform 1 0 39008 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_419
timestamp 1666199351
transform 1 0 39652 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_426
timestamp 1666199351
transform 1 0 40296 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_433
timestamp 1666199351
transform 1 0 40940 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_440
timestamp 1666199351
transform 1 0 41584 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_449
timestamp 1666199351
transform 1 0 42412 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_454
timestamp 1666199351
transform 1 0 42872 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_461
timestamp 1666199351
transform 1 0 43516 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_468
timestamp 1666199351
transform 1 0 44160 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_475
timestamp 1666199351
transform 1 0 44804 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_482
timestamp 1666199351
transform 1 0 45448 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_489
timestamp 1666199351
transform 1 0 46092 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_496
timestamp 1666199351
transform 1 0 46736 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_505
timestamp 1666199351
transform 1 0 47564 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_510
timestamp 1666199351
transform 1 0 48024 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1666199351
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1666199351
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1666199351
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_29 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_35
timestamp 1666199351
transform 1 0 4324 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_41
timestamp 1666199351
transform 1 0 4876 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_45
timestamp 1666199351
transform 1 0 5244 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_54
timestamp 1666199351
transform 1 0 6072 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_63
timestamp 1666199351
transform 1 0 6900 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_72
timestamp 1666199351
transform 1 0 7728 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_2_81
timestamp 1666199351
transform 1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1666199351
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_90
timestamp 1666199351
transform 1 0 9384 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_99
timestamp 1666199351
transform 1 0 10212 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_108
timestamp 1666199351
transform 1 0 11040 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_112
timestamp 1666199351
transform 1 0 11408 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_116
timestamp 1666199351
transform 1 0 11776 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_123
timestamp 1666199351
transform 1 0 12420 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_130
timestamp 1666199351
transform 1 0 13064 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_137
timestamp 1666199351
transform 1 0 13708 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_141
timestamp 1666199351
transform 1 0 14076 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_152
timestamp 1666199351
transform 1 0 15088 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_159
timestamp 1666199351
transform 1 0 15732 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_166
timestamp 1666199351
transform 1 0 16376 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_173
timestamp 1666199351
transform 1 0 17020 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_180
timestamp 1666199351
transform 1 0 17664 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_187
timestamp 1666199351
transform 1 0 18308 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1666199351
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_197
timestamp 1666199351
transform 1 0 19228 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_206
timestamp 1666199351
transform 1 0 20056 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_213
timestamp 1666199351
transform 1 0 20700 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_226
timestamp 1666199351
transform 1 0 21896 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_232
timestamp 1666199351
transform 1 0 22448 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_236
timestamp 1666199351
transform 1 0 22816 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_243
timestamp 1666199351
transform 1 0 23460 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1666199351
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_253
timestamp 1666199351
transform 1 0 24380 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_270
timestamp 1666199351
transform 1 0 25944 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_278
timestamp 1666199351
transform 1 0 26680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_282
timestamp 1666199351
transform 1 0 27048 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_288
timestamp 1666199351
transform 1 0 27600 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_298
timestamp 1666199351
transform 1 0 28520 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_305
timestamp 1666199351
transform 1 0 29164 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_309
timestamp 1666199351
transform 1 0 29532 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_314
timestamp 1666199351
transform 1 0 29992 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_321
timestamp 1666199351
transform 1 0 30636 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_328
timestamp 1666199351
transform 1 0 31280 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_335
timestamp 1666199351
transform 1 0 31924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_342
timestamp 1666199351
transform 1 0 32568 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_349
timestamp 1666199351
transform 1 0 33212 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_356
timestamp 1666199351
transform 1 0 33856 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_365
timestamp 1666199351
transform 1 0 34684 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_370
timestamp 1666199351
transform 1 0 35144 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_377
timestamp 1666199351
transform 1 0 35788 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_384
timestamp 1666199351
transform 1 0 36432 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_391
timestamp 1666199351
transform 1 0 37076 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_398
timestamp 1666199351
transform 1 0 37720 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_405
timestamp 1666199351
transform 1 0 38364 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_412
timestamp 1666199351
transform 1 0 39008 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_421
timestamp 1666199351
transform 1 0 39836 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_426
timestamp 1666199351
transform 1 0 40296 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_433
timestamp 1666199351
transform 1 0 40940 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_440
timestamp 1666199351
transform 1 0 41584 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_447
timestamp 1666199351
transform 1 0 42228 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_451
timestamp 1666199351
transform 1 0 42596 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_455
timestamp 1666199351
transform 1 0 42964 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_462
timestamp 1666199351
transform 1 0 43608 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_474
timestamp 1666199351
transform 1 0 44712 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_477
timestamp 1666199351
transform 1 0 44988 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_482
timestamp 1666199351
transform 1 0 45448 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_489
timestamp 1666199351
transform 1 0 46092 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_496
timestamp 1666199351
transform 1 0 46736 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_503
timestamp 1666199351
transform 1 0 47380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_510
timestamp 1666199351
transform 1 0 48024 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1666199351
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1666199351
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1666199351
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1666199351
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1666199351
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1666199351
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1666199351
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1666199351
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1666199351
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1666199351
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1666199351
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1666199351
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1666199351
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1666199351
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1666199351
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_152
timestamp 1666199351
transform 1 0 15088 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_160
timestamp 1666199351
transform 1 0 15824 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_164
timestamp 1666199351
transform 1 0 16192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_169
timestamp 1666199351
transform 1 0 16652 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_180
timestamp 1666199351
transform 1 0 17664 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_187
timestamp 1666199351
transform 1 0 18308 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_194
timestamp 1666199351
transform 1 0 18952 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_201
timestamp 1666199351
transform 1 0 19596 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_208
timestamp 1666199351
transform 1 0 20240 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_215
timestamp 1666199351
transform 1 0 20884 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1666199351
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_225
timestamp 1666199351
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_237
timestamp 1666199351
transform 1 0 22908 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_246
timestamp 1666199351
transform 1 0 23736 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_259
timestamp 1666199351
transform 1 0 24932 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_268
timestamp 1666199351
transform 1 0 25760 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_274
timestamp 1666199351
transform 1 0 26312 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_278
timestamp 1666199351
transform 1 0 26680 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_281
timestamp 1666199351
transform 1 0 26956 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_292
timestamp 1666199351
transform 1 0 27968 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_296
timestamp 1666199351
transform 1 0 28336 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_306
timestamp 1666199351
transform 1 0 29256 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_313
timestamp 1666199351
transform 1 0 29900 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_320
timestamp 1666199351
transform 1 0 30544 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_332
timestamp 1666199351
transform 1 0 31648 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1666199351
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1666199351
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1666199351
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1666199351
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1666199351
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1666199351
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1666199351
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1666199351
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1666199351
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1666199351
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1666199351
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1666199351
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1666199351
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1666199351
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1666199351
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1666199351
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1666199351
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1666199351
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_505
timestamp 1666199351
transform 1 0 47564 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_513
timestamp 1666199351
transform 1 0 48300 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1666199351
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1666199351
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1666199351
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1666199351
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1666199351
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1666199351
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1666199351
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1666199351
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1666199351
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1666199351
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1666199351
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1666199351
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1666199351
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1666199351
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1666199351
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1666199351
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1666199351
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_165
timestamp 1666199351
transform 1 0 16284 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_169
timestamp 1666199351
transform 1 0 16652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_173
timestamp 1666199351
transform 1 0 17020 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_185
timestamp 1666199351
transform 1 0 18124 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1666199351
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_197
timestamp 1666199351
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_203
timestamp 1666199351
transform 1 0 19780 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_216
timestamp 1666199351
transform 1 0 20976 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_4_231
timestamp 1666199351
transform 1 0 22356 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_237
timestamp 1666199351
transform 1 0 22908 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_247
timestamp 1666199351
transform 1 0 23828 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1666199351
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_253
timestamp 1666199351
transform 1 0 24380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_257
timestamp 1666199351
transform 1 0 24748 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_261
timestamp 1666199351
transform 1 0 25116 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_274
timestamp 1666199351
transform 1 0 26312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_281
timestamp 1666199351
transform 1 0 26956 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_288
timestamp 1666199351
transform 1 0 27600 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_296
timestamp 1666199351
transform 1 0 28336 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_306
timestamp 1666199351
transform 1 0 29256 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1666199351
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1666199351
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1666199351
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1666199351
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1666199351
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1666199351
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1666199351
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1666199351
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1666199351
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1666199351
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1666199351
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1666199351
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1666199351
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1666199351
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1666199351
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1666199351
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1666199351
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1666199351
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1666199351
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1666199351
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1666199351
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_513
timestamp 1666199351
transform 1 0 48300 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1666199351
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1666199351
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1666199351
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1666199351
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1666199351
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1666199351
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1666199351
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1666199351
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1666199351
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1666199351
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1666199351
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1666199351
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1666199351
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1666199351
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1666199351
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1666199351
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1666199351
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1666199351
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1666199351
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1666199351
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_193
timestamp 1666199351
transform 1 0 18860 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_200
timestamp 1666199351
transform 1 0 19504 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_204
timestamp 1666199351
transform 1 0 19872 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_208
timestamp 1666199351
transform 1 0 20240 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_215
timestamp 1666199351
transform 1 0 20884 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_222
timestamp 1666199351
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_225
timestamp 1666199351
transform 1 0 21804 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_229
timestamp 1666199351
transform 1 0 22172 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_233
timestamp 1666199351
transform 1 0 22540 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_246
timestamp 1666199351
transform 1 0 23736 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_252
timestamp 1666199351
transform 1 0 24288 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_262
timestamp 1666199351
transform 1 0 25208 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_271
timestamp 1666199351
transform 1 0 26036 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_278
timestamp 1666199351
transform 1 0 26680 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_281
timestamp 1666199351
transform 1 0 26956 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_292
timestamp 1666199351
transform 1 0 27968 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_305
timestamp 1666199351
transform 1 0 29164 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_312
timestamp 1666199351
transform 1 0 29808 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_324
timestamp 1666199351
transform 1 0 30912 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1666199351
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1666199351
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1666199351
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1666199351
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1666199351
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1666199351
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1666199351
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1666199351
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1666199351
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1666199351
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1666199351
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1666199351
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1666199351
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1666199351
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1666199351
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1666199351
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1666199351
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1666199351
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_505
timestamp 1666199351
transform 1 0 47564 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_513
timestamp 1666199351
transform 1 0 48300 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1666199351
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1666199351
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1666199351
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1666199351
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1666199351
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1666199351
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1666199351
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1666199351
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1666199351
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1666199351
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1666199351
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1666199351
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1666199351
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1666199351
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1666199351
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1666199351
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1666199351
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1666199351
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1666199351
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1666199351
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1666199351
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_197
timestamp 1666199351
transform 1 0 19228 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_201
timestamp 1666199351
transform 1 0 19596 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_208
timestamp 1666199351
transform 1 0 20240 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_216
timestamp 1666199351
transform 1 0 20976 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_220
timestamp 1666199351
transform 1 0 21344 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_227
timestamp 1666199351
transform 1 0 21988 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_240
timestamp 1666199351
transform 1 0 23184 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_246
timestamp 1666199351
transform 1 0 23736 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_250
timestamp 1666199351
transform 1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_253
timestamp 1666199351
transform 1 0 24380 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_262
timestamp 1666199351
transform 1 0 25208 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_275
timestamp 1666199351
transform 1 0 26404 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_282
timestamp 1666199351
transform 1 0 27048 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_289
timestamp 1666199351
transform 1 0 27692 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_296
timestamp 1666199351
transform 1 0 28336 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_303
timestamp 1666199351
transform 1 0 28980 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1666199351
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1666199351
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1666199351
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1666199351
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1666199351
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1666199351
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1666199351
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1666199351
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1666199351
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1666199351
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1666199351
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1666199351
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1666199351
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1666199351
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1666199351
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1666199351
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1666199351
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1666199351
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1666199351
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1666199351
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1666199351
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1666199351
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_513
timestamp 1666199351
transform 1 0 48300 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1666199351
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1666199351
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1666199351
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1666199351
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1666199351
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1666199351
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1666199351
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1666199351
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1666199351
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1666199351
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1666199351
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1666199351
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1666199351
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1666199351
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1666199351
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1666199351
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1666199351
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1666199351
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1666199351
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1666199351
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1666199351
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_205
timestamp 1666199351
transform 1 0 19964 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_209
timestamp 1666199351
transform 1 0 20332 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_212
timestamp 1666199351
transform 1 0 20608 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_225
timestamp 1666199351
transform 1 0 21804 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_229
timestamp 1666199351
transform 1 0 22172 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_233
timestamp 1666199351
transform 1 0 22540 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_240
timestamp 1666199351
transform 1 0 23184 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_244
timestamp 1666199351
transform 1 0 23552 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_248
timestamp 1666199351
transform 1 0 23920 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_261
timestamp 1666199351
transform 1 0 25116 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_267
timestamp 1666199351
transform 1 0 25668 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_277
timestamp 1666199351
transform 1 0 26588 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_281
timestamp 1666199351
transform 1 0 26956 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_285
timestamp 1666199351
transform 1 0 27324 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_297
timestamp 1666199351
transform 1 0 28428 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_309
timestamp 1666199351
transform 1 0 29532 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_321
timestamp 1666199351
transform 1 0 30636 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_333
timestamp 1666199351
transform 1 0 31740 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1666199351
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1666199351
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1666199351
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1666199351
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1666199351
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1666199351
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1666199351
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1666199351
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1666199351
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1666199351
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1666199351
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1666199351
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1666199351
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1666199351
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1666199351
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1666199351
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1666199351
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1666199351
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_505
timestamp 1666199351
transform 1 0 47564 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_513
timestamp 1666199351
transform 1 0 48300 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1666199351
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1666199351
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1666199351
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1666199351
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1666199351
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1666199351
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1666199351
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1666199351
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1666199351
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1666199351
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1666199351
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1666199351
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1666199351
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1666199351
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1666199351
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1666199351
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1666199351
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1666199351
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1666199351
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1666199351
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1666199351
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1666199351
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1666199351
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1666199351
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_233
timestamp 1666199351
transform 1 0 22540 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_240
timestamp 1666199351
transform 1 0 23184 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_253
timestamp 1666199351
transform 1 0 24380 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_264
timestamp 1666199351
transform 1 0 25392 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_270
timestamp 1666199351
transform 1 0 25944 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_282
timestamp 1666199351
transform 1 0 27048 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_294
timestamp 1666199351
transform 1 0 28152 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_306
timestamp 1666199351
transform 1 0 29256 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1666199351
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1666199351
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1666199351
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1666199351
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1666199351
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1666199351
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1666199351
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1666199351
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1666199351
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1666199351
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1666199351
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1666199351
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1666199351
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1666199351
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1666199351
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1666199351
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1666199351
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1666199351
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1666199351
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1666199351
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1666199351
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_513
timestamp 1666199351
transform 1 0 48300 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1666199351
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1666199351
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1666199351
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1666199351
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1666199351
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1666199351
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1666199351
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1666199351
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1666199351
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1666199351
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1666199351
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1666199351
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1666199351
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1666199351
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1666199351
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1666199351
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1666199351
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1666199351
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1666199351
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1666199351
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1666199351
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1666199351
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1666199351
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1666199351
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1666199351
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1666199351
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1666199351
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1666199351
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1666199351
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1666199351
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1666199351
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1666199351
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1666199351
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1666199351
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1666199351
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1666199351
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1666199351
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1666199351
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1666199351
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1666199351
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1666199351
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1666199351
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1666199351
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1666199351
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_417
timestamp 1666199351
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_429
timestamp 1666199351
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1666199351
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1666199351
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1666199351
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1666199351
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1666199351
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1666199351
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1666199351
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1666199351
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_505
timestamp 1666199351
transform 1 0 47564 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_513
timestamp 1666199351
transform 1 0 48300 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1666199351
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1666199351
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1666199351
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1666199351
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1666199351
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1666199351
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1666199351
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1666199351
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1666199351
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1666199351
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1666199351
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1666199351
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1666199351
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1666199351
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1666199351
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1666199351
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1666199351
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1666199351
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1666199351
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1666199351
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1666199351
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1666199351
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1666199351
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1666199351
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1666199351
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1666199351
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1666199351
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1666199351
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1666199351
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1666199351
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1666199351
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1666199351
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1666199351
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1666199351
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1666199351
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1666199351
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1666199351
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1666199351
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1666199351
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1666199351
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1666199351
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1666199351
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_401
timestamp 1666199351
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1666199351
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1666199351
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1666199351
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1666199351
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1666199351
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1666199351
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1666199351
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1666199351
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1666199351
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1666199351
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1666199351
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_513
timestamp 1666199351
transform 1 0 48300 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1666199351
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1666199351
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1666199351
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1666199351
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1666199351
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1666199351
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1666199351
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1666199351
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1666199351
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1666199351
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1666199351
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1666199351
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1666199351
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1666199351
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1666199351
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1666199351
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1666199351
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1666199351
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1666199351
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1666199351
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1666199351
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1666199351
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1666199351
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1666199351
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1666199351
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1666199351
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1666199351
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1666199351
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1666199351
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1666199351
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1666199351
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1666199351
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1666199351
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1666199351
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1666199351
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1666199351
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1666199351
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1666199351
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1666199351
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1666199351
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1666199351
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1666199351
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1666199351
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_405
timestamp 1666199351
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_417
timestamp 1666199351
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_429
timestamp 1666199351
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1666199351
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1666199351
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1666199351
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1666199351
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1666199351
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1666199351
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1666199351
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1666199351
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_505
timestamp 1666199351
transform 1 0 47564 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_513
timestamp 1666199351
transform 1 0 48300 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1666199351
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1666199351
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1666199351
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1666199351
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1666199351
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1666199351
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1666199351
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1666199351
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1666199351
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1666199351
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1666199351
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1666199351
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1666199351
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1666199351
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1666199351
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1666199351
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1666199351
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1666199351
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1666199351
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1666199351
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1666199351
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1666199351
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1666199351
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1666199351
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1666199351
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1666199351
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1666199351
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1666199351
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1666199351
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1666199351
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1666199351
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1666199351
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1666199351
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1666199351
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1666199351
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1666199351
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1666199351
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1666199351
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1666199351
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1666199351
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1666199351
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1666199351
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_401
timestamp 1666199351
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1666199351
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1666199351
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1666199351
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1666199351
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1666199351
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1666199351
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1666199351
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1666199351
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1666199351
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1666199351
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1666199351
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_513
timestamp 1666199351
transform 1 0 48300 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1666199351
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1666199351
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1666199351
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1666199351
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1666199351
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1666199351
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1666199351
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1666199351
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1666199351
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1666199351
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1666199351
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1666199351
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1666199351
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1666199351
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1666199351
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1666199351
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1666199351
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1666199351
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1666199351
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1666199351
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1666199351
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1666199351
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1666199351
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1666199351
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1666199351
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1666199351
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1666199351
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1666199351
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1666199351
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1666199351
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1666199351
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1666199351
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1666199351
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1666199351
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1666199351
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1666199351
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1666199351
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1666199351
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1666199351
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1666199351
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1666199351
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1666199351
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1666199351
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_405
timestamp 1666199351
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_417
timestamp 1666199351
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_429
timestamp 1666199351
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1666199351
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1666199351
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1666199351
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1666199351
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1666199351
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1666199351
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1666199351
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1666199351
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_505
timestamp 1666199351
transform 1 0 47564 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_513
timestamp 1666199351
transform 1 0 48300 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1666199351
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1666199351
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1666199351
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1666199351
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1666199351
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1666199351
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1666199351
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1666199351
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1666199351
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1666199351
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1666199351
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1666199351
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1666199351
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1666199351
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1666199351
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1666199351
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1666199351
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1666199351
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1666199351
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1666199351
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1666199351
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1666199351
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1666199351
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1666199351
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1666199351
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1666199351
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1666199351
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1666199351
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1666199351
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1666199351
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1666199351
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1666199351
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1666199351
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1666199351
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1666199351
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1666199351
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1666199351
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1666199351
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1666199351
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1666199351
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1666199351
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1666199351
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_401
timestamp 1666199351
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1666199351
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1666199351
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1666199351
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1666199351
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_445
timestamp 1666199351
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_457
timestamp 1666199351
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1666199351
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1666199351
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1666199351
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1666199351
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_501
timestamp 1666199351
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_513
timestamp 1666199351
transform 1 0 48300 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1666199351
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1666199351
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1666199351
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1666199351
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1666199351
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1666199351
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1666199351
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1666199351
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1666199351
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1666199351
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1666199351
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1666199351
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1666199351
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1666199351
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1666199351
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1666199351
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1666199351
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1666199351
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1666199351
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1666199351
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1666199351
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1666199351
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1666199351
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1666199351
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1666199351
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1666199351
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1666199351
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1666199351
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1666199351
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1666199351
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1666199351
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1666199351
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1666199351
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1666199351
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1666199351
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1666199351
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1666199351
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1666199351
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1666199351
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1666199351
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1666199351
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1666199351
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1666199351
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_405
timestamp 1666199351
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_417
timestamp 1666199351
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_429
timestamp 1666199351
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1666199351
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1666199351
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1666199351
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1666199351
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1666199351
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1666199351
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1666199351
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1666199351
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_505
timestamp 1666199351
transform 1 0 47564 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_513
timestamp 1666199351
transform 1 0 48300 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1666199351
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1666199351
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1666199351
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1666199351
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1666199351
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1666199351
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1666199351
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1666199351
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1666199351
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1666199351
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1666199351
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1666199351
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1666199351
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1666199351
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1666199351
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1666199351
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1666199351
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1666199351
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1666199351
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1666199351
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1666199351
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1666199351
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1666199351
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1666199351
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1666199351
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1666199351
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1666199351
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1666199351
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1666199351
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1666199351
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1666199351
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1666199351
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1666199351
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1666199351
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1666199351
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1666199351
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1666199351
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1666199351
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1666199351
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1666199351
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1666199351
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1666199351
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_401
timestamp 1666199351
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1666199351
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1666199351
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1666199351
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1666199351
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_445
timestamp 1666199351
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_457
timestamp 1666199351
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1666199351
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1666199351
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1666199351
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_489
timestamp 1666199351
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_501
timestamp 1666199351
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_513
timestamp 1666199351
transform 1 0 48300 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1666199351
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1666199351
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1666199351
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1666199351
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1666199351
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1666199351
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1666199351
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1666199351
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1666199351
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1666199351
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1666199351
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1666199351
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1666199351
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1666199351
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1666199351
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1666199351
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1666199351
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1666199351
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1666199351
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1666199351
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1666199351
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1666199351
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1666199351
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1666199351
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1666199351
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1666199351
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1666199351
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1666199351
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1666199351
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1666199351
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1666199351
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1666199351
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1666199351
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1666199351
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1666199351
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1666199351
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1666199351
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1666199351
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1666199351
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1666199351
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1666199351
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1666199351
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1666199351
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_405
timestamp 1666199351
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_417
timestamp 1666199351
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_429
timestamp 1666199351
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1666199351
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1666199351
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1666199351
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1666199351
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1666199351
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1666199351
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1666199351
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1666199351
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_505
timestamp 1666199351
transform 1 0 47564 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_513
timestamp 1666199351
transform 1 0 48300 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1666199351
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1666199351
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1666199351
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1666199351
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1666199351
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1666199351
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1666199351
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1666199351
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1666199351
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1666199351
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1666199351
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1666199351
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1666199351
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1666199351
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1666199351
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1666199351
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1666199351
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1666199351
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1666199351
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1666199351
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1666199351
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1666199351
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1666199351
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1666199351
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1666199351
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1666199351
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1666199351
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1666199351
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1666199351
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1666199351
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_289
timestamp 1666199351
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1666199351
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1666199351
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1666199351
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1666199351
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1666199351
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1666199351
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1666199351
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1666199351
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1666199351
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1666199351
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1666199351
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_401
timestamp 1666199351
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1666199351
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1666199351
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_421
timestamp 1666199351
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_433
timestamp 1666199351
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_445
timestamp 1666199351
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_457
timestamp 1666199351
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1666199351
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1666199351
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1666199351
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1666199351
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1666199351
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_513
timestamp 1666199351
transform 1 0 48300 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1666199351
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1666199351
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1666199351
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1666199351
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1666199351
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1666199351
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1666199351
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1666199351
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1666199351
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1666199351
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1666199351
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1666199351
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1666199351
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1666199351
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1666199351
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1666199351
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1666199351
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1666199351
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1666199351
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1666199351
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1666199351
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1666199351
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1666199351
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1666199351
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1666199351
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1666199351
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1666199351
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1666199351
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1666199351
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1666199351
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1666199351
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1666199351
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1666199351
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1666199351
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1666199351
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1666199351
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1666199351
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1666199351
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1666199351
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1666199351
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1666199351
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1666199351
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1666199351
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_405
timestamp 1666199351
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_417
timestamp 1666199351
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_429
timestamp 1666199351
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1666199351
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1666199351
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1666199351
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1666199351
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1666199351
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_485
timestamp 1666199351
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1666199351
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1666199351
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_505
timestamp 1666199351
transform 1 0 47564 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_513
timestamp 1666199351
transform 1 0 48300 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1666199351
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1666199351
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1666199351
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1666199351
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1666199351
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1666199351
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1666199351
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1666199351
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1666199351
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1666199351
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1666199351
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1666199351
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1666199351
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1666199351
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1666199351
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1666199351
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1666199351
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1666199351
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1666199351
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1666199351
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1666199351
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1666199351
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1666199351
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1666199351
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1666199351
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1666199351
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1666199351
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1666199351
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1666199351
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1666199351
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_289
timestamp 1666199351
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1666199351
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1666199351
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1666199351
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1666199351
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1666199351
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1666199351
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1666199351
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1666199351
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1666199351
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1666199351
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1666199351
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_401
timestamp 1666199351
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1666199351
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1666199351
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 1666199351
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_433
timestamp 1666199351
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_445
timestamp 1666199351
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_457
timestamp 1666199351
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1666199351
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1666199351
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1666199351
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1666199351
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_501
timestamp 1666199351
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_513
timestamp 1666199351
transform 1 0 48300 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1666199351
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1666199351
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1666199351
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1666199351
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1666199351
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1666199351
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1666199351
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1666199351
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1666199351
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1666199351
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1666199351
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1666199351
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1666199351
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1666199351
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1666199351
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1666199351
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1666199351
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1666199351
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1666199351
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1666199351
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1666199351
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1666199351
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1666199351
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1666199351
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1666199351
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1666199351
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1666199351
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1666199351
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1666199351
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1666199351
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1666199351
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1666199351
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1666199351
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1666199351
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1666199351
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1666199351
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1666199351
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1666199351
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1666199351
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1666199351
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1666199351
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1666199351
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1666199351
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_405
timestamp 1666199351
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_417
timestamp 1666199351
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_429
timestamp 1666199351
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1666199351
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1666199351
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1666199351
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1666199351
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_473
timestamp 1666199351
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_485
timestamp 1666199351
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1666199351
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1666199351
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_505
timestamp 1666199351
transform 1 0 47564 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_513
timestamp 1666199351
transform 1 0 48300 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1666199351
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1666199351
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1666199351
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1666199351
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1666199351
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1666199351
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1666199351
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1666199351
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1666199351
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1666199351
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1666199351
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1666199351
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1666199351
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1666199351
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1666199351
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1666199351
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1666199351
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1666199351
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1666199351
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1666199351
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1666199351
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1666199351
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1666199351
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1666199351
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1666199351
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1666199351
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1666199351
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1666199351
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1666199351
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1666199351
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_289
timestamp 1666199351
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1666199351
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1666199351
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1666199351
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1666199351
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1666199351
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1666199351
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1666199351
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1666199351
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1666199351
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1666199351
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1666199351
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_401
timestamp 1666199351
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1666199351
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1666199351
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_421
timestamp 1666199351
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_433
timestamp 1666199351
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_445
timestamp 1666199351
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_457
timestamp 1666199351
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1666199351
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1666199351
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1666199351
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1666199351
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1666199351
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_513
timestamp 1666199351
transform 1 0 48300 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1666199351
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1666199351
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1666199351
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1666199351
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1666199351
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1666199351
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1666199351
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1666199351
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1666199351
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1666199351
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1666199351
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1666199351
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1666199351
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1666199351
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1666199351
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1666199351
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1666199351
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1666199351
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1666199351
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1666199351
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1666199351
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1666199351
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1666199351
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1666199351
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1666199351
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1666199351
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_249
timestamp 1666199351
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_261
timestamp 1666199351
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1666199351
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1666199351
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1666199351
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1666199351
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1666199351
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1666199351
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1666199351
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1666199351
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1666199351
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1666199351
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1666199351
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1666199351
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1666199351
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1666199351
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1666199351
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_405
timestamp 1666199351
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_417
timestamp 1666199351
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_429
timestamp 1666199351
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1666199351
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1666199351
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1666199351
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1666199351
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1666199351
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 1666199351
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1666199351
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1666199351
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_505
timestamp 1666199351
transform 1 0 47564 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_513
timestamp 1666199351
transform 1 0 48300 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1666199351
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1666199351
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1666199351
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1666199351
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1666199351
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1666199351
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1666199351
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1666199351
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1666199351
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1666199351
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1666199351
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1666199351
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1666199351
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1666199351
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1666199351
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1666199351
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1666199351
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1666199351
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1666199351
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1666199351
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1666199351
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1666199351
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1666199351
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1666199351
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_233
timestamp 1666199351
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1666199351
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1666199351
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1666199351
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1666199351
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1666199351
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1666199351
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1666199351
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1666199351
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1666199351
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1666199351
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1666199351
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1666199351
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1666199351
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1666199351
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1666199351
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1666199351
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1666199351
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_401
timestamp 1666199351
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1666199351
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1666199351
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1666199351
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_433
timestamp 1666199351
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_445
timestamp 1666199351
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_457
timestamp 1666199351
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1666199351
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1666199351
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1666199351
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1666199351
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_501
timestamp 1666199351
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_513
timestamp 1666199351
transform 1 0 48300 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1666199351
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1666199351
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1666199351
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1666199351
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1666199351
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1666199351
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1666199351
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1666199351
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1666199351
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1666199351
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1666199351
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1666199351
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1666199351
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1666199351
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1666199351
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1666199351
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1666199351
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1666199351
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1666199351
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1666199351
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1666199351
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1666199351
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1666199351
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1666199351
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1666199351
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1666199351
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1666199351
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1666199351
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1666199351
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1666199351
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1666199351
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1666199351
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1666199351
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1666199351
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1666199351
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1666199351
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1666199351
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1666199351
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1666199351
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1666199351
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1666199351
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1666199351
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1666199351
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_405
timestamp 1666199351
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_417
timestamp 1666199351
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_429
timestamp 1666199351
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1666199351
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1666199351
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1666199351
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1666199351
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1666199351
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1666199351
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1666199351
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1666199351
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_505
timestamp 1666199351
transform 1 0 47564 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_513
timestamp 1666199351
transform 1 0 48300 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1666199351
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1666199351
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1666199351
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1666199351
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1666199351
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1666199351
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1666199351
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1666199351
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1666199351
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1666199351
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1666199351
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1666199351
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1666199351
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1666199351
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1666199351
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1666199351
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1666199351
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1666199351
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1666199351
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1666199351
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1666199351
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1666199351
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1666199351
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1666199351
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1666199351
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1666199351
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1666199351
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1666199351
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1666199351
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1666199351
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_289
timestamp 1666199351
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1666199351
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1666199351
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1666199351
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1666199351
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1666199351
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1666199351
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1666199351
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1666199351
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1666199351
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1666199351
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1666199351
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_401
timestamp 1666199351
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1666199351
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1666199351
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_421
timestamp 1666199351
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_433
timestamp 1666199351
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_445
timestamp 1666199351
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_457
timestamp 1666199351
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1666199351
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1666199351
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1666199351
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1666199351
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_501
timestamp 1666199351
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_513
timestamp 1666199351
transform 1 0 48300 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1666199351
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1666199351
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1666199351
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1666199351
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1666199351
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1666199351
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1666199351
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1666199351
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1666199351
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1666199351
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1666199351
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1666199351
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1666199351
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1666199351
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1666199351
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1666199351
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1666199351
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1666199351
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1666199351
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1666199351
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1666199351
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1666199351
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1666199351
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1666199351
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1666199351
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1666199351
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1666199351
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_261
timestamp 1666199351
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1666199351
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1666199351
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1666199351
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1666199351
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_305
timestamp 1666199351
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_317
timestamp 1666199351
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1666199351
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1666199351
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1666199351
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1666199351
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1666199351
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1666199351
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1666199351
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1666199351
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1666199351
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_405
timestamp 1666199351
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_417
timestamp 1666199351
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_429
timestamp 1666199351
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1666199351
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1666199351
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1666199351
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_461
timestamp 1666199351
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1666199351
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1666199351
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1666199351
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1666199351
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_505
timestamp 1666199351
transform 1 0 47564 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_513
timestamp 1666199351
transform 1 0 48300 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1666199351
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1666199351
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1666199351
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1666199351
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1666199351
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1666199351
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1666199351
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1666199351
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1666199351
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1666199351
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1666199351
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1666199351
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1666199351
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1666199351
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1666199351
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1666199351
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1666199351
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1666199351
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1666199351
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1666199351
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1666199351
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1666199351
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1666199351
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1666199351
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_233
timestamp 1666199351
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1666199351
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1666199351
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1666199351
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1666199351
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1666199351
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_289
timestamp 1666199351
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1666199351
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1666199351
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1666199351
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1666199351
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1666199351
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1666199351
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1666199351
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1666199351
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1666199351
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1666199351
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1666199351
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_401
timestamp 1666199351
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1666199351
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1666199351
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_421
timestamp 1666199351
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_433
timestamp 1666199351
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_445
timestamp 1666199351
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_457
timestamp 1666199351
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1666199351
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1666199351
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1666199351
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1666199351
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_501
timestamp 1666199351
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_513
timestamp 1666199351
transform 1 0 48300 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1666199351
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1666199351
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1666199351
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1666199351
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1666199351
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1666199351
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1666199351
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1666199351
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1666199351
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1666199351
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1666199351
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1666199351
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1666199351
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1666199351
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1666199351
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1666199351
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1666199351
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1666199351
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1666199351
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1666199351
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1666199351
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1666199351
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1666199351
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1666199351
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1666199351
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1666199351
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_249
timestamp 1666199351
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1666199351
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1666199351
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1666199351
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1666199351
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1666199351
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1666199351
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1666199351
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1666199351
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1666199351
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1666199351
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1666199351
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1666199351
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1666199351
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1666199351
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1666199351
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1666199351
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_405
timestamp 1666199351
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_417
timestamp 1666199351
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_429
timestamp 1666199351
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1666199351
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1666199351
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1666199351
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_461
timestamp 1666199351
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_473
timestamp 1666199351
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_485
timestamp 1666199351
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1666199351
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1666199351
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_505
timestamp 1666199351
transform 1 0 47564 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_513
timestamp 1666199351
transform 1 0 48300 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1666199351
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1666199351
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1666199351
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1666199351
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1666199351
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1666199351
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1666199351
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1666199351
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1666199351
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1666199351
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1666199351
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1666199351
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1666199351
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1666199351
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1666199351
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1666199351
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1666199351
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1666199351
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1666199351
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1666199351
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1666199351
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1666199351
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1666199351
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_221
timestamp 1666199351
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_233
timestamp 1666199351
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1666199351
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1666199351
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1666199351
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1666199351
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1666199351
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_289
timestamp 1666199351
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1666199351
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1666199351
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1666199351
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1666199351
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1666199351
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1666199351
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1666199351
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1666199351
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1666199351
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1666199351
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1666199351
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_401
timestamp 1666199351
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1666199351
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1666199351
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_421
timestamp 1666199351
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_433
timestamp 1666199351
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_445
timestamp 1666199351
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_457
timestamp 1666199351
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1666199351
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1666199351
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1666199351
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1666199351
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_501
timestamp 1666199351
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_513
timestamp 1666199351
transform 1 0 48300 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1666199351
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1666199351
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1666199351
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1666199351
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1666199351
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1666199351
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1666199351
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1666199351
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1666199351
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1666199351
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1666199351
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1666199351
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1666199351
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1666199351
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1666199351
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1666199351
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1666199351
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1666199351
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1666199351
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1666199351
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1666199351
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1666199351
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1666199351
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1666199351
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1666199351
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1666199351
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_249
timestamp 1666199351
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_261
timestamp 1666199351
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1666199351
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1666199351
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1666199351
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1666199351
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1666199351
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1666199351
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1666199351
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1666199351
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1666199351
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1666199351
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1666199351
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1666199351
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1666199351
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1666199351
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1666199351
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_405
timestamp 1666199351
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_417
timestamp 1666199351
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_429
timestamp 1666199351
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1666199351
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1666199351
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_449
timestamp 1666199351
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_461
timestamp 1666199351
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_473
timestamp 1666199351
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_485
timestamp 1666199351
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1666199351
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1666199351
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_505
timestamp 1666199351
transform 1 0 47564 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_513
timestamp 1666199351
transform 1 0 48300 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1666199351
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1666199351
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1666199351
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1666199351
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1666199351
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1666199351
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1666199351
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1666199351
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1666199351
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1666199351
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1666199351
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1666199351
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1666199351
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1666199351
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1666199351
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1666199351
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1666199351
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1666199351
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1666199351
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1666199351
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1666199351
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1666199351
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1666199351
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1666199351
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_233
timestamp 1666199351
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1666199351
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1666199351
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1666199351
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1666199351
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1666199351
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1666199351
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1666199351
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1666199351
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1666199351
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1666199351
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_333
timestamp 1666199351
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1666199351
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1666199351
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1666199351
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1666199351
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1666199351
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1666199351
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_401
timestamp 1666199351
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1666199351
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1666199351
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_421
timestamp 1666199351
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_433
timestamp 1666199351
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_445
timestamp 1666199351
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_457
timestamp 1666199351
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1666199351
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1666199351
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1666199351
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_489
timestamp 1666199351
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_501
timestamp 1666199351
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_513
timestamp 1666199351
transform 1 0 48300 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1666199351
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1666199351
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1666199351
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1666199351
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1666199351
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1666199351
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1666199351
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1666199351
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1666199351
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1666199351
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1666199351
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1666199351
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1666199351
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1666199351
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1666199351
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1666199351
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1666199351
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1666199351
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1666199351
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1666199351
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1666199351
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1666199351
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1666199351
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1666199351
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1666199351
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1666199351
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1666199351
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_261
timestamp 1666199351
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1666199351
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1666199351
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1666199351
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1666199351
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1666199351
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1666199351
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1666199351
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1666199351
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1666199351
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1666199351
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1666199351
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1666199351
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1666199351
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1666199351
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1666199351
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_405
timestamp 1666199351
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_417
timestamp 1666199351
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_429
timestamp 1666199351
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1666199351
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1666199351
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1666199351
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1666199351
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_473
timestamp 1666199351
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_485
timestamp 1666199351
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1666199351
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1666199351
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_505
timestamp 1666199351
transform 1 0 47564 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_513
timestamp 1666199351
transform 1 0 48300 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1666199351
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1666199351
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1666199351
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1666199351
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1666199351
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1666199351
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1666199351
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1666199351
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1666199351
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1666199351
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1666199351
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1666199351
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1666199351
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1666199351
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1666199351
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1666199351
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1666199351
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1666199351
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1666199351
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1666199351
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1666199351
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1666199351
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1666199351
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1666199351
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_233
timestamp 1666199351
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1666199351
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1666199351
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1666199351
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1666199351
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1666199351
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_289
timestamp 1666199351
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1666199351
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1666199351
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1666199351
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1666199351
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1666199351
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1666199351
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1666199351
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1666199351
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1666199351
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1666199351
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1666199351
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_401
timestamp 1666199351
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 1666199351
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1666199351
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_421
timestamp 1666199351
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_433
timestamp 1666199351
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_445
timestamp 1666199351
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_457
timestamp 1666199351
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1666199351
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1666199351
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1666199351
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1666199351
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_501
timestamp 1666199351
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_513
timestamp 1666199351
transform 1 0 48300 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1666199351
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1666199351
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1666199351
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1666199351
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1666199351
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1666199351
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1666199351
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1666199351
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1666199351
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1666199351
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1666199351
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1666199351
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1666199351
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1666199351
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1666199351
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1666199351
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1666199351
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1666199351
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1666199351
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1666199351
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1666199351
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_205
timestamp 1666199351
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1666199351
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1666199351
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1666199351
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1666199351
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 1666199351
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1666199351
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1666199351
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1666199351
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1666199351
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1666199351
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1666199351
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1666199351
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1666199351
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1666199351
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1666199351
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1666199351
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1666199351
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1666199351
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1666199351
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1666199351
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1666199351
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_405
timestamp 1666199351
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_417
timestamp 1666199351
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_429
timestamp 1666199351
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1666199351
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1666199351
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_449
timestamp 1666199351
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_461
timestamp 1666199351
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_473
timestamp 1666199351
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_485
timestamp 1666199351
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1666199351
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1666199351
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_505
timestamp 1666199351
transform 1 0 47564 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_513
timestamp 1666199351
transform 1 0 48300 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1666199351
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1666199351
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1666199351
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1666199351
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1666199351
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1666199351
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1666199351
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1666199351
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1666199351
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1666199351
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1666199351
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1666199351
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1666199351
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1666199351
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1666199351
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1666199351
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1666199351
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1666199351
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1666199351
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1666199351
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1666199351
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1666199351
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1666199351
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1666199351
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1666199351
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1666199351
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1666199351
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1666199351
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1666199351
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1666199351
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1666199351
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1666199351
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1666199351
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1666199351
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1666199351
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1666199351
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1666199351
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1666199351
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1666199351
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1666199351
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1666199351
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1666199351
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_401
timestamp 1666199351
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 1666199351
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1666199351
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_421
timestamp 1666199351
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_433
timestamp 1666199351
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_445
timestamp 1666199351
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_457
timestamp 1666199351
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1666199351
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1666199351
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1666199351
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1666199351
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_501
timestamp 1666199351
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_513
timestamp 1666199351
transform 1 0 48300 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1666199351
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1666199351
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1666199351
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1666199351
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1666199351
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1666199351
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1666199351
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1666199351
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1666199351
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1666199351
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1666199351
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1666199351
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1666199351
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1666199351
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1666199351
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1666199351
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1666199351
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1666199351
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1666199351
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1666199351
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1666199351
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1666199351
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1666199351
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1666199351
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1666199351
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1666199351
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1666199351
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1666199351
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1666199351
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1666199351
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1666199351
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1666199351
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1666199351
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1666199351
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1666199351
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1666199351
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1666199351
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1666199351
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1666199351
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1666199351
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1666199351
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1666199351
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_393
timestamp 1666199351
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_405
timestamp 1666199351
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_417
timestamp 1666199351
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_429
timestamp 1666199351
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 1666199351
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1666199351
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_449
timestamp 1666199351
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_461
timestamp 1666199351
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_473
timestamp 1666199351
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_485
timestamp 1666199351
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1666199351
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1666199351
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_505
timestamp 1666199351
transform 1 0 47564 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_513
timestamp 1666199351
transform 1 0 48300 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1666199351
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1666199351
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1666199351
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1666199351
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1666199351
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1666199351
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1666199351
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1666199351
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1666199351
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1666199351
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1666199351
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1666199351
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1666199351
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1666199351
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1666199351
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1666199351
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1666199351
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1666199351
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1666199351
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1666199351
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1666199351
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1666199351
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1666199351
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1666199351
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_233
timestamp 1666199351
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1666199351
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1666199351
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1666199351
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1666199351
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1666199351
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 1666199351
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1666199351
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1666199351
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1666199351
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1666199351
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1666199351
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1666199351
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1666199351
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1666199351
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1666199351
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1666199351
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1666199351
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_401
timestamp 1666199351
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1666199351
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1666199351
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_421
timestamp 1666199351
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_433
timestamp 1666199351
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_445
timestamp 1666199351
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_457
timestamp 1666199351
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1666199351
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1666199351
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1666199351
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_489
timestamp 1666199351
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_501
timestamp 1666199351
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_513
timestamp 1666199351
transform 1 0 48300 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1666199351
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1666199351
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1666199351
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1666199351
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1666199351
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1666199351
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1666199351
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1666199351
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1666199351
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1666199351
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1666199351
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1666199351
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1666199351
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1666199351
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1666199351
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1666199351
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1666199351
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1666199351
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1666199351
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1666199351
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1666199351
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1666199351
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1666199351
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1666199351
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1666199351
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1666199351
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1666199351
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1666199351
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1666199351
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1666199351
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1666199351
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1666199351
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1666199351
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_317
timestamp 1666199351
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1666199351
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1666199351
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1666199351
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1666199351
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1666199351
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1666199351
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1666199351
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1666199351
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1666199351
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_405
timestamp 1666199351
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_417
timestamp 1666199351
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_429
timestamp 1666199351
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 1666199351
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1666199351
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_449
timestamp 1666199351
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_461
timestamp 1666199351
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_473
timestamp 1666199351
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_485
timestamp 1666199351
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1666199351
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1666199351
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_505
timestamp 1666199351
transform 1 0 47564 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_513
timestamp 1666199351
transform 1 0 48300 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1666199351
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1666199351
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1666199351
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1666199351
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1666199351
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1666199351
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1666199351
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1666199351
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1666199351
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1666199351
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1666199351
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1666199351
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1666199351
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1666199351
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1666199351
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1666199351
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1666199351
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1666199351
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1666199351
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1666199351
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1666199351
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1666199351
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1666199351
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1666199351
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_233
timestamp 1666199351
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1666199351
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1666199351
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1666199351
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1666199351
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1666199351
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1666199351
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1666199351
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1666199351
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1666199351
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1666199351
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1666199351
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_345
timestamp 1666199351
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1666199351
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1666199351
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1666199351
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1666199351
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1666199351
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_401
timestamp 1666199351
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1666199351
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1666199351
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_421
timestamp 1666199351
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_433
timestamp 1666199351
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_445
timestamp 1666199351
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_457
timestamp 1666199351
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 1666199351
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1666199351
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_477
timestamp 1666199351
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_489
timestamp 1666199351
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_501
timestamp 1666199351
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_513
timestamp 1666199351
transform 1 0 48300 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1666199351
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1666199351
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1666199351
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1666199351
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1666199351
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1666199351
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1666199351
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1666199351
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1666199351
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1666199351
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1666199351
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1666199351
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1666199351
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1666199351
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1666199351
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1666199351
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1666199351
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1666199351
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1666199351
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1666199351
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1666199351
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1666199351
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1666199351
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1666199351
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1666199351
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1666199351
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1666199351
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1666199351
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1666199351
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1666199351
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1666199351
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1666199351
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1666199351
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_317
timestamp 1666199351
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1666199351
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1666199351
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1666199351
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1666199351
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1666199351
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1666199351
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1666199351
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1666199351
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1666199351
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_405
timestamp 1666199351
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_417
timestamp 1666199351
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_429
timestamp 1666199351
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 1666199351
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1666199351
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_449
timestamp 1666199351
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_461
timestamp 1666199351
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_473
timestamp 1666199351
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_485
timestamp 1666199351
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1666199351
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1666199351
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_505
timestamp 1666199351
transform 1 0 47564 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_513
timestamp 1666199351
transform 1 0 48300 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1666199351
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1666199351
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1666199351
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1666199351
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1666199351
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1666199351
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1666199351
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1666199351
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1666199351
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1666199351
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1666199351
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1666199351
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1666199351
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1666199351
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1666199351
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1666199351
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1666199351
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1666199351
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1666199351
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1666199351
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1666199351
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1666199351
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1666199351
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1666199351
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1666199351
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1666199351
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1666199351
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1666199351
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1666199351
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1666199351
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_289
timestamp 1666199351
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1666199351
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1666199351
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1666199351
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1666199351
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_333
timestamp 1666199351
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1666199351
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1666199351
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1666199351
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1666199351
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1666199351
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1666199351
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_401
timestamp 1666199351
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1666199351
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1666199351
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_421
timestamp 1666199351
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_433
timestamp 1666199351
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_445
timestamp 1666199351
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_457
timestamp 1666199351
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1666199351
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1666199351
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_477
timestamp 1666199351
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_489
timestamp 1666199351
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_501
timestamp 1666199351
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_513
timestamp 1666199351
transform 1 0 48300 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1666199351
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1666199351
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1666199351
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1666199351
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1666199351
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1666199351
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1666199351
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1666199351
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1666199351
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1666199351
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1666199351
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1666199351
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1666199351
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1666199351
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1666199351
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1666199351
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1666199351
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1666199351
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1666199351
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1666199351
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1666199351
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1666199351
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1666199351
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1666199351
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1666199351
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1666199351
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1666199351
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1666199351
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1666199351
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1666199351
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1666199351
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1666199351
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1666199351
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1666199351
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1666199351
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1666199351
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1666199351
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1666199351
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1666199351
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1666199351
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1666199351
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1666199351
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1666199351
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_405
timestamp 1666199351
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_417
timestamp 1666199351
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_429
timestamp 1666199351
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1666199351
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1666199351
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_449
timestamp 1666199351
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_461
timestamp 1666199351
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_473
timestamp 1666199351
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_485
timestamp 1666199351
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1666199351
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1666199351
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_505
timestamp 1666199351
transform 1 0 47564 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_513
timestamp 1666199351
transform 1 0 48300 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1666199351
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1666199351
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1666199351
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1666199351
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1666199351
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1666199351
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1666199351
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1666199351
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1666199351
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1666199351
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1666199351
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1666199351
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1666199351
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1666199351
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1666199351
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1666199351
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1666199351
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1666199351
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1666199351
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1666199351
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1666199351
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1666199351
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1666199351
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1666199351
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1666199351
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1666199351
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1666199351
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1666199351
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1666199351
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1666199351
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_289
timestamp 1666199351
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1666199351
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1666199351
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1666199351
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1666199351
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1666199351
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1666199351
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1666199351
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1666199351
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1666199351
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1666199351
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1666199351
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_401
timestamp 1666199351
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 1666199351
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1666199351
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_421
timestamp 1666199351
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_433
timestamp 1666199351
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_445
timestamp 1666199351
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_457
timestamp 1666199351
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1666199351
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1666199351
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_477
timestamp 1666199351
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_489
timestamp 1666199351
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_501
timestamp 1666199351
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_513
timestamp 1666199351
transform 1 0 48300 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1666199351
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1666199351
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1666199351
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1666199351
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1666199351
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1666199351
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1666199351
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1666199351
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1666199351
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1666199351
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1666199351
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1666199351
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1666199351
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1666199351
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1666199351
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1666199351
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1666199351
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1666199351
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1666199351
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1666199351
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1666199351
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1666199351
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1666199351
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1666199351
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1666199351
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1666199351
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1666199351
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1666199351
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1666199351
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1666199351
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1666199351
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1666199351
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1666199351
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1666199351
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1666199351
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1666199351
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1666199351
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1666199351
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1666199351
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1666199351
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1666199351
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1666199351
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1666199351
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_405
timestamp 1666199351
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_417
timestamp 1666199351
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_429
timestamp 1666199351
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1666199351
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1666199351
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_449
timestamp 1666199351
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_461
timestamp 1666199351
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_473
timestamp 1666199351
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_485
timestamp 1666199351
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1666199351
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1666199351
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_505
timestamp 1666199351
transform 1 0 47564 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_513
timestamp 1666199351
transform 1 0 48300 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1666199351
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1666199351
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1666199351
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1666199351
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1666199351
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1666199351
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1666199351
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1666199351
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1666199351
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1666199351
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1666199351
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1666199351
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1666199351
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1666199351
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1666199351
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1666199351
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1666199351
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1666199351
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1666199351
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1666199351
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1666199351
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1666199351
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1666199351
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1666199351
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1666199351
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1666199351
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1666199351
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1666199351
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1666199351
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1666199351
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_289
timestamp 1666199351
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1666199351
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1666199351
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1666199351
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1666199351
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1666199351
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1666199351
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1666199351
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1666199351
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1666199351
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1666199351
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1666199351
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_401
timestamp 1666199351
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1666199351
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1666199351
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_421
timestamp 1666199351
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_433
timestamp 1666199351
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_445
timestamp 1666199351
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_457
timestamp 1666199351
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1666199351
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1666199351
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_477
timestamp 1666199351
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_489
timestamp 1666199351
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_501
timestamp 1666199351
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_513
timestamp 1666199351
transform 1 0 48300 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1666199351
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1666199351
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1666199351
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1666199351
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1666199351
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1666199351
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1666199351
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1666199351
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1666199351
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1666199351
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1666199351
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1666199351
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1666199351
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1666199351
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1666199351
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1666199351
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1666199351
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1666199351
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1666199351
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1666199351
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_193
timestamp 1666199351
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_205
timestamp 1666199351
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1666199351
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1666199351
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1666199351
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1666199351
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1666199351
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1666199351
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1666199351
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1666199351
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1666199351
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1666199351
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1666199351
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1666199351
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1666199351
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1666199351
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1666199351
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1666199351
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1666199351
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1666199351
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1666199351
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1666199351
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1666199351
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_405
timestamp 1666199351
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_417
timestamp 1666199351
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_429
timestamp 1666199351
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1666199351
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1666199351
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_449
timestamp 1666199351
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_461
timestamp 1666199351
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_473
timestamp 1666199351
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_485
timestamp 1666199351
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1666199351
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1666199351
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_505
timestamp 1666199351
transform 1 0 47564 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_513
timestamp 1666199351
transform 1 0 48300 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1666199351
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1666199351
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1666199351
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1666199351
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1666199351
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1666199351
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1666199351
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1666199351
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1666199351
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1666199351
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1666199351
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1666199351
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1666199351
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1666199351
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1666199351
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1666199351
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1666199351
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_165
timestamp 1666199351
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_177
timestamp 1666199351
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1666199351
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1666199351
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1666199351
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1666199351
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1666199351
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_233
timestamp 1666199351
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1666199351
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1666199351
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1666199351
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1666199351
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1666199351
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1666199351
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1666199351
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1666199351
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1666199351
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1666199351
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1666199351
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1666199351
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1666199351
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1666199351
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1666199351
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1666199351
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1666199351
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_401
timestamp 1666199351
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1666199351
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1666199351
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_421
timestamp 1666199351
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_433
timestamp 1666199351
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_445
timestamp 1666199351
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_457
timestamp 1666199351
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1666199351
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1666199351
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_477
timestamp 1666199351
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_489
timestamp 1666199351
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_501
timestamp 1666199351
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_513
timestamp 1666199351
transform 1 0 48300 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1666199351
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1666199351
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1666199351
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1666199351
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1666199351
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1666199351
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1666199351
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1666199351
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1666199351
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1666199351
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1666199351
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1666199351
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1666199351
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1666199351
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1666199351
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1666199351
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1666199351
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1666199351
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1666199351
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1666199351
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1666199351
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_205
timestamp 1666199351
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1666199351
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1666199351
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1666199351
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1666199351
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1666199351
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 1666199351
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1666199351
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1666199351
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1666199351
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1666199351
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1666199351
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1666199351
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1666199351
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1666199351
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1666199351
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1666199351
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1666199351
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1666199351
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1666199351
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1666199351
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1666199351
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_405
timestamp 1666199351
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_417
timestamp 1666199351
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_429
timestamp 1666199351
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1666199351
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1666199351
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_449
timestamp 1666199351
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_461
timestamp 1666199351
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_473
timestamp 1666199351
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_485
timestamp 1666199351
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1666199351
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1666199351
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_505
timestamp 1666199351
transform 1 0 47564 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_513
timestamp 1666199351
transform 1 0 48300 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1666199351
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1666199351
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1666199351
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1666199351
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1666199351
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1666199351
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1666199351
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1666199351
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1666199351
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1666199351
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1666199351
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1666199351
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1666199351
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1666199351
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1666199351
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1666199351
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1666199351
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1666199351
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1666199351
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1666199351
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1666199351
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1666199351
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1666199351
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1666199351
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_233
timestamp 1666199351
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1666199351
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1666199351
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1666199351
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1666199351
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1666199351
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_289
timestamp 1666199351
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1666199351
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1666199351
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1666199351
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1666199351
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1666199351
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1666199351
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1666199351
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1666199351
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1666199351
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1666199351
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1666199351
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_401
timestamp 1666199351
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1666199351
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1666199351
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_421
timestamp 1666199351
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_433
timestamp 1666199351
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_445
timestamp 1666199351
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_457
timestamp 1666199351
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1666199351
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1666199351
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_477
timestamp 1666199351
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_489
timestamp 1666199351
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_501
timestamp 1666199351
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_513
timestamp 1666199351
transform 1 0 48300 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1666199351
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1666199351
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1666199351
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1666199351
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1666199351
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1666199351
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1666199351
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1666199351
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1666199351
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1666199351
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1666199351
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1666199351
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1666199351
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1666199351
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1666199351
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1666199351
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1666199351
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1666199351
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1666199351
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1666199351
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1666199351
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1666199351
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1666199351
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1666199351
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1666199351
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1666199351
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1666199351
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1666199351
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1666199351
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1666199351
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1666199351
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1666199351
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1666199351
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_317
timestamp 1666199351
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1666199351
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1666199351
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1666199351
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1666199351
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1666199351
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1666199351
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1666199351
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1666199351
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_393
timestamp 1666199351
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_405
timestamp 1666199351
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_417
timestamp 1666199351
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_429
timestamp 1666199351
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1666199351
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1666199351
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_449
timestamp 1666199351
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_461
timestamp 1666199351
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_473
timestamp 1666199351
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_485
timestamp 1666199351
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1666199351
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1666199351
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_505
timestamp 1666199351
transform 1 0 47564 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_513
timestamp 1666199351
transform 1 0 48300 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1666199351
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1666199351
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1666199351
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1666199351
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1666199351
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1666199351
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1666199351
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1666199351
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1666199351
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1666199351
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1666199351
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1666199351
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1666199351
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1666199351
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1666199351
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1666199351
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1666199351
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1666199351
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1666199351
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1666199351
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1666199351
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1666199351
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1666199351
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1666199351
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_233
timestamp 1666199351
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1666199351
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1666199351
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1666199351
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1666199351
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1666199351
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1666199351
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1666199351
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1666199351
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1666199351
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1666199351
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1666199351
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1666199351
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1666199351
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1666199351
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1666199351
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1666199351
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1666199351
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_401
timestamp 1666199351
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 1666199351
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1666199351
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_421
timestamp 1666199351
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_433
timestamp 1666199351
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_445
timestamp 1666199351
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_457
timestamp 1666199351
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1666199351
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1666199351
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_477
timestamp 1666199351
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_489
timestamp 1666199351
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_501
timestamp 1666199351
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_513
timestamp 1666199351
transform 1 0 48300 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1666199351
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1666199351
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1666199351
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1666199351
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1666199351
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1666199351
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1666199351
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1666199351
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1666199351
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1666199351
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1666199351
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1666199351
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1666199351
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1666199351
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1666199351
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1666199351
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1666199351
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1666199351
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1666199351
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1666199351
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1666199351
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1666199351
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1666199351
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1666199351
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1666199351
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1666199351
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1666199351
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_261
timestamp 1666199351
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1666199351
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1666199351
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1666199351
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1666199351
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1666199351
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1666199351
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1666199351
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1666199351
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1666199351
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1666199351
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1666199351
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1666199351
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1666199351
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1666199351
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1666199351
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_405
timestamp 1666199351
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_417
timestamp 1666199351
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_429
timestamp 1666199351
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1666199351
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1666199351
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_449
timestamp 1666199351
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_461
timestamp 1666199351
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_473
timestamp 1666199351
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_485
timestamp 1666199351
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1666199351
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1666199351
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_505
timestamp 1666199351
transform 1 0 47564 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_513
timestamp 1666199351
transform 1 0 48300 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1666199351
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1666199351
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1666199351
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1666199351
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1666199351
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1666199351
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1666199351
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1666199351
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1666199351
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1666199351
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1666199351
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1666199351
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1666199351
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1666199351
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1666199351
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1666199351
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1666199351
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1666199351
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1666199351
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1666199351
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1666199351
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1666199351
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1666199351
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1666199351
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1666199351
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1666199351
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1666199351
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1666199351
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1666199351
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1666199351
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1666199351
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1666199351
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1666199351
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1666199351
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1666199351
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1666199351
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1666199351
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1666199351
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1666199351
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1666199351
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1666199351
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1666199351
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_401
timestamp 1666199351
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1666199351
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1666199351
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_421
timestamp 1666199351
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_433
timestamp 1666199351
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_445
timestamp 1666199351
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_457
timestamp 1666199351
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1666199351
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1666199351
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_477
timestamp 1666199351
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_489
timestamp 1666199351
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_501
timestamp 1666199351
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_513
timestamp 1666199351
transform 1 0 48300 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1666199351
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1666199351
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1666199351
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1666199351
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1666199351
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1666199351
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1666199351
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1666199351
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1666199351
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1666199351
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1666199351
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1666199351
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1666199351
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1666199351
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1666199351
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1666199351
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1666199351
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1666199351
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1666199351
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1666199351
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1666199351
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1666199351
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1666199351
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1666199351
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1666199351
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1666199351
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1666199351
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1666199351
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1666199351
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1666199351
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1666199351
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1666199351
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1666199351
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1666199351
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1666199351
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1666199351
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1666199351
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1666199351
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1666199351
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1666199351
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1666199351
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1666199351
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_393
timestamp 1666199351
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_405
timestamp 1666199351
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_417
timestamp 1666199351
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_429
timestamp 1666199351
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1666199351
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1666199351
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_449
timestamp 1666199351
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_461
timestamp 1666199351
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_473
timestamp 1666199351
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_485
timestamp 1666199351
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1666199351
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1666199351
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_505
timestamp 1666199351
transform 1 0 47564 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_513
timestamp 1666199351
transform 1 0 48300 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1666199351
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1666199351
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1666199351
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1666199351
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1666199351
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1666199351
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1666199351
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1666199351
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1666199351
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1666199351
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1666199351
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1666199351
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1666199351
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1666199351
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1666199351
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1666199351
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1666199351
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1666199351
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1666199351
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1666199351
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1666199351
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1666199351
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1666199351
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1666199351
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1666199351
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1666199351
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1666199351
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1666199351
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1666199351
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1666199351
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1666199351
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1666199351
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1666199351
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1666199351
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1666199351
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1666199351
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1666199351
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1666199351
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1666199351
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1666199351
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1666199351
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1666199351
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_401
timestamp 1666199351
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1666199351
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1666199351
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_421
timestamp 1666199351
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_433
timestamp 1666199351
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_445
timestamp 1666199351
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_457
timestamp 1666199351
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1666199351
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1666199351
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_477
timestamp 1666199351
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_489
timestamp 1666199351
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_501
timestamp 1666199351
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_513
timestamp 1666199351
transform 1 0 48300 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1666199351
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1666199351
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1666199351
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1666199351
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1666199351
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1666199351
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1666199351
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1666199351
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1666199351
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1666199351
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1666199351
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1666199351
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1666199351
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1666199351
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1666199351
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1666199351
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1666199351
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1666199351
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1666199351
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1666199351
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1666199351
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1666199351
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1666199351
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1666199351
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1666199351
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1666199351
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1666199351
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1666199351
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1666199351
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1666199351
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1666199351
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1666199351
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1666199351
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1666199351
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1666199351
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1666199351
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1666199351
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1666199351
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1666199351
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1666199351
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1666199351
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1666199351
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1666199351
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_405
timestamp 1666199351
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_417
timestamp 1666199351
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_429
timestamp 1666199351
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1666199351
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1666199351
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_449
timestamp 1666199351
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_461
timestamp 1666199351
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_473
timestamp 1666199351
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_485
timestamp 1666199351
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1666199351
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1666199351
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_505
timestamp 1666199351
transform 1 0 47564 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_513
timestamp 1666199351
transform 1 0 48300 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1666199351
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1666199351
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1666199351
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1666199351
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1666199351
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1666199351
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1666199351
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1666199351
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1666199351
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1666199351
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1666199351
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1666199351
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1666199351
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1666199351
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1666199351
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1666199351
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1666199351
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1666199351
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1666199351
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1666199351
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1666199351
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1666199351
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1666199351
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1666199351
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1666199351
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1666199351
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1666199351
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1666199351
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1666199351
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1666199351
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1666199351
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1666199351
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1666199351
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1666199351
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1666199351
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1666199351
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1666199351
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1666199351
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1666199351
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1666199351
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1666199351
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1666199351
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_401
timestamp 1666199351
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1666199351
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1666199351
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_421
timestamp 1666199351
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_433
timestamp 1666199351
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_445
timestamp 1666199351
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_457
timestamp 1666199351
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1666199351
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1666199351
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_477
timestamp 1666199351
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_489
timestamp 1666199351
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_501
timestamp 1666199351
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_513
timestamp 1666199351
transform 1 0 48300 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1666199351
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1666199351
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1666199351
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1666199351
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1666199351
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1666199351
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1666199351
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1666199351
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1666199351
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1666199351
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1666199351
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1666199351
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1666199351
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1666199351
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1666199351
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1666199351
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1666199351
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1666199351
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1666199351
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1666199351
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1666199351
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1666199351
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1666199351
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1666199351
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1666199351
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1666199351
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1666199351
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1666199351
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1666199351
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1666199351
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1666199351
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1666199351
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1666199351
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1666199351
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1666199351
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1666199351
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1666199351
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1666199351
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1666199351
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1666199351
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1666199351
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1666199351
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1666199351
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_405
timestamp 1666199351
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_417
timestamp 1666199351
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_429
timestamp 1666199351
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1666199351
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1666199351
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_449
timestamp 1666199351
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_461
timestamp 1666199351
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_473
timestamp 1666199351
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_485
timestamp 1666199351
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1666199351
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1666199351
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_505
timestamp 1666199351
transform 1 0 47564 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_513
timestamp 1666199351
transform 1 0 48300 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1666199351
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1666199351
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1666199351
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1666199351
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1666199351
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1666199351
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1666199351
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1666199351
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1666199351
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1666199351
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1666199351
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1666199351
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1666199351
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1666199351
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1666199351
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1666199351
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1666199351
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1666199351
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1666199351
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1666199351
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1666199351
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1666199351
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1666199351
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1666199351
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1666199351
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1666199351
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1666199351
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1666199351
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1666199351
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1666199351
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1666199351
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1666199351
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1666199351
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1666199351
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1666199351
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1666199351
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1666199351
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1666199351
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1666199351
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1666199351
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1666199351
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1666199351
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_401
timestamp 1666199351
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1666199351
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1666199351
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_421
timestamp 1666199351
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_433
timestamp 1666199351
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_445
timestamp 1666199351
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_457
timestamp 1666199351
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1666199351
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1666199351
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_477
timestamp 1666199351
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_489
timestamp 1666199351
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_501
timestamp 1666199351
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_513
timestamp 1666199351
transform 1 0 48300 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1666199351
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1666199351
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1666199351
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1666199351
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1666199351
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1666199351
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1666199351
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1666199351
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1666199351
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1666199351
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1666199351
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1666199351
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1666199351
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1666199351
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1666199351
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1666199351
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1666199351
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1666199351
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1666199351
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1666199351
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1666199351
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1666199351
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1666199351
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1666199351
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1666199351
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1666199351
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1666199351
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1666199351
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1666199351
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1666199351
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1666199351
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1666199351
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1666199351
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1666199351
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1666199351
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1666199351
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1666199351
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1666199351
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1666199351
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1666199351
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1666199351
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1666199351
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1666199351
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_405
timestamp 1666199351
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_417
timestamp 1666199351
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_429
timestamp 1666199351
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1666199351
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1666199351
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_449
timestamp 1666199351
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_461
timestamp 1666199351
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_473
timestamp 1666199351
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_485
timestamp 1666199351
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1666199351
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1666199351
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_505
timestamp 1666199351
transform 1 0 47564 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_513
timestamp 1666199351
transform 1 0 48300 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1666199351
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1666199351
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1666199351
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1666199351
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1666199351
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1666199351
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1666199351
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1666199351
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1666199351
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1666199351
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1666199351
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1666199351
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1666199351
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1666199351
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1666199351
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1666199351
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1666199351
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1666199351
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1666199351
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1666199351
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1666199351
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1666199351
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1666199351
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1666199351
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1666199351
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1666199351
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1666199351
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1666199351
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1666199351
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1666199351
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1666199351
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1666199351
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1666199351
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1666199351
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1666199351
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1666199351
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1666199351
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1666199351
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1666199351
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1666199351
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1666199351
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_389
timestamp 1666199351
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_401
timestamp 1666199351
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1666199351
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1666199351
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_421
timestamp 1666199351
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_433
timestamp 1666199351
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_445
timestamp 1666199351
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_457
timestamp 1666199351
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1666199351
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1666199351
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_477
timestamp 1666199351
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_489
timestamp 1666199351
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_501
timestamp 1666199351
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_513
timestamp 1666199351
transform 1 0 48300 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1666199351
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1666199351
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1666199351
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1666199351
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1666199351
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1666199351
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1666199351
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1666199351
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1666199351
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1666199351
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1666199351
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1666199351
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1666199351
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1666199351
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1666199351
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1666199351
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1666199351
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1666199351
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1666199351
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1666199351
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1666199351
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_205
timestamp 1666199351
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1666199351
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1666199351
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1666199351
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_237
timestamp 1666199351
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_249
timestamp 1666199351
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_261
timestamp 1666199351
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1666199351
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1666199351
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1666199351
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1666199351
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_305
timestamp 1666199351
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_317
timestamp 1666199351
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1666199351
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1666199351
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1666199351
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1666199351
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1666199351
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_373
timestamp 1666199351
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1666199351
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1666199351
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_393
timestamp 1666199351
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_405
timestamp 1666199351
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_417
timestamp 1666199351
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_429
timestamp 1666199351
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1666199351
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1666199351
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_449
timestamp 1666199351
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_461
timestamp 1666199351
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_473
timestamp 1666199351
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_485
timestamp 1666199351
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1666199351
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1666199351
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_505
timestamp 1666199351
transform 1 0 47564 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_513
timestamp 1666199351
transform 1 0 48300 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1666199351
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1666199351
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1666199351
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1666199351
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1666199351
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1666199351
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_65
timestamp 1666199351
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1666199351
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1666199351
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1666199351
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1666199351
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1666199351
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_121
timestamp 1666199351
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1666199351
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1666199351
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1666199351
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1666199351
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_165
timestamp 1666199351
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_177
timestamp 1666199351
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1666199351
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1666199351
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_197
timestamp 1666199351
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_209
timestamp 1666199351
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_221
timestamp 1666199351
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_233
timestamp 1666199351
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1666199351
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1666199351
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_253
timestamp 1666199351
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_265
timestamp 1666199351
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_277
timestamp 1666199351
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_289
timestamp 1666199351
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1666199351
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1666199351
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_309
timestamp 1666199351
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_321
timestamp 1666199351
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_333
timestamp 1666199351
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_345
timestamp 1666199351
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1666199351
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1666199351
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_365
timestamp 1666199351
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_377
timestamp 1666199351
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_389
timestamp 1666199351
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_401
timestamp 1666199351
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1666199351
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1666199351
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_421
timestamp 1666199351
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_433
timestamp 1666199351
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_445
timestamp 1666199351
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_457
timestamp 1666199351
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1666199351
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1666199351
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_477
timestamp 1666199351
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_489
timestamp 1666199351
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_501
timestamp 1666199351
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_513
timestamp 1666199351
transform 1 0 48300 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1666199351
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1666199351
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1666199351
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_39
timestamp 1666199351
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1666199351
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1666199351
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1666199351
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_69
timestamp 1666199351
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_81
timestamp 1666199351
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_93
timestamp 1666199351
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1666199351
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1666199351
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1666199351
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_125
timestamp 1666199351
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_137
timestamp 1666199351
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_149
timestamp 1666199351
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1666199351
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1666199351
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_169
timestamp 1666199351
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_181
timestamp 1666199351
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_193
timestamp 1666199351
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_205
timestamp 1666199351
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1666199351
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1666199351
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_225
timestamp 1666199351
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_237
timestamp 1666199351
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_249
timestamp 1666199351
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_261
timestamp 1666199351
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_273
timestamp 1666199351
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1666199351
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_281
timestamp 1666199351
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_293
timestamp 1666199351
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_305
timestamp 1666199351
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_317
timestamp 1666199351
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 1666199351
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1666199351
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_337
timestamp 1666199351
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_349
timestamp 1666199351
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_361
timestamp 1666199351
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_373
timestamp 1666199351
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1666199351
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1666199351
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_393
timestamp 1666199351
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_405
timestamp 1666199351
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_417
timestamp 1666199351
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_429
timestamp 1666199351
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1666199351
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1666199351
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_449
timestamp 1666199351
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_461
timestamp 1666199351
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_473
timestamp 1666199351
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_485
timestamp 1666199351
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1666199351
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1666199351
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_505
timestamp 1666199351
transform 1 0 47564 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_513
timestamp 1666199351
transform 1 0 48300 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1666199351
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1666199351
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1666199351
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1666199351
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1666199351
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1666199351
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1666199351
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1666199351
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1666199351
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1666199351
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1666199351
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1666199351
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1666199351
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1666199351
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1666199351
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1666199351
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_153
timestamp 1666199351
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_165
timestamp 1666199351
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_177
timestamp 1666199351
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1666199351
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1666199351
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_197
timestamp 1666199351
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_209
timestamp 1666199351
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_221
timestamp 1666199351
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_233
timestamp 1666199351
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1666199351
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1666199351
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_253
timestamp 1666199351
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_265
timestamp 1666199351
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_277
timestamp 1666199351
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_289
timestamp 1666199351
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_301
timestamp 1666199351
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1666199351
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_309
timestamp 1666199351
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_321
timestamp 1666199351
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_333
timestamp 1666199351
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_345
timestamp 1666199351
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1666199351
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1666199351
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_365
timestamp 1666199351
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_377
timestamp 1666199351
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_389
timestamp 1666199351
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_401
timestamp 1666199351
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1666199351
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1666199351
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_421
timestamp 1666199351
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_433
timestamp 1666199351
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_445
timestamp 1666199351
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_457
timestamp 1666199351
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1666199351
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1666199351
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_477
timestamp 1666199351
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_489
timestamp 1666199351
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_501
timestamp 1666199351
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_513
timestamp 1666199351
transform 1 0 48300 0 1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1666199351
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1666199351
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1666199351
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_39
timestamp 1666199351
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1666199351
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1666199351
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1666199351
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1666199351
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1666199351
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1666199351
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1666199351
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1666199351
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1666199351
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1666199351
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 1666199351
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_149
timestamp 1666199351
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1666199351
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1666199351
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_169
timestamp 1666199351
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_181
timestamp 1666199351
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_193
timestamp 1666199351
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_205
timestamp 1666199351
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1666199351
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1666199351
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_225
timestamp 1666199351
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_237
timestamp 1666199351
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_249
timestamp 1666199351
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_261
timestamp 1666199351
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_273
timestamp 1666199351
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1666199351
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_281
timestamp 1666199351
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_293
timestamp 1666199351
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_305
timestamp 1666199351
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_317
timestamp 1666199351
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1666199351
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1666199351
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_337
timestamp 1666199351
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_349
timestamp 1666199351
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_361
timestamp 1666199351
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_373
timestamp 1666199351
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1666199351
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1666199351
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_393
timestamp 1666199351
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_405
timestamp 1666199351
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_417
timestamp 1666199351
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_429
timestamp 1666199351
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1666199351
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1666199351
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_449
timestamp 1666199351
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_461
timestamp 1666199351
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_473
timestamp 1666199351
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_485
timestamp 1666199351
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1666199351
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1666199351
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_505
timestamp 1666199351
transform 1 0 47564 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_513
timestamp 1666199351
transform 1 0 48300 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1666199351
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1666199351
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1666199351
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1666199351
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1666199351
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1666199351
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1666199351
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1666199351
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1666199351
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1666199351
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1666199351
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_109
timestamp 1666199351
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_121
timestamp 1666199351
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1666199351
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1666199351
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1666199351
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1666199351
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_165
timestamp 1666199351
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_177
timestamp 1666199351
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1666199351
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1666199351
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_197
timestamp 1666199351
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_209
timestamp 1666199351
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_221
timestamp 1666199351
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_233
timestamp 1666199351
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_245
timestamp 1666199351
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1666199351
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_253
timestamp 1666199351
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_265
timestamp 1666199351
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_277
timestamp 1666199351
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_289
timestamp 1666199351
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 1666199351
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1666199351
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_309
timestamp 1666199351
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_321
timestamp 1666199351
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_333
timestamp 1666199351
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_345
timestamp 1666199351
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1666199351
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1666199351
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_365
timestamp 1666199351
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_377
timestamp 1666199351
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_389
timestamp 1666199351
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_401
timestamp 1666199351
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1666199351
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1666199351
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_421
timestamp 1666199351
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_433
timestamp 1666199351
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_445
timestamp 1666199351
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_457
timestamp 1666199351
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1666199351
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1666199351
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_477
timestamp 1666199351
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_489
timestamp 1666199351
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_501
timestamp 1666199351
transform 1 0 47196 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_513
timestamp 1666199351
transform 1 0 48300 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1666199351
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1666199351
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1666199351
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1666199351
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1666199351
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1666199351
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1666199351
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1666199351
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1666199351
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1666199351
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1666199351
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1666199351
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1666199351
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_125
timestamp 1666199351
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_137
timestamp 1666199351
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_149
timestamp 1666199351
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1666199351
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1666199351
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_169
timestamp 1666199351
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_181
timestamp 1666199351
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_193
timestamp 1666199351
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_205
timestamp 1666199351
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1666199351
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1666199351
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_225
timestamp 1666199351
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_237
timestamp 1666199351
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_249
timestamp 1666199351
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_261
timestamp 1666199351
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1666199351
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1666199351
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_281
timestamp 1666199351
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_293
timestamp 1666199351
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_305
timestamp 1666199351
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_317
timestamp 1666199351
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1666199351
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1666199351
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_337
timestamp 1666199351
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_349
timestamp 1666199351
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_361
timestamp 1666199351
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_373
timestamp 1666199351
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1666199351
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1666199351
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_393
timestamp 1666199351
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_405
timestamp 1666199351
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_417
timestamp 1666199351
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_429
timestamp 1666199351
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1666199351
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1666199351
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_449
timestamp 1666199351
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_461
timestamp 1666199351
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_473
timestamp 1666199351
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_485
timestamp 1666199351
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1666199351
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1666199351
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_505
timestamp 1666199351
transform 1 0 47564 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_513
timestamp 1666199351
transform 1 0 48300 0 -1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1666199351
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1666199351
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1666199351
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1666199351
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1666199351
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1666199351
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1666199351
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1666199351
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1666199351
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1666199351
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1666199351
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_109
timestamp 1666199351
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_121
timestamp 1666199351
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1666199351
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1666199351
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1666199351
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_153
timestamp 1666199351
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_165
timestamp 1666199351
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_177
timestamp 1666199351
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1666199351
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1666199351
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_197
timestamp 1666199351
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_209
timestamp 1666199351
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_221
timestamp 1666199351
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_233
timestamp 1666199351
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1666199351
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1666199351
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_253
timestamp 1666199351
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_265
timestamp 1666199351
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_277
timestamp 1666199351
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_289
timestamp 1666199351
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_301
timestamp 1666199351
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1666199351
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_309
timestamp 1666199351
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_321
timestamp 1666199351
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_333
timestamp 1666199351
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_345
timestamp 1666199351
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1666199351
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1666199351
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_365
timestamp 1666199351
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_377
timestamp 1666199351
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_389
timestamp 1666199351
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_401
timestamp 1666199351
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1666199351
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1666199351
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_421
timestamp 1666199351
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_433
timestamp 1666199351
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_445
timestamp 1666199351
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_457
timestamp 1666199351
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1666199351
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1666199351
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_477
timestamp 1666199351
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_489
timestamp 1666199351
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_501
timestamp 1666199351
transform 1 0 47196 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_513
timestamp 1666199351
transform 1 0 48300 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1666199351
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1666199351
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1666199351
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_39
timestamp 1666199351
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1666199351
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1666199351
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1666199351
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1666199351
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1666199351
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 1666199351
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1666199351
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1666199351
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1666199351
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1666199351
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_137
timestamp 1666199351
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_149
timestamp 1666199351
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1666199351
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1666199351
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_169
timestamp 1666199351
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_181
timestamp 1666199351
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_193
timestamp 1666199351
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_205
timestamp 1666199351
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1666199351
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1666199351
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_225
timestamp 1666199351
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_237
timestamp 1666199351
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_249
timestamp 1666199351
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_261
timestamp 1666199351
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1666199351
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1666199351
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_281
timestamp 1666199351
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_293
timestamp 1666199351
transform 1 0 28060 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_297
timestamp 1666199351
transform 1 0 28428 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_300
timestamp 1666199351
transform 1 0 28704 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_312
timestamp 1666199351
transform 1 0 29808 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_324
timestamp 1666199351
transform 1 0 30912 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_337
timestamp 1666199351
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_349
timestamp 1666199351
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_361
timestamp 1666199351
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_373
timestamp 1666199351
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1666199351
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1666199351
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_393
timestamp 1666199351
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_405
timestamp 1666199351
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_417
timestamp 1666199351
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_429
timestamp 1666199351
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1666199351
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1666199351
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_449
timestamp 1666199351
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_461
timestamp 1666199351
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_473
timestamp 1666199351
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_485
timestamp 1666199351
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_497
timestamp 1666199351
transform 1 0 46828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_503
timestamp 1666199351
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_505
timestamp 1666199351
transform 1 0 47564 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_513
timestamp 1666199351
transform 1 0 48300 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1666199351
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1666199351
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1666199351
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1666199351
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1666199351
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1666199351
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1666199351
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1666199351
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1666199351
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1666199351
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1666199351
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_109
timestamp 1666199351
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_121
timestamp 1666199351
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1666199351
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1666199351
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1666199351
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_153
timestamp 1666199351
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_165
timestamp 1666199351
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_177
timestamp 1666199351
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1666199351
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1666199351
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_197
timestamp 1666199351
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_209
timestamp 1666199351
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_221
timestamp 1666199351
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_233
timestamp 1666199351
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1666199351
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1666199351
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_253
timestamp 1666199351
transform 1 0 24380 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_261
timestamp 1666199351
transform 1 0 25116 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_72_265
timestamp 1666199351
transform 1 0 25484 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_271
timestamp 1666199351
transform 1 0 26036 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_274
timestamp 1666199351
transform 1 0 26312 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_72_282
timestamp 1666199351
transform 1 0 27048 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_290
timestamp 1666199351
transform 1 0 27784 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_294
timestamp 1666199351
transform 1 0 28152 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_298
timestamp 1666199351
transform 1 0 28520 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1666199351
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1666199351
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_309
timestamp 1666199351
transform 1 0 29532 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_313
timestamp 1666199351
transform 1 0 29900 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_319
timestamp 1666199351
transform 1 0 30452 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_325
timestamp 1666199351
transform 1 0 31004 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_337
timestamp 1666199351
transform 1 0 32108 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_349
timestamp 1666199351
transform 1 0 33212 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_72_361
timestamp 1666199351
transform 1 0 34316 0 1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_72_365
timestamp 1666199351
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_377
timestamp 1666199351
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_389
timestamp 1666199351
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_401
timestamp 1666199351
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1666199351
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1666199351
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_421
timestamp 1666199351
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_433
timestamp 1666199351
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_445
timestamp 1666199351
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_457
timestamp 1666199351
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1666199351
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1666199351
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_477
timestamp 1666199351
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_489
timestamp 1666199351
transform 1 0 46092 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_501
timestamp 1666199351
transform 1 0 47196 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_72_513
timestamp 1666199351
transform 1 0 48300 0 1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1666199351
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1666199351
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1666199351
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1666199351
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1666199351
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1666199351
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1666199351
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1666199351
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_81
timestamp 1666199351
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_93
timestamp 1666199351
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1666199351
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1666199351
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_113
timestamp 1666199351
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_125
timestamp 1666199351
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_137
timestamp 1666199351
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_149
timestamp 1666199351
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1666199351
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1666199351
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1666199351
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_181
timestamp 1666199351
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_193
timestamp 1666199351
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_205
timestamp 1666199351
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1666199351
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1666199351
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_225
timestamp 1666199351
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_237
timestamp 1666199351
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_251
timestamp 1666199351
transform 1 0 24196 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_259
timestamp 1666199351
transform 1 0 24932 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_262
timestamp 1666199351
transform 1 0 25208 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_268
timestamp 1666199351
transform 1 0 25760 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_73_274
timestamp 1666199351
transform 1 0 26312 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_73_281
timestamp 1666199351
transform 1 0 26956 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_285
timestamp 1666199351
transform 1 0 27324 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_73_291
timestamp 1666199351
transform 1 0 27876 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_297
timestamp 1666199351
transform 1 0 28428 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_300
timestamp 1666199351
transform 1 0 28704 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_306
timestamp 1666199351
transform 1 0 29256 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_73_312
timestamp 1666199351
transform 1 0 29808 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_73_320
timestamp 1666199351
transform 1 0 30544 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_326
timestamp 1666199351
transform 1 0 31096 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_332
timestamp 1666199351
transform 1 0 31648 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_337
timestamp 1666199351
transform 1 0 32108 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_341
timestamp 1666199351
transform 1 0 32476 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_345
timestamp 1666199351
transform 1 0 32844 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_348
timestamp 1666199351
transform 1 0 33120 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_354
timestamp 1666199351
transform 1 0 33672 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_73_364
timestamp 1666199351
transform 1 0 34592 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_73_370
timestamp 1666199351
transform 1 0 35144 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_73_378
timestamp 1666199351
transform 1 0 35880 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_384
timestamp 1666199351
transform 1 0 36432 0 -1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_73_393
timestamp 1666199351
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_405
timestamp 1666199351
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_417
timestamp 1666199351
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_429
timestamp 1666199351
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1666199351
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1666199351
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_449
timestamp 1666199351
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_461
timestamp 1666199351
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_473
timestamp 1666199351
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_485
timestamp 1666199351
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_497
timestamp 1666199351
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1666199351
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_505
timestamp 1666199351
transform 1 0 47564 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_73_513
timestamp 1666199351
transform 1 0 48300 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1666199351
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1666199351
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1666199351
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1666199351
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1666199351
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1666199351
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1666199351
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1666199351
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1666199351
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_85
timestamp 1666199351
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_97
timestamp 1666199351
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_109
timestamp 1666199351
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_121
timestamp 1666199351
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1666199351
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1666199351
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1666199351
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1666199351
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_165
timestamp 1666199351
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_177
timestamp 1666199351
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1666199351
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1666199351
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_197
timestamp 1666199351
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_209
timestamp 1666199351
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_221
timestamp 1666199351
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_233
timestamp 1666199351
transform 1 0 22540 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_74_239
timestamp 1666199351
transform 1 0 23092 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_247
timestamp 1666199351
transform 1 0 23828 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_250
timestamp 1666199351
transform 1 0 24104 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_253
timestamp 1666199351
transform 1 0 24380 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_260
timestamp 1666199351
transform 1 0 25024 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_266
timestamp 1666199351
transform 1 0 25576 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_272
timestamp 1666199351
transform 1 0 26128 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_278
timestamp 1666199351
transform 1 0 26680 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_74_284
timestamp 1666199351
transform 1 0 27232 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_74_292
timestamp 1666199351
transform 1 0 27968 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_296
timestamp 1666199351
transform 1 0 28336 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_299
timestamp 1666199351
transform 1 0 28612 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_74_305
timestamp 1666199351
transform 1 0 29164 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_74_309
timestamp 1666199351
transform 1 0 29532 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_313
timestamp 1666199351
transform 1 0 29900 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_319
timestamp 1666199351
transform 1 0 30452 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_325
timestamp 1666199351
transform 1 0 31004 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_331
timestamp 1666199351
transform 1 0 31556 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_337
timestamp 1666199351
transform 1 0 32108 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_343
timestamp 1666199351
transform 1 0 32660 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_74_349
timestamp 1666199351
transform 1 0 33212 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1666199351
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1666199351
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_365
timestamp 1666199351
transform 1 0 34684 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_369
timestamp 1666199351
transform 1 0 35052 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_375
timestamp 1666199351
transform 1 0 35604 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_381
timestamp 1666199351
transform 1 0 36156 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_387
timestamp 1666199351
transform 1 0 36708 0 1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_74_393
timestamp 1666199351
transform 1 0 37260 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_405
timestamp 1666199351
transform 1 0 38364 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_74_417
timestamp 1666199351
transform 1 0 39468 0 1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_74_421
timestamp 1666199351
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_433
timestamp 1666199351
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_445
timestamp 1666199351
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_457
timestamp 1666199351
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1666199351
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1666199351
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_477
timestamp 1666199351
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_489
timestamp 1666199351
transform 1 0 46092 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_501
timestamp 1666199351
transform 1 0 47196 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_74_513
timestamp 1666199351
transform 1 0 48300 0 1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1666199351
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1666199351
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_27
timestamp 1666199351
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_39
timestamp 1666199351
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1666199351
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1666199351
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1666199351
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1666199351
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1666199351
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1666199351
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1666199351
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1666199351
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1666199351
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1666199351
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_137
timestamp 1666199351
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_149
timestamp 1666199351
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1666199351
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1666199351
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1666199351
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_181
timestamp 1666199351
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_193
timestamp 1666199351
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_205
timestamp 1666199351
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1666199351
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1666199351
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_225
timestamp 1666199351
transform 1 0 21804 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_233
timestamp 1666199351
transform 1 0 22540 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_75_238
timestamp 1666199351
transform 1 0 23000 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_244
timestamp 1666199351
transform 1 0 23552 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_250
timestamp 1666199351
transform 1 0 24104 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_260
timestamp 1666199351
transform 1 0 25024 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_267
timestamp 1666199351
transform 1 0 25668 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1666199351
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1666199351
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_75_281
timestamp 1666199351
transform 1 0 26956 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_290
timestamp 1666199351
transform 1 0 27784 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_297
timestamp 1666199351
transform 1 0 28428 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_303
timestamp 1666199351
transform 1 0 28980 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_309
timestamp 1666199351
transform 1 0 29532 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_315
timestamp 1666199351
transform 1 0 30084 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_75_321
timestamp 1666199351
transform 1 0 30636 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_75_332
timestamp 1666199351
transform 1 0 31648 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_337
timestamp 1666199351
transform 1 0 32108 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_341
timestamp 1666199351
transform 1 0 32476 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_75_347
timestamp 1666199351
transform 1 0 33028 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_75_356
timestamp 1666199351
transform 1 0 33856 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_362
timestamp 1666199351
transform 1 0 34408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_368
timestamp 1666199351
transform 1 0 34960 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_374
timestamp 1666199351
transform 1 0 35512 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_380
timestamp 1666199351
transform 1 0 36064 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_75_386
timestamp 1666199351
transform 1 0 36616 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_75_393
timestamp 1666199351
transform 1 0 37260 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_397
timestamp 1666199351
transform 1 0 37628 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_403
timestamp 1666199351
transform 1 0 38180 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_409
timestamp 1666199351
transform 1 0 38732 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_415
timestamp 1666199351
transform 1 0 39284 0 -1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_75_421
timestamp 1666199351
transform 1 0 39836 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_433
timestamp 1666199351
transform 1 0 40940 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_445
timestamp 1666199351
transform 1 0 42044 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_75_449
timestamp 1666199351
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_461
timestamp 1666199351
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_473
timestamp 1666199351
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_485
timestamp 1666199351
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_497
timestamp 1666199351
transform 1 0 46828 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_503
timestamp 1666199351
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_505
timestamp 1666199351
transform 1 0 47564 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_513
timestamp 1666199351
transform 1 0 48300 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1666199351
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1666199351
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1666199351
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1666199351
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1666199351
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1666199351
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1666199351
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1666199351
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1666199351
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1666199351
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1666199351
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_109
timestamp 1666199351
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_121
timestamp 1666199351
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1666199351
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1666199351
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1666199351
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1666199351
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1666199351
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_177
timestamp 1666199351
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1666199351
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1666199351
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_197
timestamp 1666199351
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_76_209
timestamp 1666199351
transform 1 0 20332 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_76_214
timestamp 1666199351
transform 1 0 20792 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_220
timestamp 1666199351
transform 1 0 21344 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_224
timestamp 1666199351
transform 1 0 21712 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_227
timestamp 1666199351
transform 1 0 21988 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_233
timestamp 1666199351
transform 1 0 22540 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_239
timestamp 1666199351
transform 1 0 23092 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_250
timestamp 1666199351
transform 1 0 24104 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_253
timestamp 1666199351
transform 1 0 24380 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_270
timestamp 1666199351
transform 1 0 25944 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_274
timestamp 1666199351
transform 1 0 26312 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_288
timestamp 1666199351
transform 1 0 27600 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_299
timestamp 1666199351
transform 1 0 28612 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_306
timestamp 1666199351
transform 1 0 29256 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_309
timestamp 1666199351
transform 1 0 29532 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_318
timestamp 1666199351
transform 1 0 30360 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_325
timestamp 1666199351
transform 1 0 31004 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_76_332
timestamp 1666199351
transform 1 0 31648 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_76_343
timestamp 1666199351
transform 1 0 32660 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_76_356
timestamp 1666199351
transform 1 0 33856 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_362
timestamp 1666199351
transform 1 0 34408 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_365
timestamp 1666199351
transform 1 0 34684 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_374
timestamp 1666199351
transform 1 0 35512 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_384
timestamp 1666199351
transform 1 0 36432 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_390
timestamp 1666199351
transform 1 0 36984 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_396
timestamp 1666199351
transform 1 0 37536 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_402
timestamp 1666199351
transform 1 0 38088 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_408
timestamp 1666199351
transform 1 0 38640 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_76_414
timestamp 1666199351
transform 1 0 39192 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_76_421
timestamp 1666199351
transform 1 0 39836 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_425
timestamp 1666199351
transform 1 0 40204 0 1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_76_431
timestamp 1666199351
transform 1 0 40756 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_443
timestamp 1666199351
transform 1 0 41860 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_455
timestamp 1666199351
transform 1 0 42964 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_467
timestamp 1666199351
transform 1 0 44068 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1666199351
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_477
timestamp 1666199351
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_489
timestamp 1666199351
transform 1 0 46092 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_501
timestamp 1666199351
transform 1 0 47196 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_76_513
timestamp 1666199351
transform 1 0 48300 0 1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1666199351
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1666199351
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1666199351
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1666199351
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1666199351
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1666199351
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1666199351
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1666199351
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_81
timestamp 1666199351
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_93
timestamp 1666199351
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1666199351
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1666199351
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1666199351
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 1666199351
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_137
timestamp 1666199351
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_149
timestamp 1666199351
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1666199351
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1666199351
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1666199351
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_181
timestamp 1666199351
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_193
timestamp 1666199351
transform 1 0 18860 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_77_203
timestamp 1666199351
transform 1 0 19780 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_207
timestamp 1666199351
transform 1 0 20148 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_210
timestamp 1666199351
transform 1 0 20424 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1666199351
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1666199351
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_77_225
timestamp 1666199351
transform 1 0 21804 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_229
timestamp 1666199351
transform 1 0 22172 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_236
timestamp 1666199351
transform 1 0 22816 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_253
timestamp 1666199351
transform 1 0 24380 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_259
timestamp 1666199351
transform 1 0 24932 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_267
timestamp 1666199351
transform 1 0 25668 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_278
timestamp 1666199351
transform 1 0 26680 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_281
timestamp 1666199351
transform 1 0 26956 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_285
timestamp 1666199351
transform 1 0 27324 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_295
timestamp 1666199351
transform 1 0 28244 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_312
timestamp 1666199351
transform 1 0 29808 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_325
timestamp 1666199351
transform 1 0 31004 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_332
timestamp 1666199351
transform 1 0 31648 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_337
timestamp 1666199351
transform 1 0 32108 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_77_345
timestamp 1666199351
transform 1 0 32844 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_351
timestamp 1666199351
transform 1 0 33396 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_359
timestamp 1666199351
transform 1 0 34132 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_376
timestamp 1666199351
transform 1 0 35696 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_387
timestamp 1666199351
transform 1 0 36708 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1666199351
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_77_393
timestamp 1666199351
transform 1 0 37260 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_402
timestamp 1666199351
transform 1 0 38088 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_408
timestamp 1666199351
transform 1 0 38640 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_414
timestamp 1666199351
transform 1 0 39192 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_420
timestamp 1666199351
transform 1 0 39744 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_426
timestamp 1666199351
transform 1 0 40296 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_77_432
timestamp 1666199351
transform 1 0 40848 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_444
timestamp 1666199351
transform 1 0 41952 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_77_449
timestamp 1666199351
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_461
timestamp 1666199351
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_473
timestamp 1666199351
transform 1 0 44620 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_485
timestamp 1666199351
transform 1 0 45724 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_497
timestamp 1666199351
transform 1 0 46828 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_503
timestamp 1666199351
transform 1 0 47380 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_505
timestamp 1666199351
transform 1 0 47564 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_77_513
timestamp 1666199351
transform 1 0 48300 0 -1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1666199351
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1666199351
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1666199351
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1666199351
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1666199351
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1666199351
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1666199351
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1666199351
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1666199351
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_85
timestamp 1666199351
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_97
timestamp 1666199351
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_109
timestamp 1666199351
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_121
timestamp 1666199351
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1666199351
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1666199351
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1666199351
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_153
timestamp 1666199351
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_165
timestamp 1666199351
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_177
timestamp 1666199351
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_78_189
timestamp 1666199351
transform 1 0 18492 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_78_194
timestamp 1666199351
transform 1 0 18952 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_78_197
timestamp 1666199351
transform 1 0 19228 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_78_206
timestamp 1666199351
transform 1 0 20056 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_210
timestamp 1666199351
transform 1 0 20424 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_217
timestamp 1666199351
transform 1 0 21068 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_78_228
timestamp 1666199351
transform 1 0 22080 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_237
timestamp 1666199351
transform 1 0 22908 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_248
timestamp 1666199351
transform 1 0 23920 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_253
timestamp 1666199351
transform 1 0 24380 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_78_263
timestamp 1666199351
transform 1 0 25300 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_78_276
timestamp 1666199351
transform 1 0 26496 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_280
timestamp 1666199351
transform 1 0 26864 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_284
timestamp 1666199351
transform 1 0 27232 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_296
timestamp 1666199351
transform 1 0 28336 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_306
timestamp 1666199351
transform 1 0 29256 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_309
timestamp 1666199351
transform 1 0 29532 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_318
timestamp 1666199351
transform 1 0 30360 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_78_325
timestamp 1666199351
transform 1 0 31004 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_331
timestamp 1666199351
transform 1 0 31556 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_338
timestamp 1666199351
transform 1 0 32200 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_355
timestamp 1666199351
transform 1 0 33764 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_362
timestamp 1666199351
transform 1 0 34408 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_365
timestamp 1666199351
transform 1 0 34684 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_370
timestamp 1666199351
transform 1 0 35144 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_374
timestamp 1666199351
transform 1 0 35512 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_384
timestamp 1666199351
transform 1 0 36432 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_401
timestamp 1666199351
transform 1 0 37996 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_408
timestamp 1666199351
transform 1 0 38640 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_78_414
timestamp 1666199351
transform 1 0 39192 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_78_421
timestamp 1666199351
transform 1 0 39836 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_425
timestamp 1666199351
transform 1 0 40204 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_431
timestamp 1666199351
transform 1 0 40756 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_437
timestamp 1666199351
transform 1 0 41308 0 1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_443
timestamp 1666199351
transform 1 0 41860 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_455
timestamp 1666199351
transform 1 0 42964 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_467
timestamp 1666199351
transform 1 0 44068 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_475
timestamp 1666199351
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_477
timestamp 1666199351
transform 1 0 44988 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_489
timestamp 1666199351
transform 1 0 46092 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_501
timestamp 1666199351
transform 1 0 47196 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_78_513
timestamp 1666199351
transform 1 0 48300 0 1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1666199351
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1666199351
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1666199351
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1666199351
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1666199351
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1666199351
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1666199351
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1666199351
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_81
timestamp 1666199351
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_93
timestamp 1666199351
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1666199351
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1666199351
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 1666199351
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_125
timestamp 1666199351
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_137
timestamp 1666199351
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_149
timestamp 1666199351
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1666199351
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1666199351
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1666199351
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_181
timestamp 1666199351
transform 1 0 17756 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_189
timestamp 1666199351
transform 1 0 18492 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_193
timestamp 1666199351
transform 1 0 18860 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_200
timestamp 1666199351
transform 1 0 19504 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_207
timestamp 1666199351
transform 1 0 20148 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_220
timestamp 1666199351
transform 1 0 21344 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_79_225
timestamp 1666199351
transform 1 0 21804 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_233
timestamp 1666199351
transform 1 0 22540 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_237
timestamp 1666199351
transform 1 0 22908 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_245
timestamp 1666199351
transform 1 0 23644 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_251
timestamp 1666199351
transform 1 0 24196 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_262
timestamp 1666199351
transform 1 0 25208 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_275
timestamp 1666199351
transform 1 0 26404 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 1666199351
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_281
timestamp 1666199351
transform 1 0 26956 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_288
timestamp 1666199351
transform 1 0 27600 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_292
timestamp 1666199351
transform 1 0 27968 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_306
timestamp 1666199351
transform 1 0 29256 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_312
timestamp 1666199351
transform 1 0 29808 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1666199351
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1666199351
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_337
timestamp 1666199351
transform 1 0 32108 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_347
timestamp 1666199351
transform 1 0 33028 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_360
timestamp 1666199351
transform 1 0 34224 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_371
timestamp 1666199351
transform 1 0 35236 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_377
timestamp 1666199351
transform 1 0 35788 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_79_386
timestamp 1666199351
transform 1 0 36616 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_79_393
timestamp 1666199351
transform 1 0 37260 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_403
timestamp 1666199351
transform 1 0 38180 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_414
timestamp 1666199351
transform 1 0 39192 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_421
timestamp 1666199351
transform 1 0 39836 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_427
timestamp 1666199351
transform 1 0 40388 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_433
timestamp 1666199351
transform 1 0 40940 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_439
timestamp 1666199351
transform 1 0 41492 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_79_445
timestamp 1666199351
transform 1 0 42044 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_79_449
timestamp 1666199351
transform 1 0 42412 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_453
timestamp 1666199351
transform 1 0 42780 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_465
timestamp 1666199351
transform 1 0 43884 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_477
timestamp 1666199351
transform 1 0 44988 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_489
timestamp 1666199351
transform 1 0 46092 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_501
timestamp 1666199351
transform 1 0 47196 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_79_505
timestamp 1666199351
transform 1 0 47564 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_513
timestamp 1666199351
transform 1 0 48300 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 1666199351
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1666199351
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1666199351
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1666199351
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1666199351
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1666199351
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_65
timestamp 1666199351
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1666199351
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1666199351
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1666199351
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_97
timestamp 1666199351
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_109
timestamp 1666199351
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_121
timestamp 1666199351
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1666199351
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1666199351
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_141
timestamp 1666199351
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_153
timestamp 1666199351
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_165
timestamp 1666199351
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_177
timestamp 1666199351
transform 1 0 17388 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_180
timestamp 1666199351
transform 1 0 17664 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_187
timestamp 1666199351
transform 1 0 18308 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_194
timestamp 1666199351
transform 1 0 18952 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_197
timestamp 1666199351
transform 1 0 19228 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_207
timestamp 1666199351
transform 1 0 20148 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_216
timestamp 1666199351
transform 1 0 20976 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_226
timestamp 1666199351
transform 1 0 21896 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_238
timestamp 1666199351
transform 1 0 23000 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_80_249
timestamp 1666199351
transform 1 0 24012 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_80_253
timestamp 1666199351
transform 1 0 24380 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_258
timestamp 1666199351
transform 1 0 24840 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_269
timestamp 1666199351
transform 1 0 25852 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_280
timestamp 1666199351
transform 1 0 26864 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_292
timestamp 1666199351
transform 1 0 27968 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_80_306
timestamp 1666199351
transform 1 0 29256 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_309
timestamp 1666199351
transform 1 0 29532 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_318
timestamp 1666199351
transform 1 0 30360 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_329
timestamp 1666199351
transform 1 0 31372 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_340
timestamp 1666199351
transform 1 0 32384 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_351
timestamp 1666199351
transform 1 0 33396 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_362
timestamp 1666199351
transform 1 0 34408 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_365
timestamp 1666199351
transform 1 0 34684 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_369
timestamp 1666199351
transform 1 0 35052 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_381
timestamp 1666199351
transform 1 0 36156 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_387
timestamp 1666199351
transform 1 0 36708 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_404
timestamp 1666199351
transform 1 0 38272 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_415
timestamp 1666199351
transform 1 0 39284 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_419
timestamp 1666199351
transform 1 0 39652 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_421
timestamp 1666199351
transform 1 0 39836 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_426
timestamp 1666199351
transform 1 0 40296 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_433
timestamp 1666199351
transform 1 0 40940 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_440
timestamp 1666199351
transform 1 0 41584 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_447
timestamp 1666199351
transform 1 0 42228 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_453
timestamp 1666199351
transform 1 0 42780 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_459
timestamp 1666199351
transform 1 0 43332 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_465
timestamp 1666199351
transform 1 0 43884 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_473
timestamp 1666199351
transform 1 0 44620 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_477
timestamp 1666199351
transform 1 0 44988 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_489
timestamp 1666199351
transform 1 0 46092 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_501
timestamp 1666199351
transform 1 0 47196 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_513
timestamp 1666199351
transform 1 0 48300 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1666199351
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1666199351
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1666199351
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1666199351
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1666199351
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1666199351
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_57
timestamp 1666199351
transform 1 0 6348 0 -1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_81_64
timestamp 1666199351
transform 1 0 6992 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_76
timestamp 1666199351
transform 1 0 8096 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_88
timestamp 1666199351
transform 1 0 9200 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_100
timestamp 1666199351
transform 1 0 10304 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_113
timestamp 1666199351
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_125
timestamp 1666199351
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_137
timestamp 1666199351
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_149
timestamp 1666199351
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_161
timestamp 1666199351
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1666199351
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_81_169
timestamp 1666199351
transform 1 0 16652 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_81_178
timestamp 1666199351
transform 1 0 17480 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_185
timestamp 1666199351
transform 1 0 18124 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_192
timestamp 1666199351
transform 1 0 18768 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_199
timestamp 1666199351
transform 1 0 19412 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_209
timestamp 1666199351
transform 1 0 20332 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_222
timestamp 1666199351
transform 1 0 21528 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_225
timestamp 1666199351
transform 1 0 21804 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_237
timestamp 1666199351
transform 1 0 22908 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_243
timestamp 1666199351
transform 1 0 23460 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_256
timestamp 1666199351
transform 1 0 24656 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_265
timestamp 1666199351
transform 1 0 25484 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_278
timestamp 1666199351
transform 1 0 26680 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_281
timestamp 1666199351
transform 1 0 26956 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_290
timestamp 1666199351
transform 1 0 27784 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_299
timestamp 1666199351
transform 1 0 28612 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_311
timestamp 1666199351
transform 1 0 29716 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_325
timestamp 1666199351
transform 1 0 31004 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_334
timestamp 1666199351
transform 1 0 31832 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_337
timestamp 1666199351
transform 1 0 32108 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_346
timestamp 1666199351
transform 1 0 32936 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_353
timestamp 1666199351
transform 1 0 33580 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_366
timestamp 1666199351
transform 1 0 34776 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_373
timestamp 1666199351
transform 1 0 35420 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_387
timestamp 1666199351
transform 1 0 36708 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1666199351
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_81_393
timestamp 1666199351
transform 1 0 37260 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_402
timestamp 1666199351
transform 1 0 38088 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_413
timestamp 1666199351
transform 1 0 39100 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_420
timestamp 1666199351
transform 1 0 39744 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_427
timestamp 1666199351
transform 1 0 40388 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_434
timestamp 1666199351
transform 1 0 41032 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_81_441
timestamp 1666199351
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 1666199351
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_81_449
timestamp 1666199351
transform 1 0 42412 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_81_454
timestamp 1666199351
transform 1 0 42872 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_460
timestamp 1666199351
transform 1 0 43424 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_464
timestamp 1666199351
transform 1 0 43792 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_468
timestamp 1666199351
transform 1 0 44160 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_472
timestamp 1666199351
transform 1 0 44528 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_484
timestamp 1666199351
transform 1 0 45632 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_496
timestamp 1666199351
transform 1 0 46736 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_81_505
timestamp 1666199351
transform 1 0 47564 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_513
timestamp 1666199351
transform 1 0 48300 0 -1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1666199351
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1666199351
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1666199351
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_29
timestamp 1666199351
transform 1 0 3772 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_82_40
timestamp 1666199351
transform 1 0 4784 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_47
timestamp 1666199351
transform 1 0 5428 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_54
timestamp 1666199351
transform 1 0 6072 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_82_57
timestamp 1666199351
transform 1 0 6348 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_82_66
timestamp 1666199351
transform 1 0 7176 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_73
timestamp 1666199351
transform 1 0 7820 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_80
timestamp 1666199351
transform 1 0 8464 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_85
timestamp 1666199351
transform 1 0 8924 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_82_90
timestamp 1666199351
transform 1 0 9384 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_96
timestamp 1666199351
transform 1 0 9936 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_82_100
timestamp 1666199351
transform 1 0 10304 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_106
timestamp 1666199351
transform 1 0 10856 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_110
timestamp 1666199351
transform 1 0 11224 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_82_113
timestamp 1666199351
transform 1 0 11500 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_82_124
timestamp 1666199351
transform 1 0 12512 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_132
timestamp 1666199351
transform 1 0 13248 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_136
timestamp 1666199351
transform 1 0 13616 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_141
timestamp 1666199351
transform 1 0 14076 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_148
timestamp 1666199351
transform 1 0 14720 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_82_159
timestamp 1666199351
transform 1 0 15732 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_166
timestamp 1666199351
transform 1 0 16376 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_169
timestamp 1666199351
transform 1 0 16652 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_173
timestamp 1666199351
transform 1 0 17020 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_180
timestamp 1666199351
transform 1 0 17664 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_187
timestamp 1666199351
transform 1 0 18308 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_194
timestamp 1666199351
transform 1 0 18952 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_197
timestamp 1666199351
transform 1 0 19228 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_82_208
timestamp 1666199351
transform 1 0 20240 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_216
timestamp 1666199351
transform 1 0 20976 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_222
timestamp 1666199351
transform 1 0 21528 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_225
timestamp 1666199351
transform 1 0 21804 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_82_233
timestamp 1666199351
transform 1 0 22540 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_250
timestamp 1666199351
transform 1 0 24104 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_253
timestamp 1666199351
transform 1 0 24380 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_261
timestamp 1666199351
transform 1 0 25116 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_272
timestamp 1666199351
transform 1 0 26128 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_278
timestamp 1666199351
transform 1 0 26680 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_281
timestamp 1666199351
transform 1 0 26956 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_286
timestamp 1666199351
transform 1 0 27416 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_290
timestamp 1666199351
transform 1 0 27784 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_298
timestamp 1666199351
transform 1 0 28520 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_82_305
timestamp 1666199351
transform 1 0 29164 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_82_309
timestamp 1666199351
transform 1 0 29532 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_318
timestamp 1666199351
transform 1 0 30360 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_327
timestamp 1666199351
transform 1 0 31188 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_334
timestamp 1666199351
transform 1 0 31832 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_337
timestamp 1666199351
transform 1 0 32108 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_346
timestamp 1666199351
transform 1 0 32936 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_357
timestamp 1666199351
transform 1 0 33948 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_363
timestamp 1666199351
transform 1 0 34500 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_365
timestamp 1666199351
transform 1 0 34684 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_374
timestamp 1666199351
transform 1 0 35512 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_385
timestamp 1666199351
transform 1 0 36524 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_391
timestamp 1666199351
transform 1 0 37076 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_393
timestamp 1666199351
transform 1 0 37260 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_402
timestamp 1666199351
transform 1 0 38088 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_409
timestamp 1666199351
transform 1 0 38732 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_416
timestamp 1666199351
transform 1 0 39376 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_421
timestamp 1666199351
transform 1 0 39836 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_426
timestamp 1666199351
transform 1 0 40296 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_433
timestamp 1666199351
transform 1 0 40940 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_440
timestamp 1666199351
transform 1 0 41584 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_446
timestamp 1666199351
transform 1 0 42136 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_449
timestamp 1666199351
transform 1 0 42412 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_454
timestamp 1666199351
transform 1 0 42872 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_461
timestamp 1666199351
transform 1 0 43516 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_468
timestamp 1666199351
transform 1 0 44160 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_474
timestamp 1666199351
transform 1 0 44712 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_477
timestamp 1666199351
transform 1 0 44988 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_482
timestamp 1666199351
transform 1 0 45448 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_489
timestamp 1666199351
transform 1 0 46092 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_496
timestamp 1666199351
transform 1 0 46736 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_82_505
timestamp 1666199351
transform 1 0 47564 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_513
timestamp 1666199351
transform 1 0 48300 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1666199351
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1666199351
transform -1 0 48852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1666199351
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1666199351
transform -1 0 48852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1666199351
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1666199351
transform -1 0 48852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1666199351
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1666199351
transform -1 0 48852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1666199351
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1666199351
transform -1 0 48852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1666199351
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1666199351
transform -1 0 48852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1666199351
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1666199351
transform -1 0 48852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1666199351
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1666199351
transform -1 0 48852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1666199351
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1666199351
transform -1 0 48852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1666199351
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1666199351
transform -1 0 48852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1666199351
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1666199351
transform -1 0 48852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1666199351
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1666199351
transform -1 0 48852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1666199351
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1666199351
transform -1 0 48852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1666199351
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1666199351
transform -1 0 48852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1666199351
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1666199351
transform -1 0 48852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1666199351
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1666199351
transform -1 0 48852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1666199351
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1666199351
transform -1 0 48852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1666199351
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1666199351
transform -1 0 48852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1666199351
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1666199351
transform -1 0 48852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1666199351
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1666199351
transform -1 0 48852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1666199351
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1666199351
transform -1 0 48852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1666199351
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1666199351
transform -1 0 48852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1666199351
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1666199351
transform -1 0 48852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1666199351
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1666199351
transform -1 0 48852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1666199351
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1666199351
transform -1 0 48852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1666199351
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1666199351
transform -1 0 48852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1666199351
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1666199351
transform -1 0 48852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1666199351
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1666199351
transform -1 0 48852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1666199351
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1666199351
transform -1 0 48852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1666199351
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1666199351
transform -1 0 48852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1666199351
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1666199351
transform -1 0 48852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1666199351
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1666199351
transform -1 0 48852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1666199351
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1666199351
transform -1 0 48852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1666199351
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1666199351
transform -1 0 48852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1666199351
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1666199351
transform -1 0 48852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1666199351
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1666199351
transform -1 0 48852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1666199351
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1666199351
transform -1 0 48852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1666199351
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1666199351
transform -1 0 48852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1666199351
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1666199351
transform -1 0 48852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1666199351
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1666199351
transform -1 0 48852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1666199351
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1666199351
transform -1 0 48852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1666199351
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1666199351
transform -1 0 48852 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1666199351
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1666199351
transform -1 0 48852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1666199351
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1666199351
transform -1 0 48852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1666199351
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1666199351
transform -1 0 48852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1666199351
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1666199351
transform -1 0 48852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1666199351
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1666199351
transform -1 0 48852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1666199351
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1666199351
transform -1 0 48852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1666199351
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1666199351
transform -1 0 48852 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1666199351
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1666199351
transform -1 0 48852 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1666199351
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1666199351
transform -1 0 48852 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1666199351
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1666199351
transform -1 0 48852 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1666199351
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1666199351
transform -1 0 48852 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1666199351
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1666199351
transform -1 0 48852 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1666199351
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1666199351
transform -1 0 48852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1666199351
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1666199351
transform -1 0 48852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1666199351
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1666199351
transform -1 0 48852 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1666199351
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1666199351
transform -1 0 48852 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1666199351
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1666199351
transform -1 0 48852 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1666199351
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1666199351
transform -1 0 48852 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1666199351
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1666199351
transform -1 0 48852 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1666199351
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1666199351
transform -1 0 48852 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1666199351
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1666199351
transform -1 0 48852 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1666199351
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1666199351
transform -1 0 48852 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1666199351
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1666199351
transform -1 0 48852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1666199351
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1666199351
transform -1 0 48852 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1666199351
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1666199351
transform -1 0 48852 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1666199351
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1666199351
transform -1 0 48852 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1666199351
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1666199351
transform -1 0 48852 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1666199351
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1666199351
transform -1 0 48852 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1666199351
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1666199351
transform -1 0 48852 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1666199351
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1666199351
transform -1 0 48852 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1666199351
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1666199351
transform -1 0 48852 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1666199351
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1666199351
transform -1 0 48852 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1666199351
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1666199351
transform -1 0 48852 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1666199351
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1666199351
transform -1 0 48852 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1666199351
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1666199351
transform -1 0 48852 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1666199351
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1666199351
transform -1 0 48852 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1666199351
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1666199351
transform -1 0 48852 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1666199351
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1666199351
transform -1 0 48852 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1666199351
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1666199351
transform -1 0 48852 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1666199351
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1666199351
transform -1 0 48852 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1666199351
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1666199351
transform -1 0 48852 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1666199351
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1666199351
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1666199351
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1666199351
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1666199351
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1666199351
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1666199351
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1666199351
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1666199351
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1666199351
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1666199351
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1666199351
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1666199351
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1666199351
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1666199351
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1666199351
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1666199351
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1666199351
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1666199351
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1666199351
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1666199351
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1666199351
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1666199351
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1666199351
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1666199351
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1666199351
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1666199351
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1666199351
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1666199351
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1666199351
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1666199351
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1666199351
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1666199351
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1666199351
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1666199351
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1666199351
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1666199351
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1666199351
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1666199351
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1666199351
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1666199351
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1666199351
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1666199351
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1666199351
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1666199351
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1666199351
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1666199351
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1666199351
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1666199351
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1666199351
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1666199351
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1666199351
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1666199351
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1666199351
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1666199351
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1666199351
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1666199351
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1666199351
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1666199351
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1666199351
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1666199351
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1666199351
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1666199351
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1666199351
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1666199351
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1666199351
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1666199351
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1666199351
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1666199351
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1666199351
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1666199351
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1666199351
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1666199351
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1666199351
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1666199351
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1666199351
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1666199351
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1666199351
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1666199351
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1666199351
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1666199351
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1666199351
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1666199351
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1666199351
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1666199351
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1666199351
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1666199351
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1666199351
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1666199351
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1666199351
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1666199351
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1666199351
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1666199351
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1666199351
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1666199351
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1666199351
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1666199351
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1666199351
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1666199351
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1666199351
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1666199351
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1666199351
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1666199351
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1666199351
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1666199351
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1666199351
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1666199351
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1666199351
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1666199351
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1666199351
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1666199351
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1666199351
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1666199351
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1666199351
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1666199351
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1666199351
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1666199351
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1666199351
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1666199351
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1666199351
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1666199351
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1666199351
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1666199351
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1666199351
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1666199351
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1666199351
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1666199351
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1666199351
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1666199351
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1666199351
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1666199351
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1666199351
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1666199351
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1666199351
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1666199351
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1666199351
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1666199351
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1666199351
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1666199351
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1666199351
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1666199351
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1666199351
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1666199351
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1666199351
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1666199351
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1666199351
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1666199351
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1666199351
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1666199351
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1666199351
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1666199351
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1666199351
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1666199351
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1666199351
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1666199351
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1666199351
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1666199351
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1666199351
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1666199351
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1666199351
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1666199351
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1666199351
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1666199351
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1666199351
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1666199351
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1666199351
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1666199351
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1666199351
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1666199351
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1666199351
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1666199351
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1666199351
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1666199351
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1666199351
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1666199351
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1666199351
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1666199351
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1666199351
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1666199351
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1666199351
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1666199351
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1666199351
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1666199351
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1666199351
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1666199351
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1666199351
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1666199351
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1666199351
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1666199351
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1666199351
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1666199351
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1666199351
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1666199351
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1666199351
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1666199351
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1666199351
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1666199351
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1666199351
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1666199351
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1666199351
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1666199351
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1666199351
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1666199351
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1666199351
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1666199351
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1666199351
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1666199351
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1666199351
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1666199351
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1666199351
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1666199351
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1666199351
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1666199351
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1666199351
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1666199351
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1666199351
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1666199351
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1666199351
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1666199351
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1666199351
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1666199351
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1666199351
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1666199351
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1666199351
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1666199351
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1666199351
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1666199351
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1666199351
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1666199351
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1666199351
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1666199351
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1666199351
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1666199351
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1666199351
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1666199351
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1666199351
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1666199351
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1666199351
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1666199351
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1666199351
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1666199351
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1666199351
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1666199351
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1666199351
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1666199351
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1666199351
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1666199351
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1666199351
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1666199351
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1666199351
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1666199351
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1666199351
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1666199351
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1666199351
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1666199351
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1666199351
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1666199351
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1666199351
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1666199351
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1666199351
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1666199351
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1666199351
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1666199351
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1666199351
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1666199351
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1666199351
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1666199351
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1666199351
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1666199351
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1666199351
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1666199351
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1666199351
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1666199351
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1666199351
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1666199351
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1666199351
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1666199351
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1666199351
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1666199351
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1666199351
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1666199351
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1666199351
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1666199351
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1666199351
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1666199351
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1666199351
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1666199351
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1666199351
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1666199351
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1666199351
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1666199351
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1666199351
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1666199351
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1666199351
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1666199351
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1666199351
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1666199351
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1666199351
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1666199351
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1666199351
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1666199351
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1666199351
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1666199351
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1666199351
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1666199351
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1666199351
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1666199351
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1666199351
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1666199351
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1666199351
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1666199351
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1666199351
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1666199351
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1666199351
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1666199351
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1666199351
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1666199351
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1666199351
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1666199351
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1666199351
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1666199351
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1666199351
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1666199351
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1666199351
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1666199351
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1666199351
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1666199351
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1666199351
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1666199351
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1666199351
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1666199351
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1666199351
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1666199351
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1666199351
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1666199351
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1666199351
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1666199351
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1666199351
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1666199351
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1666199351
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1666199351
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1666199351
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1666199351
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1666199351
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1666199351
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1666199351
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1666199351
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1666199351
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1666199351
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1666199351
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1666199351
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1666199351
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1666199351
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1666199351
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1666199351
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1666199351
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1666199351
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1666199351
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1666199351
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1666199351
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1666199351
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1666199351
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1666199351
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1666199351
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1666199351
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1666199351
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1666199351
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1666199351
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1666199351
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1666199351
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1666199351
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1666199351
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1666199351
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1666199351
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1666199351
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1666199351
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1666199351
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1666199351
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1666199351
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1666199351
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1666199351
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1666199351
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1666199351
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1666199351
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1666199351
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1666199351
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1666199351
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1666199351
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1666199351
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1666199351
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1666199351
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1666199351
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1666199351
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1666199351
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1666199351
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1666199351
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1666199351
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1666199351
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1666199351
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1666199351
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1666199351
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1666199351
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1666199351
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1666199351
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1666199351
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1666199351
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1666199351
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1666199351
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1666199351
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1666199351
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1666199351
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1666199351
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1666199351
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1666199351
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1666199351
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1666199351
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1666199351
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1666199351
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1666199351
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1666199351
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1666199351
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1666199351
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1666199351
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1666199351
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1666199351
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1666199351
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1666199351
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1666199351
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1666199351
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1666199351
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1666199351
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1666199351
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1666199351
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1666199351
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1666199351
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1666199351
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1666199351
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1666199351
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1666199351
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1666199351
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1666199351
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1666199351
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1666199351
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1666199351
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1666199351
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1666199351
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1666199351
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1666199351
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1666199351
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1666199351
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1666199351
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1666199351
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1666199351
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1666199351
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1666199351
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1666199351
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1666199351
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1666199351
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1666199351
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1666199351
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1666199351
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1666199351
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1666199351
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1666199351
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1666199351
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1666199351
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1666199351
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1666199351
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1666199351
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1666199351
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1666199351
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1666199351
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1666199351
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1666199351
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1666199351
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1666199351
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1666199351
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1666199351
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1666199351
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1666199351
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1666199351
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1666199351
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1666199351
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1666199351
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1666199351
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1666199351
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1666199351
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1666199351
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1666199351
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1666199351
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1666199351
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1666199351
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1666199351
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1666199351
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1666199351
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1666199351
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1666199351
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1666199351
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1666199351
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1666199351
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1666199351
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1666199351
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1666199351
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1666199351
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1666199351
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1666199351
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1666199351
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1666199351
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1666199351
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1666199351
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1666199351
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1666199351
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1666199351
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1666199351
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1666199351
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1666199351
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1666199351
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1666199351
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1666199351
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1666199351
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1666199351
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1666199351
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1666199351
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1666199351
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1666199351
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1666199351
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1666199351
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1666199351
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1666199351
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1666199351
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1666199351
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1666199351
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1666199351
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1666199351
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1666199351
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1666199351
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1666199351
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1666199351
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1666199351
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1666199351
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1666199351
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1666199351
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1666199351
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1666199351
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1666199351
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1666199351
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1666199351
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1666199351
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1666199351
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1666199351
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1666199351
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1666199351
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1666199351
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1666199351
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1666199351
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1666199351
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1666199351
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1666199351
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1666199351
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1666199351
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1666199351
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1666199351
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1666199351
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1666199351
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1666199351
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1666199351
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1666199351
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1666199351
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1666199351
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1666199351
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1666199351
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1666199351
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1666199351
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1666199351
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1666199351
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1666199351
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1666199351
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1666199351
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1666199351
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1666199351
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1666199351
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1666199351
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1666199351
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1666199351
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1666199351
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1666199351
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1666199351
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1666199351
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1666199351
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1666199351
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1666199351
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1666199351
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1666199351
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1666199351
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1666199351
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1666199351
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1666199351
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1666199351
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1666199351
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1666199351
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1666199351
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1666199351
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1666199351
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1666199351
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1666199351
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1666199351
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1666199351
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1666199351
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1666199351
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1666199351
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1666199351
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1666199351
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1666199351
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1666199351
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1666199351
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1666199351
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1666199351
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1666199351
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1666199351
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1666199351
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1666199351
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1666199351
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1666199351
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1666199351
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1666199351
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1666199351
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1666199351
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1666199351
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1666199351
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1666199351
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1666199351
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1666199351
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1666199351
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1666199351
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1666199351
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1666199351
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1666199351
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1666199351
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1666199351
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1666199351
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1666199351
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1666199351
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1666199351
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1666199351
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1666199351
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1666199351
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1666199351
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1666199351
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1666199351
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1666199351
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1666199351
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1666199351
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1666199351
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1666199351
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1666199351
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1666199351
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1666199351
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1666199351
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1666199351
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1666199351
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1666199351
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1666199351
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1666199351
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1666199351
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1666199351
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1666199351
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1666199351
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1666199351
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1666199351
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1666199351
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1666199351
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1666199351
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1666199351
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1666199351
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1666199351
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1666199351
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1666199351
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1666199351
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1666199351
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1666199351
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1666199351
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1666199351
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1666199351
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1666199351
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1666199351
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1666199351
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1666199351
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1666199351
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1666199351
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1666199351
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1666199351
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1666199351
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1666199351
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1666199351
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1666199351
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1666199351
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1666199351
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1666199351
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1666199351
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1666199351
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1666199351
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1666199351
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1666199351
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1666199351
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1666199351
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1666199351
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1666199351
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1666199351
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1666199351
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1666199351
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1666199351
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1666199351
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1666199351
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1666199351
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1666199351
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1666199351
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1666199351
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1666199351
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1666199351
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1666199351
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1666199351
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1666199351
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1666199351
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1666199351
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1666199351
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1666199351
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1666199351
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1666199351
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1666199351
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1666199351
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1666199351
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1666199351
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1666199351
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1666199351
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1666199351
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1666199351
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1666199351
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1666199351
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1666199351
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1666199351
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1666199351
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1666199351
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1666199351
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1666199351
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1666199351
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1666199351
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1666199351
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1666199351
transform 1 0 6256 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1666199351
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1666199351
transform 1 0 11408 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1666199351
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1666199351
transform 1 0 16560 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1666199351
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1666199351
transform 1 0 21712 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1666199351
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1666199351
transform 1 0 26864 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1666199351
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1666199351
transform 1 0 32016 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1666199351
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1666199351
transform 1 0 37168 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1666199351
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1666199351
transform 1 0 42320 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1666199351
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1666199351
transform 1 0 47472 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _157_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 19872 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _158_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 19780 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _159_
timestamp 1666199351
transform -1 0 26956 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _160_
timestamp 1666199351
transform 1 0 31372 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _161_
timestamp 1666199351
transform -1 0 29900 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _162_
timestamp 1666199351
transform -1 0 29808 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _163_
timestamp 1666199351
transform -1 0 30636 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _164_
timestamp 1666199351
transform -1 0 30636 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _165_
timestamp 1666199351
transform 1 0 28060 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _166_
timestamp 1666199351
transform -1 0 27692 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _167_
timestamp 1666199351
transform 1 0 26772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _168_
timestamp 1666199351
transform -1 0 29256 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _169_
timestamp 1666199351
transform -1 0 24104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _170_
timestamp 1666199351
transform -1 0 25392 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _171_
timestamp 1666199351
transform 1 0 24932 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _172_
timestamp 1666199351
transform 1 0 26772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _173_
timestamp 1666199351
transform 1 0 25484 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _174_
timestamp 1666199351
transform 1 0 22172 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _175_
timestamp 1666199351
transform 1 0 23184 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _176_
timestamp 1666199351
transform 1 0 23460 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _177_
timestamp 1666199351
transform 1 0 23644 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _178_
timestamp 1666199351
transform 1 0 23828 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _179_
timestamp 1666199351
transform 1 0 20056 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _180_
timestamp 1666199351
transform 1 0 20056 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _181_
timestamp 1666199351
transform 1 0 20608 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _182_
timestamp 1666199351
transform 1 0 19780 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _183_
timestamp 1666199351
transform 1 0 22908 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _184_
timestamp 1666199351
transform 1 0 22908 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _185_
timestamp 1666199351
transform 1 0 22264 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _186_
timestamp 1666199351
transform 1 0 19412 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _187_
timestamp 1666199351
transform 1 0 19964 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _188_
timestamp 1666199351
transform 1 0 21068 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _189_
timestamp 1666199351
transform -1 0 18308 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _190_
timestamp 1666199351
transform -1 0 18400 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _191_
timestamp 1666199351
transform 1 0 18676 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _192_
timestamp 1666199351
transform 1 0 19964 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_2  _193_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform -1 0 30360 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_2  _194_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 28520 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _195_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform -1 0 29256 0 -1 45696
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_2  _196_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform -1 0 25484 0 -1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_2  _197_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 29716 0 1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _198_
timestamp 1666199351
transform -1 0 29808 0 -1 44608
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_2  _199_
timestamp 1666199351
transform -1 0 25024 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__nand3b_2  _200_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 27416 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_2  _201_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform -1 0 28336 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_2  _202_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 27968 0 1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_2  _203_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 25852 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__and3_2  _204_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform -1 0 29256 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_2  _205_
timestamp 1666199351
transform 1 0 26036 0 -1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _206_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform -1 0 25116 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _207_
timestamp 1666199351
transform -1 0 25024 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_2  _208_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform -1 0 25300 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _209_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 27876 0 1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _210_
timestamp 1666199351
transform 1 0 23000 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  _211_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 23368 0 1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _212_
timestamp 1666199351
transform -1 0 20976 0 1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _213_
timestamp 1666199351
transform -1 0 39192 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_2  _214_
timestamp 1666199351
transform -1 0 38180 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _215_
timestamp 1666199351
transform -1 0 38272 0 1 45696
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_2  _216_
timestamp 1666199351
transform -1 0 31832 0 -1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_2  _217_
timestamp 1666199351
transform 1 0 37444 0 -1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _218_
timestamp 1666199351
transform -1 0 37996 0 1 44608
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_2  _219_
timestamp 1666199351
transform -1 0 32660 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__nand3b_2  _220_
timestamp 1666199351
transform 1 0 35604 0 1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_2  _221_
timestamp 1666199351
transform 1 0 35880 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_2  _222_
timestamp 1666199351
transform -1 0 36708 0 -1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_2  _223_
timestamp 1666199351
transform -1 0 35236 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__and3_2  _224_
timestamp 1666199351
transform -1 0 36432 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_2  _225_
timestamp 1666199351
transform 1 0 33488 0 -1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _226_
timestamp 1666199351
transform 1 0 32292 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _227_
timestamp 1666199351
transform -1 0 32200 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_2  _228_
timestamp 1666199351
transform -1 0 33028 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _229_
timestamp 1666199351
transform -1 0 39284 0 1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _230_
timestamp 1666199351
transform 1 0 32292 0 -1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  _231_
timestamp 1666199351
transform 1 0 32292 0 1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _232_
timestamp 1666199351
transform -1 0 31188 0 1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_2  _233_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 28980 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_2  _234_
timestamp 1666199351
transform -1 0 23000 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_2  _235_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 22172 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _236_
timestamp 1666199351
transform -1 0 31832 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_2  _237_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 25852 0 -1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_2  _238_
timestamp 1666199351
transform 1 0 25484 0 1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  _239_
timestamp 1666199351
transform 1 0 24564 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _240_
timestamp 1666199351
transform -1 0 35144 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_2  _241_
timestamp 1666199351
transform -1 0 34776 0 -1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_2  _242_
timestamp 1666199351
transform 1 0 35880 0 1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  _243_
timestamp 1666199351
transform 1 0 33304 0 1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _244_
timestamp 1666199351
transform -1 0 20148 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _245_
timestamp 1666199351
transform -1 0 18124 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _246_
timestamp 1666199351
transform -1 0 20332 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _247_
timestamp 1666199351
transform 1 0 19228 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_2  _248_
timestamp 1666199351
transform -1 0 20240 0 1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__or2b_2  _249_
timestamp 1666199351
transform -1 0 27784 0 -1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _250_
timestamp 1666199351
transform 1 0 26404 0 1 43520
box -38 -48 1234 592
use sky130_fd_sc_hd__o21a_2  _251_
timestamp 1666199351
transform 1 0 29716 0 1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_2  _252_
timestamp 1666199351
transform 1 0 27232 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_2  _253_
timestamp 1666199351
transform 1 0 27140 0 -1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_2  _254_
timestamp 1666199351
transform -1 0 35512 0 1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _255_
timestamp 1666199351
transform 1 0 34500 0 -1 44608
box -38 -48 1234 592
use sky130_fd_sc_hd__o21a_2  _256_
timestamp 1666199351
transform 1 0 37444 0 1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_2  _257_
timestamp 1666199351
transform 1 0 35420 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_2  _258_
timestamp 1666199351
transform 1 0 37444 0 -1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _259_
timestamp 1666199351
transform -1 0 22540 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _260_
timestamp 1666199351
transform -1 0 18952 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _261_
timestamp 1666199351
transform -1 0 21896 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _262_
timestamp 1666199351
transform 1 0 18492 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_2  _263_
timestamp 1666199351
transform -1 0 21528 0 -1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_2  _264_
timestamp 1666199351
transform 1 0 26220 0 1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _265_
timestamp 1666199351
transform 1 0 28152 0 -1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_2  _266_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 24748 0 1 43520
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_2  _267_
timestamp 1666199351
transform 1 0 27140 0 -1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _268_
timestamp 1666199351
transform -1 0 25668 0 -1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_2  _269_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 25576 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_2  _270_
timestamp 1666199351
transform 1 0 34868 0 1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _271_
timestamp 1666199351
transform -1 0 34960 0 -1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_2  _272_
timestamp 1666199351
transform 1 0 32568 0 1 44608
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_2  _273_
timestamp 1666199351
transform 1 0 33396 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _274_
timestamp 1666199351
transform 1 0 33764 0 1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_2  _275_
timestamp 1666199351
transform 1 0 33396 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__and2_2  _276_
timestamp 1666199351
transform 1 0 20516 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _277_
timestamp 1666199351
transform 1 0 20792 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _278_
timestamp 1666199351
transform -1 0 22540 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _279_
timestamp 1666199351
transform -1 0 22080 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_2  _280_
timestamp 1666199351
transform 1 0 20516 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_2  _281_
timestamp 1666199351
transform 1 0 23460 0 1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_2  _282_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform -1 0 23920 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _283_
timestamp 1666199351
transform -1 0 24380 0 -1 44608
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_2  _284_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 21068 0 1 46784
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_2  _285_
timestamp 1666199351
transform 1 0 25208 0 1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _286_
timestamp 1666199351
transform 1 0 29716 0 1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _287_
timestamp 1666199351
transform -1 0 22908 0 1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_2  _288_
timestamp 1666199351
transform 1 0 31740 0 1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_2  _289_
timestamp 1666199351
transform -1 0 33396 0 1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _290_
timestamp 1666199351
transform -1 0 31372 0 -1 45696
box -38 -48 1234 592
use sky130_fd_sc_hd__o21a_2  _291_
timestamp 1666199351
transform 1 0 38456 0 -1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_2  _292_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 35788 0 -1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_2  _293_
timestamp 1666199351
transform 1 0 30728 0 1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_2  _294_
timestamp 1666199351
transform 1 0 30084 0 -1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_2  _295_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform -1 0 24656 0 -1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__o32a_2  _296_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 23276 0 1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _297_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform -1 0 41584 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _298_
timestamp 1666199351
transform -1 0 42872 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _299_
timestamp 1666199351
transform -1 0 44160 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _300_
timestamp 1666199351
transform 1 0 44252 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _301_
timestamp 1666199351
transform -1 0 46092 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _302_
timestamp 1666199351
transform 1 0 5796 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _303_
timestamp 1666199351
transform 1 0 6900 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _304_
timestamp 1666199351
transform 1 0 8188 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _305_
timestamp 1666199351
transform -1 0 25668 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _306_
timestamp 1666199351
transform -1 0 27416 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _307_
timestamp 1666199351
transform 1 0 26956 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _308_
timestamp 1666199351
transform -1 0 31004 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _309_
timestamp 1666199351
transform 1 0 28980 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _310_
timestamp 1666199351
transform -1 0 35420 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _311_
timestamp 1666199351
transform 1 0 31372 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _312_
timestamp 1666199351
transform -1 0 38732 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _313_
timestamp 1666199351
transform 1 0 33580 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _314_
timestamp 1666199351
transform -1 0 40296 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _315_
timestamp 1666199351
transform -1 0 40388 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _316_
timestamp 1666199351
transform -1 0 41584 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _317_
timestamp 1666199351
transform -1 0 39836 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _318_
timestamp 1666199351
transform -1 0 40940 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _319_
timestamp 1666199351
transform -1 0 42872 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _320_
timestamp 1666199351
transform -1 0 42228 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _321_
timestamp 1666199351
transform -1 0 43516 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _322_
timestamp 1666199351
transform 1 0 43516 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _323_
timestamp 1666199351
transform -1 0 45448 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _324_
timestamp 1666199351
transform -1 0 46736 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _325_
timestamp 1666199351
transform 1 0 10304 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _326_
timestamp 1666199351
transform 1 0 12144 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _327_
timestamp 1666199351
transform 1 0 10948 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _328_
timestamp 1666199351
transform 1 0 12788 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _329_
timestamp 1666199351
transform 1 0 12236 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _330_
timestamp 1666199351
transform 1 0 13432 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _331_
timestamp 1666199351
transform 1 0 12880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _332_
timestamp 1666199351
transform 1 0 12236 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _333_
timestamp 1666199351
transform 1 0 13524 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _334_
timestamp 1666199351
transform 1 0 12880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _335_
timestamp 1666199351
transform 1 0 14812 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _336_
timestamp 1666199351
transform 1 0 14168 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _337_
timestamp 1666199351
transform 1 0 13524 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _338_
timestamp 1666199351
transform 1 0 14812 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _339_
timestamp 1666199351
transform 1 0 15916 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _340_
timestamp 1666199351
transform 1 0 15456 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _341_
timestamp 1666199351
transform 1 0 14812 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _342_
timestamp 1666199351
transform 1 0 16744 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _343_
timestamp 1666199351
transform 1 0 16100 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _344_
timestamp 1666199351
transform 1 0 15456 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _345_
timestamp 1666199351
transform 1 0 14812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _346_
timestamp 1666199351
transform 1 0 17388 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _347_
timestamp 1666199351
transform 1 0 15456 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _348_
timestamp 1666199351
transform 1 0 16744 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _349_
timestamp 1666199351
transform 1 0 16100 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _350_
timestamp 1666199351
transform 1 0 18032 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _351_
timestamp 1666199351
transform 1 0 19228 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _352_
timestamp 1666199351
transform 1 0 18676 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _353_
timestamp 1666199351
transform 1 0 16100 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _354_
timestamp 1666199351
transform 1 0 17388 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _355_
timestamp 1666199351
transform 1 0 16836 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _356_
timestamp 1666199351
transform 1 0 18032 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _357_
timestamp 1666199351
transform -1 0 30544 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _358_
timestamp 1666199351
transform -1 0 31280 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _359_
timestamp 1666199351
transform -1 0 33212 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _360_
timestamp 1666199351
transform -1 0 32568 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _361_
timestamp 1666199351
transform -1 0 31924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _362_
timestamp 1666199351
transform -1 0 33856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _363_
timestamp 1666199351
transform -1 0 33212 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _364_
timestamp 1666199351
transform -1 0 32568 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _365_
timestamp 1666199351
transform -1 0 33856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _366_
timestamp 1666199351
transform -1 0 33212 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _367_
timestamp 1666199351
transform -1 0 34500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _368_
timestamp 1666199351
transform -1 0 33856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _369_
timestamp 1666199351
transform -1 0 35144 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _370_
timestamp 1666199351
transform -1 0 35144 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _371_
timestamp 1666199351
transform -1 0 35788 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _372_
timestamp 1666199351
transform -1 0 35788 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _373_
timestamp 1666199351
transform -1 0 35144 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _374_
timestamp 1666199351
transform -1 0 36432 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _375_
timestamp 1666199351
transform -1 0 35788 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _376_
timestamp 1666199351
transform -1 0 36432 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _377_
timestamp 1666199351
transform -1 0 37720 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _378_
timestamp 1666199351
transform -1 0 36432 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _379_
timestamp 1666199351
transform -1 0 37720 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _380_
timestamp 1666199351
transform -1 0 37076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _381_
timestamp 1666199351
transform -1 0 38364 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _382_
timestamp 1666199351
transform -1 0 37720 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _383_
timestamp 1666199351
transform -1 0 38364 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _384_
timestamp 1666199351
transform -1 0 39008 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _385_
timestamp 1666199351
transform -1 0 38364 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _386_
timestamp 1666199351
transform -1 0 39008 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _387_
timestamp 1666199351
transform -1 0 39008 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _388_
timestamp 1666199351
transform -1 0 40296 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _389_
timestamp 1666199351
transform -1 0 39652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _390_
timestamp 1666199351
transform -1 0 40296 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _391_
timestamp 1666199351
transform -1 0 40940 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _392_
timestamp 1666199351
transform -1 0 40296 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _393_
timestamp 1666199351
transform -1 0 41584 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _394_
timestamp 1666199351
transform -1 0 40940 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _395_
timestamp 1666199351
transform -1 0 40940 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _396_
timestamp 1666199351
transform -1 0 41584 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _397_
timestamp 1666199351
transform -1 0 41584 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _398_
timestamp 1666199351
transform -1 0 42872 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _399_
timestamp 1666199351
transform -1 0 42228 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _400_
timestamp 1666199351
transform -1 0 43516 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _401_
timestamp 1666199351
transform -1 0 42872 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _402_
timestamp 1666199351
transform -1 0 44160 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _403_
timestamp 1666199351
transform -1 0 43516 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _404_
timestamp 1666199351
transform 1 0 42688 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _405_
timestamp 1666199351
transform -1 0 43608 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _406_
timestamp 1666199351
transform -1 0 44160 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _407_
timestamp 1666199351
transform -1 0 45448 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _408_
timestamp 1666199351
transform -1 0 44804 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _409_
timestamp 1666199351
transform -1 0 46092 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _410_
timestamp 1666199351
transform -1 0 45448 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _411_
timestamp 1666199351
transform -1 0 45448 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _412_
timestamp 1666199351
transform -1 0 46736 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _413_
timestamp 1666199351
transform -1 0 46092 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _414_
timestamp 1666199351
transform -1 0 46092 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _415_
timestamp 1666199351
transform -1 0 46736 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _416_
timestamp 1666199351
transform -1 0 48024 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _417_
timestamp 1666199351
transform -1 0 46736 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _418_
timestamp 1666199351
transform -1 0 47380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _419_
timestamp 1666199351
transform -1 0 48024 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _420_
timestamp 1666199351
transform -1 0 48024 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _421_
timestamp 1666199351
transform 1 0 1932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _422_
timestamp 1666199351
transform 1 0 2576 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _423_
timestamp 1666199351
transform 1 0 2576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _424_
timestamp 1666199351
transform 1 0 3220 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _425_
timestamp 1666199351
transform 1 0 4048 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _426_
timestamp 1666199351
transform 1 0 3220 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _427_
timestamp 1666199351
transform 1 0 3864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _428_
timestamp 1666199351
transform 1 0 4968 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _429_
timestamp 1666199351
transform 1 0 4508 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _430_
timestamp 1666199351
transform 1 0 4508 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _431_
timestamp 1666199351
transform 1 0 5796 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _432_
timestamp 1666199351
transform 1 0 5152 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _433_
timestamp 1666199351
transform 1 0 5796 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _434_
timestamp 1666199351
transform 1 0 6624 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _435_
timestamp 1666199351
transform 1 0 5152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _436_
timestamp 1666199351
transform 1 0 5796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _437_
timestamp 1666199351
transform 1 0 7452 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _438_
timestamp 1666199351
transform 1 0 7084 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _439_
timestamp 1666199351
transform 1 0 7084 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _440_
timestamp 1666199351
transform 1 0 8280 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _441_
timestamp 1666199351
transform 1 0 7728 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _442_
timestamp 1666199351
transform 1 0 8372 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _443_
timestamp 1666199351
transform 1 0 9108 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _444_
timestamp 1666199351
transform 1 0 7728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _445_
timestamp 1666199351
transform 1 0 9016 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _446_
timestamp 1666199351
transform 1 0 9936 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _447_
timestamp 1666199351
transform 1 0 8372 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _448_
timestamp 1666199351
transform 1 0 9660 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _449_
timestamp 1666199351
transform 1 0 10764 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _450_
timestamp 1666199351
transform 1 0 10304 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _451_
timestamp 1666199351
transform 1 0 9660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _452_
timestamp 1666199351
transform 1 0 11500 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _453_
timestamp 1666199351
transform 1 0 10948 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _454_
timestamp 1666199351
transform 1 0 19964 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _455_
timestamp 1666199351
transform 1 0 18676 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _456_
timestamp 1666199351
transform 1 0 17480 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _457_
timestamp 1666199351
transform 1 0 17388 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _458_
timestamp 1666199351
transform 1 0 19504 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _459_
timestamp 1666199351
transform 1 0 19320 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _460_
timestamp 1666199351
transform 1 0 18768 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _461_
timestamp 1666199351
transform 1 0 21712 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _462_
timestamp 1666199351
transform 1 0 21252 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _463_
timestamp 1666199351
transform 1 0 20608 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _464_
timestamp 1666199351
transform 1 0 18676 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _465_
timestamp 1666199351
transform 1 0 19412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _466_
timestamp 1666199351
transform 1 0 20424 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _467_
timestamp 1666199351
transform 1 0 21252 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _468_
timestamp 1666199351
transform 1 0 23828 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _469_
timestamp 1666199351
transform 1 0 22264 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _470_
timestamp 1666199351
transform 1 0 22540 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _471_
timestamp 1666199351
transform -1 0 29992 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _472_
timestamp 1666199351
transform 1 0 24840 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _473_
timestamp 1666199351
transform -1 0 26680 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _474_
timestamp 1666199351
transform -1 0 26036 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _475_
timestamp 1666199351
transform 1 0 26128 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _476_
timestamp 1666199351
transform -1 0 28612 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _477_
timestamp 1666199351
transform -1 0 29164 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _478_
timestamp 1666199351
transform -1 0 27600 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _479_
timestamp 1666199351
transform 1 0 26404 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _480_
timestamp 1666199351
transform -1 0 31004 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _481_
timestamp 1666199351
transform -1 0 31280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _482_
timestamp 1666199351
transform 1 0 28704 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _483_
timestamp 1666199351
transform -1 0 29992 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _484_
timestamp 1666199351
transform -1 0 32568 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _485_
timestamp 1666199351
transform -1 0 31648 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _486_
timestamp 1666199351
transform 1 0 4508 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _487_
timestamp 1666199351
transform 1 0 5152 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _488_
timestamp 1666199351
transform 1 0 6716 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _489_
timestamp 1666199351
transform 1 0 7544 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _490_
timestamp 1666199351
transform -1 0 9384 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _491_
timestamp 1666199351
transform 1 0 10028 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _492_
timestamp 1666199351
transform 1 0 10948 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _493_
timestamp 1666199351
transform 1 0 12236 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _494_
timestamp 1666199351
transform 1 0 13340 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _495_
timestamp 1666199351
transform 1 0 14444 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _496_
timestamp 1666199351
transform 1 0 15456 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _497_
timestamp 1666199351
transform 1 0 16100 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _498_
timestamp 1666199351
transform 1 0 17204 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _499_
timestamp 1666199351
transform 1 0 18032 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _500_
timestamp 1666199351
transform 1 0 17388 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _501_
timestamp 1666199351
transform 1 0 18032 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _502_
timestamp 1666199351
transform 1 0 19136 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _503_
timestamp 1666199351
transform 1 0 18676 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _504_
timestamp 1666199351
transform 1 0 22540 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _505_
timestamp 1666199351
transform 1 0 24564 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _506_
timestamp 1666199351
transform -1 0 29164 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _507_
timestamp 1666199351
transform -1 0 28428 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _508_
timestamp 1666199351
transform -1 0 33580 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _509_
timestamp 1666199351
transform -1 0 31004 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _510_
timestamp 1666199351
transform -1 0 31648 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _511_
timestamp 1666199351
transform -1 0 34408 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _512_
timestamp 1666199351
transform -1 0 39376 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _513_
timestamp 1666199351
transform -1 0 39744 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _514_
timestamp 1666199351
transform -1 0 40940 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _515_
timestamp 1666199351
transform -1 0 40296 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _516_
timestamp 1666199351
transform -1 0 38640 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _517_
timestamp 1666199351
transform -1 0 41032 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _518_
timestamp 1666199351
transform -1 0 41676 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _519_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666199351
transform 1 0 20148 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _520_
timestamp 1666199351
transform 1 0 21068 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _521_
timestamp 1666199351
transform 1 0 20700 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _522_
timestamp 1666199351
transform 1 0 20700 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _523_
timestamp 1666199351
transform 1 0 21528 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _524_
timestamp 1666199351
transform 1 0 22080 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _525_
timestamp 1666199351
transform 1 0 22356 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _526_
timestamp 1666199351
transform 1 0 22356 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _527_
timestamp 1666199351
transform 1 0 22908 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _528_
timestamp 1666199351
transform 1 0 23000 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _529_
timestamp 1666199351
transform 1 0 22816 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _530_
timestamp 1666199351
transform 1 0 24564 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _531_
timestamp 1666199351
transform 1 0 24012 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _532_
timestamp 1666199351
transform 1 0 24104 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _533_
timestamp 1666199351
transform 1 0 24288 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _534_
timestamp 1666199351
transform 1 0 24380 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _535_
timestamp 1666199351
transform 1 0 25116 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _536_
timestamp 1666199351
transform -1 0 26220 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _537_
timestamp 1666199351
transform 1 0 25484 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _538_
timestamp 1666199351
transform -1 0 26404 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _539_
timestamp 1666199351
transform 1 0 25760 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _540_
timestamp 1666199351
transform 1 0 27140 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _541_
timestamp 1666199351
transform -1 0 27968 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _542_
timestamp 1666199351
transform -1 0 27968 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _543_
timestamp 1666199351
transform 1 0 27140 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _544_
timestamp 1666199351
transform 1 0 28336 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _545_
timestamp 1666199351
transform -1 0 28520 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _546_
timestamp 1666199351
transform -1 0 29164 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _547_
timestamp 1666199351
transform -1 0 29256 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _548_
timestamp 1666199351
transform -1 0 29256 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _549_
timestamp 1666199351
transform -1 0 30360 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _550_
timestamp 1666199351
transform -1 0 31004 0 -1 44608
box -38 -48 866 592
<< labels >>
flabel metal2 s 3974 49200 4030 50000 0 FreeSans 224 90 0 0 io_active
port 0 nsew signal input
flabel metal2 s 4342 49200 4398 50000 0 FreeSans 224 90 0 0 io_in[0]
port 1 nsew signal input
flabel metal2 s 15382 49200 15438 50000 0 FreeSans 224 90 0 0 io_in[10]
port 2 nsew signal input
flabel metal2 s 16486 49200 16542 50000 0 FreeSans 224 90 0 0 io_in[11]
port 3 nsew signal input
flabel metal2 s 17590 49200 17646 50000 0 FreeSans 224 90 0 0 io_in[12]
port 4 nsew signal input
flabel metal2 s 18694 49200 18750 50000 0 FreeSans 224 90 0 0 io_in[13]
port 5 nsew signal input
flabel metal2 s 19798 49200 19854 50000 0 FreeSans 224 90 0 0 io_in[14]
port 6 nsew signal input
flabel metal2 s 20902 49200 20958 50000 0 FreeSans 224 90 0 0 io_in[15]
port 7 nsew signal input
flabel metal2 s 22006 49200 22062 50000 0 FreeSans 224 90 0 0 io_in[16]
port 8 nsew signal input
flabel metal2 s 23110 49200 23166 50000 0 FreeSans 224 90 0 0 io_in[17]
port 9 nsew signal input
flabel metal2 s 24214 49200 24270 50000 0 FreeSans 224 90 0 0 io_in[18]
port 10 nsew signal input
flabel metal2 s 25318 49200 25374 50000 0 FreeSans 224 90 0 0 io_in[19]
port 11 nsew signal input
flabel metal2 s 5446 49200 5502 50000 0 FreeSans 224 90 0 0 io_in[1]
port 12 nsew signal input
flabel metal2 s 26422 49200 26478 50000 0 FreeSans 224 90 0 0 io_in[20]
port 13 nsew signal input
flabel metal2 s 27526 49200 27582 50000 0 FreeSans 224 90 0 0 io_in[21]
port 14 nsew signal input
flabel metal2 s 28630 49200 28686 50000 0 FreeSans 224 90 0 0 io_in[22]
port 15 nsew signal input
flabel metal2 s 29734 49200 29790 50000 0 FreeSans 224 90 0 0 io_in[23]
port 16 nsew signal input
flabel metal2 s 30838 49200 30894 50000 0 FreeSans 224 90 0 0 io_in[24]
port 17 nsew signal input
flabel metal2 s 31942 49200 31998 50000 0 FreeSans 224 90 0 0 io_in[25]
port 18 nsew signal input
flabel metal2 s 33046 49200 33102 50000 0 FreeSans 224 90 0 0 io_in[26]
port 19 nsew signal input
flabel metal2 s 34150 49200 34206 50000 0 FreeSans 224 90 0 0 io_in[27]
port 20 nsew signal input
flabel metal2 s 35254 49200 35310 50000 0 FreeSans 224 90 0 0 io_in[28]
port 21 nsew signal input
flabel metal2 s 36358 49200 36414 50000 0 FreeSans 224 90 0 0 io_in[29]
port 22 nsew signal input
flabel metal2 s 6550 49200 6606 50000 0 FreeSans 224 90 0 0 io_in[2]
port 23 nsew signal input
flabel metal2 s 37462 49200 37518 50000 0 FreeSans 224 90 0 0 io_in[30]
port 24 nsew signal input
flabel metal2 s 38566 49200 38622 50000 0 FreeSans 224 90 0 0 io_in[31]
port 25 nsew signal input
flabel metal2 s 39670 49200 39726 50000 0 FreeSans 224 90 0 0 io_in[32]
port 26 nsew signal input
flabel metal2 s 40774 49200 40830 50000 0 FreeSans 224 90 0 0 io_in[33]
port 27 nsew signal input
flabel metal2 s 41878 49200 41934 50000 0 FreeSans 224 90 0 0 io_in[34]
port 28 nsew signal input
flabel metal2 s 42982 49200 43038 50000 0 FreeSans 224 90 0 0 io_in[35]
port 29 nsew signal input
flabel metal2 s 44086 49200 44142 50000 0 FreeSans 224 90 0 0 io_in[36]
port 30 nsew signal input
flabel metal2 s 45190 49200 45246 50000 0 FreeSans 224 90 0 0 io_in[37]
port 31 nsew signal input
flabel metal2 s 7654 49200 7710 50000 0 FreeSans 224 90 0 0 io_in[3]
port 32 nsew signal input
flabel metal2 s 8758 49200 8814 50000 0 FreeSans 224 90 0 0 io_in[4]
port 33 nsew signal input
flabel metal2 s 9862 49200 9918 50000 0 FreeSans 224 90 0 0 io_in[5]
port 34 nsew signal input
flabel metal2 s 10966 49200 11022 50000 0 FreeSans 224 90 0 0 io_in[6]
port 35 nsew signal input
flabel metal2 s 12070 49200 12126 50000 0 FreeSans 224 90 0 0 io_in[7]
port 36 nsew signal input
flabel metal2 s 13174 49200 13230 50000 0 FreeSans 224 90 0 0 io_in[8]
port 37 nsew signal input
flabel metal2 s 14278 49200 14334 50000 0 FreeSans 224 90 0 0 io_in[9]
port 38 nsew signal input
flabel metal2 s 4710 49200 4766 50000 0 FreeSans 224 90 0 0 io_oeb[0]
port 39 nsew signal tristate
flabel metal2 s 15750 49200 15806 50000 0 FreeSans 224 90 0 0 io_oeb[10]
port 40 nsew signal tristate
flabel metal2 s 16854 49200 16910 50000 0 FreeSans 224 90 0 0 io_oeb[11]
port 41 nsew signal tristate
flabel metal2 s 17958 49200 18014 50000 0 FreeSans 224 90 0 0 io_oeb[12]
port 42 nsew signal tristate
flabel metal2 s 19062 49200 19118 50000 0 FreeSans 224 90 0 0 io_oeb[13]
port 43 nsew signal tristate
flabel metal2 s 20166 49200 20222 50000 0 FreeSans 224 90 0 0 io_oeb[14]
port 44 nsew signal tristate
flabel metal2 s 21270 49200 21326 50000 0 FreeSans 224 90 0 0 io_oeb[15]
port 45 nsew signal tristate
flabel metal2 s 22374 49200 22430 50000 0 FreeSans 224 90 0 0 io_oeb[16]
port 46 nsew signal tristate
flabel metal2 s 23478 49200 23534 50000 0 FreeSans 224 90 0 0 io_oeb[17]
port 47 nsew signal tristate
flabel metal2 s 24582 49200 24638 50000 0 FreeSans 224 90 0 0 io_oeb[18]
port 48 nsew signal tristate
flabel metal2 s 25686 49200 25742 50000 0 FreeSans 224 90 0 0 io_oeb[19]
port 49 nsew signal tristate
flabel metal2 s 5814 49200 5870 50000 0 FreeSans 224 90 0 0 io_oeb[1]
port 50 nsew signal tristate
flabel metal2 s 26790 49200 26846 50000 0 FreeSans 224 90 0 0 io_oeb[20]
port 51 nsew signal tristate
flabel metal2 s 27894 49200 27950 50000 0 FreeSans 224 90 0 0 io_oeb[21]
port 52 nsew signal tristate
flabel metal2 s 28998 49200 29054 50000 0 FreeSans 224 90 0 0 io_oeb[22]
port 53 nsew signal tristate
flabel metal2 s 30102 49200 30158 50000 0 FreeSans 224 90 0 0 io_oeb[23]
port 54 nsew signal tristate
flabel metal2 s 31206 49200 31262 50000 0 FreeSans 224 90 0 0 io_oeb[24]
port 55 nsew signal tristate
flabel metal2 s 32310 49200 32366 50000 0 FreeSans 224 90 0 0 io_oeb[25]
port 56 nsew signal tristate
flabel metal2 s 33414 49200 33470 50000 0 FreeSans 224 90 0 0 io_oeb[26]
port 57 nsew signal tristate
flabel metal2 s 34518 49200 34574 50000 0 FreeSans 224 90 0 0 io_oeb[27]
port 58 nsew signal tristate
flabel metal2 s 35622 49200 35678 50000 0 FreeSans 224 90 0 0 io_oeb[28]
port 59 nsew signal tristate
flabel metal2 s 36726 49200 36782 50000 0 FreeSans 224 90 0 0 io_oeb[29]
port 60 nsew signal tristate
flabel metal2 s 6918 49200 6974 50000 0 FreeSans 224 90 0 0 io_oeb[2]
port 61 nsew signal tristate
flabel metal2 s 37830 49200 37886 50000 0 FreeSans 224 90 0 0 io_oeb[30]
port 62 nsew signal tristate
flabel metal2 s 38934 49200 38990 50000 0 FreeSans 224 90 0 0 io_oeb[31]
port 63 nsew signal tristate
flabel metal2 s 40038 49200 40094 50000 0 FreeSans 224 90 0 0 io_oeb[32]
port 64 nsew signal tristate
flabel metal2 s 41142 49200 41198 50000 0 FreeSans 224 90 0 0 io_oeb[33]
port 65 nsew signal tristate
flabel metal2 s 42246 49200 42302 50000 0 FreeSans 224 90 0 0 io_oeb[34]
port 66 nsew signal tristate
flabel metal2 s 43350 49200 43406 50000 0 FreeSans 224 90 0 0 io_oeb[35]
port 67 nsew signal tristate
flabel metal2 s 44454 49200 44510 50000 0 FreeSans 224 90 0 0 io_oeb[36]
port 68 nsew signal tristate
flabel metal2 s 45558 49200 45614 50000 0 FreeSans 224 90 0 0 io_oeb[37]
port 69 nsew signal tristate
flabel metal2 s 8022 49200 8078 50000 0 FreeSans 224 90 0 0 io_oeb[3]
port 70 nsew signal tristate
flabel metal2 s 9126 49200 9182 50000 0 FreeSans 224 90 0 0 io_oeb[4]
port 71 nsew signal tristate
flabel metal2 s 10230 49200 10286 50000 0 FreeSans 224 90 0 0 io_oeb[5]
port 72 nsew signal tristate
flabel metal2 s 11334 49200 11390 50000 0 FreeSans 224 90 0 0 io_oeb[6]
port 73 nsew signal tristate
flabel metal2 s 12438 49200 12494 50000 0 FreeSans 224 90 0 0 io_oeb[7]
port 74 nsew signal tristate
flabel metal2 s 13542 49200 13598 50000 0 FreeSans 224 90 0 0 io_oeb[8]
port 75 nsew signal tristate
flabel metal2 s 14646 49200 14702 50000 0 FreeSans 224 90 0 0 io_oeb[9]
port 76 nsew signal tristate
flabel metal2 s 5078 49200 5134 50000 0 FreeSans 224 90 0 0 io_out[0]
port 77 nsew signal tristate
flabel metal2 s 16118 49200 16174 50000 0 FreeSans 224 90 0 0 io_out[10]
port 78 nsew signal tristate
flabel metal2 s 17222 49200 17278 50000 0 FreeSans 224 90 0 0 io_out[11]
port 79 nsew signal tristate
flabel metal2 s 18326 49200 18382 50000 0 FreeSans 224 90 0 0 io_out[12]
port 80 nsew signal tristate
flabel metal2 s 19430 49200 19486 50000 0 FreeSans 224 90 0 0 io_out[13]
port 81 nsew signal tristate
flabel metal2 s 20534 49200 20590 50000 0 FreeSans 224 90 0 0 io_out[14]
port 82 nsew signal tristate
flabel metal2 s 21638 49200 21694 50000 0 FreeSans 224 90 0 0 io_out[15]
port 83 nsew signal tristate
flabel metal2 s 22742 49200 22798 50000 0 FreeSans 224 90 0 0 io_out[16]
port 84 nsew signal tristate
flabel metal2 s 23846 49200 23902 50000 0 FreeSans 224 90 0 0 io_out[17]
port 85 nsew signal tristate
flabel metal2 s 24950 49200 25006 50000 0 FreeSans 224 90 0 0 io_out[18]
port 86 nsew signal tristate
flabel metal2 s 26054 49200 26110 50000 0 FreeSans 224 90 0 0 io_out[19]
port 87 nsew signal tristate
flabel metal2 s 6182 49200 6238 50000 0 FreeSans 224 90 0 0 io_out[1]
port 88 nsew signal tristate
flabel metal2 s 27158 49200 27214 50000 0 FreeSans 224 90 0 0 io_out[20]
port 89 nsew signal tristate
flabel metal2 s 28262 49200 28318 50000 0 FreeSans 224 90 0 0 io_out[21]
port 90 nsew signal tristate
flabel metal2 s 29366 49200 29422 50000 0 FreeSans 224 90 0 0 io_out[22]
port 91 nsew signal tristate
flabel metal2 s 30470 49200 30526 50000 0 FreeSans 224 90 0 0 io_out[23]
port 92 nsew signal tristate
flabel metal2 s 31574 49200 31630 50000 0 FreeSans 224 90 0 0 io_out[24]
port 93 nsew signal tristate
flabel metal2 s 32678 49200 32734 50000 0 FreeSans 224 90 0 0 io_out[25]
port 94 nsew signal tristate
flabel metal2 s 33782 49200 33838 50000 0 FreeSans 224 90 0 0 io_out[26]
port 95 nsew signal tristate
flabel metal2 s 34886 49200 34942 50000 0 FreeSans 224 90 0 0 io_out[27]
port 96 nsew signal tristate
flabel metal2 s 35990 49200 36046 50000 0 FreeSans 224 90 0 0 io_out[28]
port 97 nsew signal tristate
flabel metal2 s 37094 49200 37150 50000 0 FreeSans 224 90 0 0 io_out[29]
port 98 nsew signal tristate
flabel metal2 s 7286 49200 7342 50000 0 FreeSans 224 90 0 0 io_out[2]
port 99 nsew signal tristate
flabel metal2 s 38198 49200 38254 50000 0 FreeSans 224 90 0 0 io_out[30]
port 100 nsew signal tristate
flabel metal2 s 39302 49200 39358 50000 0 FreeSans 224 90 0 0 io_out[31]
port 101 nsew signal tristate
flabel metal2 s 40406 49200 40462 50000 0 FreeSans 224 90 0 0 io_out[32]
port 102 nsew signal tristate
flabel metal2 s 41510 49200 41566 50000 0 FreeSans 224 90 0 0 io_out[33]
port 103 nsew signal tristate
flabel metal2 s 42614 49200 42670 50000 0 FreeSans 224 90 0 0 io_out[34]
port 104 nsew signal tristate
flabel metal2 s 43718 49200 43774 50000 0 FreeSans 224 90 0 0 io_out[35]
port 105 nsew signal tristate
flabel metal2 s 44822 49200 44878 50000 0 FreeSans 224 90 0 0 io_out[36]
port 106 nsew signal tristate
flabel metal2 s 45926 49200 45982 50000 0 FreeSans 224 90 0 0 io_out[37]
port 107 nsew signal tristate
flabel metal2 s 8390 49200 8446 50000 0 FreeSans 224 90 0 0 io_out[3]
port 108 nsew signal tristate
flabel metal2 s 9494 49200 9550 50000 0 FreeSans 224 90 0 0 io_out[4]
port 109 nsew signal tristate
flabel metal2 s 10598 49200 10654 50000 0 FreeSans 224 90 0 0 io_out[5]
port 110 nsew signal tristate
flabel metal2 s 11702 49200 11758 50000 0 FreeSans 224 90 0 0 io_out[6]
port 111 nsew signal tristate
flabel metal2 s 12806 49200 12862 50000 0 FreeSans 224 90 0 0 io_out[7]
port 112 nsew signal tristate
flabel metal2 s 13910 49200 13966 50000 0 FreeSans 224 90 0 0 io_out[8]
port 113 nsew signal tristate
flabel metal2 s 15014 49200 15070 50000 0 FreeSans 224 90 0 0 io_out[9]
port 114 nsew signal tristate
flabel metal2 s 12162 0 12218 800 0 FreeSans 224 90 0 0 la_data_in[0]
port 115 nsew signal input
flabel metal2 s 39762 0 39818 800 0 FreeSans 224 90 0 0 la_data_in[100]
port 116 nsew signal input
flabel metal2 s 40038 0 40094 800 0 FreeSans 224 90 0 0 la_data_in[101]
port 117 nsew signal input
flabel metal2 s 40314 0 40370 800 0 FreeSans 224 90 0 0 la_data_in[102]
port 118 nsew signal input
flabel metal2 s 40590 0 40646 800 0 FreeSans 224 90 0 0 la_data_in[103]
port 119 nsew signal input
flabel metal2 s 40866 0 40922 800 0 FreeSans 224 90 0 0 la_data_in[104]
port 120 nsew signal input
flabel metal2 s 41142 0 41198 800 0 FreeSans 224 90 0 0 la_data_in[105]
port 121 nsew signal input
flabel metal2 s 41418 0 41474 800 0 FreeSans 224 90 0 0 la_data_in[106]
port 122 nsew signal input
flabel metal2 s 41694 0 41750 800 0 FreeSans 224 90 0 0 la_data_in[107]
port 123 nsew signal input
flabel metal2 s 41970 0 42026 800 0 FreeSans 224 90 0 0 la_data_in[108]
port 124 nsew signal input
flabel metal2 s 42246 0 42302 800 0 FreeSans 224 90 0 0 la_data_in[109]
port 125 nsew signal input
flabel metal2 s 14922 0 14978 800 0 FreeSans 224 90 0 0 la_data_in[10]
port 126 nsew signal input
flabel metal2 s 42522 0 42578 800 0 FreeSans 224 90 0 0 la_data_in[110]
port 127 nsew signal input
flabel metal2 s 42798 0 42854 800 0 FreeSans 224 90 0 0 la_data_in[111]
port 128 nsew signal input
flabel metal2 s 43074 0 43130 800 0 FreeSans 224 90 0 0 la_data_in[112]
port 129 nsew signal input
flabel metal2 s 43350 0 43406 800 0 FreeSans 224 90 0 0 la_data_in[113]
port 130 nsew signal input
flabel metal2 s 43626 0 43682 800 0 FreeSans 224 90 0 0 la_data_in[114]
port 131 nsew signal input
flabel metal2 s 43902 0 43958 800 0 FreeSans 224 90 0 0 la_data_in[115]
port 132 nsew signal input
flabel metal2 s 44178 0 44234 800 0 FreeSans 224 90 0 0 la_data_in[116]
port 133 nsew signal input
flabel metal2 s 44454 0 44510 800 0 FreeSans 224 90 0 0 la_data_in[117]
port 134 nsew signal input
flabel metal2 s 44730 0 44786 800 0 FreeSans 224 90 0 0 la_data_in[118]
port 135 nsew signal input
flabel metal2 s 45006 0 45062 800 0 FreeSans 224 90 0 0 la_data_in[119]
port 136 nsew signal input
flabel metal2 s 15198 0 15254 800 0 FreeSans 224 90 0 0 la_data_in[11]
port 137 nsew signal input
flabel metal2 s 45282 0 45338 800 0 FreeSans 224 90 0 0 la_data_in[120]
port 138 nsew signal input
flabel metal2 s 45558 0 45614 800 0 FreeSans 224 90 0 0 la_data_in[121]
port 139 nsew signal input
flabel metal2 s 45834 0 45890 800 0 FreeSans 224 90 0 0 la_data_in[122]
port 140 nsew signal input
flabel metal2 s 46110 0 46166 800 0 FreeSans 224 90 0 0 la_data_in[123]
port 141 nsew signal input
flabel metal2 s 46386 0 46442 800 0 FreeSans 224 90 0 0 la_data_in[124]
port 142 nsew signal input
flabel metal2 s 46662 0 46718 800 0 FreeSans 224 90 0 0 la_data_in[125]
port 143 nsew signal input
flabel metal2 s 46938 0 46994 800 0 FreeSans 224 90 0 0 la_data_in[126]
port 144 nsew signal input
flabel metal2 s 47214 0 47270 800 0 FreeSans 224 90 0 0 la_data_in[127]
port 145 nsew signal input
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 la_data_in[12]
port 146 nsew signal input
flabel metal2 s 15750 0 15806 800 0 FreeSans 224 90 0 0 la_data_in[13]
port 147 nsew signal input
flabel metal2 s 16026 0 16082 800 0 FreeSans 224 90 0 0 la_data_in[14]
port 148 nsew signal input
flabel metal2 s 16302 0 16358 800 0 FreeSans 224 90 0 0 la_data_in[15]
port 149 nsew signal input
flabel metal2 s 16578 0 16634 800 0 FreeSans 224 90 0 0 la_data_in[16]
port 150 nsew signal input
flabel metal2 s 16854 0 16910 800 0 FreeSans 224 90 0 0 la_data_in[17]
port 151 nsew signal input
flabel metal2 s 17130 0 17186 800 0 FreeSans 224 90 0 0 la_data_in[18]
port 152 nsew signal input
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 la_data_in[19]
port 153 nsew signal input
flabel metal2 s 12438 0 12494 800 0 FreeSans 224 90 0 0 la_data_in[1]
port 154 nsew signal input
flabel metal2 s 17682 0 17738 800 0 FreeSans 224 90 0 0 la_data_in[20]
port 155 nsew signal input
flabel metal2 s 17958 0 18014 800 0 FreeSans 224 90 0 0 la_data_in[21]
port 156 nsew signal input
flabel metal2 s 18234 0 18290 800 0 FreeSans 224 90 0 0 la_data_in[22]
port 157 nsew signal input
flabel metal2 s 18510 0 18566 800 0 FreeSans 224 90 0 0 la_data_in[23]
port 158 nsew signal input
flabel metal2 s 18786 0 18842 800 0 FreeSans 224 90 0 0 la_data_in[24]
port 159 nsew signal input
flabel metal2 s 19062 0 19118 800 0 FreeSans 224 90 0 0 la_data_in[25]
port 160 nsew signal input
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 la_data_in[26]
port 161 nsew signal input
flabel metal2 s 19614 0 19670 800 0 FreeSans 224 90 0 0 la_data_in[27]
port 162 nsew signal input
flabel metal2 s 19890 0 19946 800 0 FreeSans 224 90 0 0 la_data_in[28]
port 163 nsew signal input
flabel metal2 s 20166 0 20222 800 0 FreeSans 224 90 0 0 la_data_in[29]
port 164 nsew signal input
flabel metal2 s 12714 0 12770 800 0 FreeSans 224 90 0 0 la_data_in[2]
port 165 nsew signal input
flabel metal2 s 20442 0 20498 800 0 FreeSans 224 90 0 0 la_data_in[30]
port 166 nsew signal input
flabel metal2 s 20718 0 20774 800 0 FreeSans 224 90 0 0 la_data_in[31]
port 167 nsew signal input
flabel metal2 s 20994 0 21050 800 0 FreeSans 224 90 0 0 la_data_in[32]
port 168 nsew signal input
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 la_data_in[33]
port 169 nsew signal input
flabel metal2 s 21546 0 21602 800 0 FreeSans 224 90 0 0 la_data_in[34]
port 170 nsew signal input
flabel metal2 s 21822 0 21878 800 0 FreeSans 224 90 0 0 la_data_in[35]
port 171 nsew signal input
flabel metal2 s 22098 0 22154 800 0 FreeSans 224 90 0 0 la_data_in[36]
port 172 nsew signal input
flabel metal2 s 22374 0 22430 800 0 FreeSans 224 90 0 0 la_data_in[37]
port 173 nsew signal input
flabel metal2 s 22650 0 22706 800 0 FreeSans 224 90 0 0 la_data_in[38]
port 174 nsew signal input
flabel metal2 s 22926 0 22982 800 0 FreeSans 224 90 0 0 la_data_in[39]
port 175 nsew signal input
flabel metal2 s 12990 0 13046 800 0 FreeSans 224 90 0 0 la_data_in[3]
port 176 nsew signal input
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 la_data_in[40]
port 177 nsew signal input
flabel metal2 s 23478 0 23534 800 0 FreeSans 224 90 0 0 la_data_in[41]
port 178 nsew signal input
flabel metal2 s 23754 0 23810 800 0 FreeSans 224 90 0 0 la_data_in[42]
port 179 nsew signal input
flabel metal2 s 24030 0 24086 800 0 FreeSans 224 90 0 0 la_data_in[43]
port 180 nsew signal input
flabel metal2 s 24306 0 24362 800 0 FreeSans 224 90 0 0 la_data_in[44]
port 181 nsew signal input
flabel metal2 s 24582 0 24638 800 0 FreeSans 224 90 0 0 la_data_in[45]
port 182 nsew signal input
flabel metal2 s 24858 0 24914 800 0 FreeSans 224 90 0 0 la_data_in[46]
port 183 nsew signal input
flabel metal2 s 25134 0 25190 800 0 FreeSans 224 90 0 0 la_data_in[47]
port 184 nsew signal input
flabel metal2 s 25410 0 25466 800 0 FreeSans 224 90 0 0 la_data_in[48]
port 185 nsew signal input
flabel metal2 s 25686 0 25742 800 0 FreeSans 224 90 0 0 la_data_in[49]
port 186 nsew signal input
flabel metal2 s 13266 0 13322 800 0 FreeSans 224 90 0 0 la_data_in[4]
port 187 nsew signal input
flabel metal2 s 25962 0 26018 800 0 FreeSans 224 90 0 0 la_data_in[50]
port 188 nsew signal input
flabel metal2 s 26238 0 26294 800 0 FreeSans 224 90 0 0 la_data_in[51]
port 189 nsew signal input
flabel metal2 s 26514 0 26570 800 0 FreeSans 224 90 0 0 la_data_in[52]
port 190 nsew signal input
flabel metal2 s 26790 0 26846 800 0 FreeSans 224 90 0 0 la_data_in[53]
port 191 nsew signal input
flabel metal2 s 27066 0 27122 800 0 FreeSans 224 90 0 0 la_data_in[54]
port 192 nsew signal input
flabel metal2 s 27342 0 27398 800 0 FreeSans 224 90 0 0 la_data_in[55]
port 193 nsew signal input
flabel metal2 s 27618 0 27674 800 0 FreeSans 224 90 0 0 la_data_in[56]
port 194 nsew signal input
flabel metal2 s 27894 0 27950 800 0 FreeSans 224 90 0 0 la_data_in[57]
port 195 nsew signal input
flabel metal2 s 28170 0 28226 800 0 FreeSans 224 90 0 0 la_data_in[58]
port 196 nsew signal input
flabel metal2 s 28446 0 28502 800 0 FreeSans 224 90 0 0 la_data_in[59]
port 197 nsew signal input
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 la_data_in[5]
port 198 nsew signal input
flabel metal2 s 28722 0 28778 800 0 FreeSans 224 90 0 0 la_data_in[60]
port 199 nsew signal input
flabel metal2 s 28998 0 29054 800 0 FreeSans 224 90 0 0 la_data_in[61]
port 200 nsew signal input
flabel metal2 s 29274 0 29330 800 0 FreeSans 224 90 0 0 la_data_in[62]
port 201 nsew signal input
flabel metal2 s 29550 0 29606 800 0 FreeSans 224 90 0 0 la_data_in[63]
port 202 nsew signal input
flabel metal2 s 29826 0 29882 800 0 FreeSans 224 90 0 0 la_data_in[64]
port 203 nsew signal input
flabel metal2 s 30102 0 30158 800 0 FreeSans 224 90 0 0 la_data_in[65]
port 204 nsew signal input
flabel metal2 s 30378 0 30434 800 0 FreeSans 224 90 0 0 la_data_in[66]
port 205 nsew signal input
flabel metal2 s 30654 0 30710 800 0 FreeSans 224 90 0 0 la_data_in[67]
port 206 nsew signal input
flabel metal2 s 30930 0 30986 800 0 FreeSans 224 90 0 0 la_data_in[68]
port 207 nsew signal input
flabel metal2 s 31206 0 31262 800 0 FreeSans 224 90 0 0 la_data_in[69]
port 208 nsew signal input
flabel metal2 s 13818 0 13874 800 0 FreeSans 224 90 0 0 la_data_in[6]
port 209 nsew signal input
flabel metal2 s 31482 0 31538 800 0 FreeSans 224 90 0 0 la_data_in[70]
port 210 nsew signal input
flabel metal2 s 31758 0 31814 800 0 FreeSans 224 90 0 0 la_data_in[71]
port 211 nsew signal input
flabel metal2 s 32034 0 32090 800 0 FreeSans 224 90 0 0 la_data_in[72]
port 212 nsew signal input
flabel metal2 s 32310 0 32366 800 0 FreeSans 224 90 0 0 la_data_in[73]
port 213 nsew signal input
flabel metal2 s 32586 0 32642 800 0 FreeSans 224 90 0 0 la_data_in[74]
port 214 nsew signal input
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 la_data_in[75]
port 215 nsew signal input
flabel metal2 s 33138 0 33194 800 0 FreeSans 224 90 0 0 la_data_in[76]
port 216 nsew signal input
flabel metal2 s 33414 0 33470 800 0 FreeSans 224 90 0 0 la_data_in[77]
port 217 nsew signal input
flabel metal2 s 33690 0 33746 800 0 FreeSans 224 90 0 0 la_data_in[78]
port 218 nsew signal input
flabel metal2 s 33966 0 34022 800 0 FreeSans 224 90 0 0 la_data_in[79]
port 219 nsew signal input
flabel metal2 s 14094 0 14150 800 0 FreeSans 224 90 0 0 la_data_in[7]
port 220 nsew signal input
flabel metal2 s 34242 0 34298 800 0 FreeSans 224 90 0 0 la_data_in[80]
port 221 nsew signal input
flabel metal2 s 34518 0 34574 800 0 FreeSans 224 90 0 0 la_data_in[81]
port 222 nsew signal input
flabel metal2 s 34794 0 34850 800 0 FreeSans 224 90 0 0 la_data_in[82]
port 223 nsew signal input
flabel metal2 s 35070 0 35126 800 0 FreeSans 224 90 0 0 la_data_in[83]
port 224 nsew signal input
flabel metal2 s 35346 0 35402 800 0 FreeSans 224 90 0 0 la_data_in[84]
port 225 nsew signal input
flabel metal2 s 35622 0 35678 800 0 FreeSans 224 90 0 0 la_data_in[85]
port 226 nsew signal input
flabel metal2 s 35898 0 35954 800 0 FreeSans 224 90 0 0 la_data_in[86]
port 227 nsew signal input
flabel metal2 s 36174 0 36230 800 0 FreeSans 224 90 0 0 la_data_in[87]
port 228 nsew signal input
flabel metal2 s 36450 0 36506 800 0 FreeSans 224 90 0 0 la_data_in[88]
port 229 nsew signal input
flabel metal2 s 36726 0 36782 800 0 FreeSans 224 90 0 0 la_data_in[89]
port 230 nsew signal input
flabel metal2 s 14370 0 14426 800 0 FreeSans 224 90 0 0 la_data_in[8]
port 231 nsew signal input
flabel metal2 s 37002 0 37058 800 0 FreeSans 224 90 0 0 la_data_in[90]
port 232 nsew signal input
flabel metal2 s 37278 0 37334 800 0 FreeSans 224 90 0 0 la_data_in[91]
port 233 nsew signal input
flabel metal2 s 37554 0 37610 800 0 FreeSans 224 90 0 0 la_data_in[92]
port 234 nsew signal input
flabel metal2 s 37830 0 37886 800 0 FreeSans 224 90 0 0 la_data_in[93]
port 235 nsew signal input
flabel metal2 s 38106 0 38162 800 0 FreeSans 224 90 0 0 la_data_in[94]
port 236 nsew signal input
flabel metal2 s 38382 0 38438 800 0 FreeSans 224 90 0 0 la_data_in[95]
port 237 nsew signal input
flabel metal2 s 38658 0 38714 800 0 FreeSans 224 90 0 0 la_data_in[96]
port 238 nsew signal input
flabel metal2 s 38934 0 38990 800 0 FreeSans 224 90 0 0 la_data_in[97]
port 239 nsew signal input
flabel metal2 s 39210 0 39266 800 0 FreeSans 224 90 0 0 la_data_in[98]
port 240 nsew signal input
flabel metal2 s 39486 0 39542 800 0 FreeSans 224 90 0 0 la_data_in[99]
port 241 nsew signal input
flabel metal2 s 14646 0 14702 800 0 FreeSans 224 90 0 0 la_data_in[9]
port 242 nsew signal input
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 la_data_out[0]
port 243 nsew signal tristate
flabel metal2 s 39854 0 39910 800 0 FreeSans 224 90 0 0 la_data_out[100]
port 244 nsew signal tristate
flabel metal2 s 40130 0 40186 800 0 FreeSans 224 90 0 0 la_data_out[101]
port 245 nsew signal tristate
flabel metal2 s 40406 0 40462 800 0 FreeSans 224 90 0 0 la_data_out[102]
port 246 nsew signal tristate
flabel metal2 s 40682 0 40738 800 0 FreeSans 224 90 0 0 la_data_out[103]
port 247 nsew signal tristate
flabel metal2 s 40958 0 41014 800 0 FreeSans 224 90 0 0 la_data_out[104]
port 248 nsew signal tristate
flabel metal2 s 41234 0 41290 800 0 FreeSans 224 90 0 0 la_data_out[105]
port 249 nsew signal tristate
flabel metal2 s 41510 0 41566 800 0 FreeSans 224 90 0 0 la_data_out[106]
port 250 nsew signal tristate
flabel metal2 s 41786 0 41842 800 0 FreeSans 224 90 0 0 la_data_out[107]
port 251 nsew signal tristate
flabel metal2 s 42062 0 42118 800 0 FreeSans 224 90 0 0 la_data_out[108]
port 252 nsew signal tristate
flabel metal2 s 42338 0 42394 800 0 FreeSans 224 90 0 0 la_data_out[109]
port 253 nsew signal tristate
flabel metal2 s 15014 0 15070 800 0 FreeSans 224 90 0 0 la_data_out[10]
port 254 nsew signal tristate
flabel metal2 s 42614 0 42670 800 0 FreeSans 224 90 0 0 la_data_out[110]
port 255 nsew signal tristate
flabel metal2 s 42890 0 42946 800 0 FreeSans 224 90 0 0 la_data_out[111]
port 256 nsew signal tristate
flabel metal2 s 43166 0 43222 800 0 FreeSans 224 90 0 0 la_data_out[112]
port 257 nsew signal tristate
flabel metal2 s 43442 0 43498 800 0 FreeSans 224 90 0 0 la_data_out[113]
port 258 nsew signal tristate
flabel metal2 s 43718 0 43774 800 0 FreeSans 224 90 0 0 la_data_out[114]
port 259 nsew signal tristate
flabel metal2 s 43994 0 44050 800 0 FreeSans 224 90 0 0 la_data_out[115]
port 260 nsew signal tristate
flabel metal2 s 44270 0 44326 800 0 FreeSans 224 90 0 0 la_data_out[116]
port 261 nsew signal tristate
flabel metal2 s 44546 0 44602 800 0 FreeSans 224 90 0 0 la_data_out[117]
port 262 nsew signal tristate
flabel metal2 s 44822 0 44878 800 0 FreeSans 224 90 0 0 la_data_out[118]
port 263 nsew signal tristate
flabel metal2 s 45098 0 45154 800 0 FreeSans 224 90 0 0 la_data_out[119]
port 264 nsew signal tristate
flabel metal2 s 15290 0 15346 800 0 FreeSans 224 90 0 0 la_data_out[11]
port 265 nsew signal tristate
flabel metal2 s 45374 0 45430 800 0 FreeSans 224 90 0 0 la_data_out[120]
port 266 nsew signal tristate
flabel metal2 s 45650 0 45706 800 0 FreeSans 224 90 0 0 la_data_out[121]
port 267 nsew signal tristate
flabel metal2 s 45926 0 45982 800 0 FreeSans 224 90 0 0 la_data_out[122]
port 268 nsew signal tristate
flabel metal2 s 46202 0 46258 800 0 FreeSans 224 90 0 0 la_data_out[123]
port 269 nsew signal tristate
flabel metal2 s 46478 0 46534 800 0 FreeSans 224 90 0 0 la_data_out[124]
port 270 nsew signal tristate
flabel metal2 s 46754 0 46810 800 0 FreeSans 224 90 0 0 la_data_out[125]
port 271 nsew signal tristate
flabel metal2 s 47030 0 47086 800 0 FreeSans 224 90 0 0 la_data_out[126]
port 272 nsew signal tristate
flabel metal2 s 47306 0 47362 800 0 FreeSans 224 90 0 0 la_data_out[127]
port 273 nsew signal tristate
flabel metal2 s 15566 0 15622 800 0 FreeSans 224 90 0 0 la_data_out[12]
port 274 nsew signal tristate
flabel metal2 s 15842 0 15898 800 0 FreeSans 224 90 0 0 la_data_out[13]
port 275 nsew signal tristate
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 la_data_out[14]
port 276 nsew signal tristate
flabel metal2 s 16394 0 16450 800 0 FreeSans 224 90 0 0 la_data_out[15]
port 277 nsew signal tristate
flabel metal2 s 16670 0 16726 800 0 FreeSans 224 90 0 0 la_data_out[16]
port 278 nsew signal tristate
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 la_data_out[17]
port 279 nsew signal tristate
flabel metal2 s 17222 0 17278 800 0 FreeSans 224 90 0 0 la_data_out[18]
port 280 nsew signal tristate
flabel metal2 s 17498 0 17554 800 0 FreeSans 224 90 0 0 la_data_out[19]
port 281 nsew signal tristate
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 la_data_out[1]
port 282 nsew signal tristate
flabel metal2 s 17774 0 17830 800 0 FreeSans 224 90 0 0 la_data_out[20]
port 283 nsew signal tristate
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 la_data_out[21]
port 284 nsew signal tristate
flabel metal2 s 18326 0 18382 800 0 FreeSans 224 90 0 0 la_data_out[22]
port 285 nsew signal tristate
flabel metal2 s 18602 0 18658 800 0 FreeSans 224 90 0 0 la_data_out[23]
port 286 nsew signal tristate
flabel metal2 s 18878 0 18934 800 0 FreeSans 224 90 0 0 la_data_out[24]
port 287 nsew signal tristate
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 la_data_out[25]
port 288 nsew signal tristate
flabel metal2 s 19430 0 19486 800 0 FreeSans 224 90 0 0 la_data_out[26]
port 289 nsew signal tristate
flabel metal2 s 19706 0 19762 800 0 FreeSans 224 90 0 0 la_data_out[27]
port 290 nsew signal tristate
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 la_data_out[28]
port 291 nsew signal tristate
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 la_data_out[29]
port 292 nsew signal tristate
flabel metal2 s 12806 0 12862 800 0 FreeSans 224 90 0 0 la_data_out[2]
port 293 nsew signal tristate
flabel metal2 s 20534 0 20590 800 0 FreeSans 224 90 0 0 la_data_out[30]
port 294 nsew signal tristate
flabel metal2 s 20810 0 20866 800 0 FreeSans 224 90 0 0 la_data_out[31]
port 295 nsew signal tristate
flabel metal2 s 21086 0 21142 800 0 FreeSans 224 90 0 0 la_data_out[32]
port 296 nsew signal tristate
flabel metal2 s 21362 0 21418 800 0 FreeSans 224 90 0 0 la_data_out[33]
port 297 nsew signal tristate
flabel metal2 s 21638 0 21694 800 0 FreeSans 224 90 0 0 la_data_out[34]
port 298 nsew signal tristate
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 la_data_out[35]
port 299 nsew signal tristate
flabel metal2 s 22190 0 22246 800 0 FreeSans 224 90 0 0 la_data_out[36]
port 300 nsew signal tristate
flabel metal2 s 22466 0 22522 800 0 FreeSans 224 90 0 0 la_data_out[37]
port 301 nsew signal tristate
flabel metal2 s 22742 0 22798 800 0 FreeSans 224 90 0 0 la_data_out[38]
port 302 nsew signal tristate
flabel metal2 s 23018 0 23074 800 0 FreeSans 224 90 0 0 la_data_out[39]
port 303 nsew signal tristate
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 la_data_out[3]
port 304 nsew signal tristate
flabel metal2 s 23294 0 23350 800 0 FreeSans 224 90 0 0 la_data_out[40]
port 305 nsew signal tristate
flabel metal2 s 23570 0 23626 800 0 FreeSans 224 90 0 0 la_data_out[41]
port 306 nsew signal tristate
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 la_data_out[42]
port 307 nsew signal tristate
flabel metal2 s 24122 0 24178 800 0 FreeSans 224 90 0 0 la_data_out[43]
port 308 nsew signal tristate
flabel metal2 s 24398 0 24454 800 0 FreeSans 224 90 0 0 la_data_out[44]
port 309 nsew signal tristate
flabel metal2 s 24674 0 24730 800 0 FreeSans 224 90 0 0 la_data_out[45]
port 310 nsew signal tristate
flabel metal2 s 24950 0 25006 800 0 FreeSans 224 90 0 0 la_data_out[46]
port 311 nsew signal tristate
flabel metal2 s 25226 0 25282 800 0 FreeSans 224 90 0 0 la_data_out[47]
port 312 nsew signal tristate
flabel metal2 s 25502 0 25558 800 0 FreeSans 224 90 0 0 la_data_out[48]
port 313 nsew signal tristate
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 la_data_out[49]
port 314 nsew signal tristate
flabel metal2 s 13358 0 13414 800 0 FreeSans 224 90 0 0 la_data_out[4]
port 315 nsew signal tristate
flabel metal2 s 26054 0 26110 800 0 FreeSans 224 90 0 0 la_data_out[50]
port 316 nsew signal tristate
flabel metal2 s 26330 0 26386 800 0 FreeSans 224 90 0 0 la_data_out[51]
port 317 nsew signal tristate
flabel metal2 s 26606 0 26662 800 0 FreeSans 224 90 0 0 la_data_out[52]
port 318 nsew signal tristate
flabel metal2 s 26882 0 26938 800 0 FreeSans 224 90 0 0 la_data_out[53]
port 319 nsew signal tristate
flabel metal2 s 27158 0 27214 800 0 FreeSans 224 90 0 0 la_data_out[54]
port 320 nsew signal tristate
flabel metal2 s 27434 0 27490 800 0 FreeSans 224 90 0 0 la_data_out[55]
port 321 nsew signal tristate
flabel metal2 s 27710 0 27766 800 0 FreeSans 224 90 0 0 la_data_out[56]
port 322 nsew signal tristate
flabel metal2 s 27986 0 28042 800 0 FreeSans 224 90 0 0 la_data_out[57]
port 323 nsew signal tristate
flabel metal2 s 28262 0 28318 800 0 FreeSans 224 90 0 0 la_data_out[58]
port 324 nsew signal tristate
flabel metal2 s 28538 0 28594 800 0 FreeSans 224 90 0 0 la_data_out[59]
port 325 nsew signal tristate
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 la_data_out[5]
port 326 nsew signal tristate
flabel metal2 s 28814 0 28870 800 0 FreeSans 224 90 0 0 la_data_out[60]
port 327 nsew signal tristate
flabel metal2 s 29090 0 29146 800 0 FreeSans 224 90 0 0 la_data_out[61]
port 328 nsew signal tristate
flabel metal2 s 29366 0 29422 800 0 FreeSans 224 90 0 0 la_data_out[62]
port 329 nsew signal tristate
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 la_data_out[63]
port 330 nsew signal tristate
flabel metal2 s 29918 0 29974 800 0 FreeSans 224 90 0 0 la_data_out[64]
port 331 nsew signal tristate
flabel metal2 s 30194 0 30250 800 0 FreeSans 224 90 0 0 la_data_out[65]
port 332 nsew signal tristate
flabel metal2 s 30470 0 30526 800 0 FreeSans 224 90 0 0 la_data_out[66]
port 333 nsew signal tristate
flabel metal2 s 30746 0 30802 800 0 FreeSans 224 90 0 0 la_data_out[67]
port 334 nsew signal tristate
flabel metal2 s 31022 0 31078 800 0 FreeSans 224 90 0 0 la_data_out[68]
port 335 nsew signal tristate
flabel metal2 s 31298 0 31354 800 0 FreeSans 224 90 0 0 la_data_out[69]
port 336 nsew signal tristate
flabel metal2 s 13910 0 13966 800 0 FreeSans 224 90 0 0 la_data_out[6]
port 337 nsew signal tristate
flabel metal2 s 31574 0 31630 800 0 FreeSans 224 90 0 0 la_data_out[70]
port 338 nsew signal tristate
flabel metal2 s 31850 0 31906 800 0 FreeSans 224 90 0 0 la_data_out[71]
port 339 nsew signal tristate
flabel metal2 s 32126 0 32182 800 0 FreeSans 224 90 0 0 la_data_out[72]
port 340 nsew signal tristate
flabel metal2 s 32402 0 32458 800 0 FreeSans 224 90 0 0 la_data_out[73]
port 341 nsew signal tristate
flabel metal2 s 32678 0 32734 800 0 FreeSans 224 90 0 0 la_data_out[74]
port 342 nsew signal tristate
flabel metal2 s 32954 0 33010 800 0 FreeSans 224 90 0 0 la_data_out[75]
port 343 nsew signal tristate
flabel metal2 s 33230 0 33286 800 0 FreeSans 224 90 0 0 la_data_out[76]
port 344 nsew signal tristate
flabel metal2 s 33506 0 33562 800 0 FreeSans 224 90 0 0 la_data_out[77]
port 345 nsew signal tristate
flabel metal2 s 33782 0 33838 800 0 FreeSans 224 90 0 0 la_data_out[78]
port 346 nsew signal tristate
flabel metal2 s 34058 0 34114 800 0 FreeSans 224 90 0 0 la_data_out[79]
port 347 nsew signal tristate
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 la_data_out[7]
port 348 nsew signal tristate
flabel metal2 s 34334 0 34390 800 0 FreeSans 224 90 0 0 la_data_out[80]
port 349 nsew signal tristate
flabel metal2 s 34610 0 34666 800 0 FreeSans 224 90 0 0 la_data_out[81]
port 350 nsew signal tristate
flabel metal2 s 34886 0 34942 800 0 FreeSans 224 90 0 0 la_data_out[82]
port 351 nsew signal tristate
flabel metal2 s 35162 0 35218 800 0 FreeSans 224 90 0 0 la_data_out[83]
port 352 nsew signal tristate
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 la_data_out[84]
port 353 nsew signal tristate
flabel metal2 s 35714 0 35770 800 0 FreeSans 224 90 0 0 la_data_out[85]
port 354 nsew signal tristate
flabel metal2 s 35990 0 36046 800 0 FreeSans 224 90 0 0 la_data_out[86]
port 355 nsew signal tristate
flabel metal2 s 36266 0 36322 800 0 FreeSans 224 90 0 0 la_data_out[87]
port 356 nsew signal tristate
flabel metal2 s 36542 0 36598 800 0 FreeSans 224 90 0 0 la_data_out[88]
port 357 nsew signal tristate
flabel metal2 s 36818 0 36874 800 0 FreeSans 224 90 0 0 la_data_out[89]
port 358 nsew signal tristate
flabel metal2 s 14462 0 14518 800 0 FreeSans 224 90 0 0 la_data_out[8]
port 359 nsew signal tristate
flabel metal2 s 37094 0 37150 800 0 FreeSans 224 90 0 0 la_data_out[90]
port 360 nsew signal tristate
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 la_data_out[91]
port 361 nsew signal tristate
flabel metal2 s 37646 0 37702 800 0 FreeSans 224 90 0 0 la_data_out[92]
port 362 nsew signal tristate
flabel metal2 s 37922 0 37978 800 0 FreeSans 224 90 0 0 la_data_out[93]
port 363 nsew signal tristate
flabel metal2 s 38198 0 38254 800 0 FreeSans 224 90 0 0 la_data_out[94]
port 364 nsew signal tristate
flabel metal2 s 38474 0 38530 800 0 FreeSans 224 90 0 0 la_data_out[95]
port 365 nsew signal tristate
flabel metal2 s 38750 0 38806 800 0 FreeSans 224 90 0 0 la_data_out[96]
port 366 nsew signal tristate
flabel metal2 s 39026 0 39082 800 0 FreeSans 224 90 0 0 la_data_out[97]
port 367 nsew signal tristate
flabel metal2 s 39302 0 39358 800 0 FreeSans 224 90 0 0 la_data_out[98]
port 368 nsew signal tristate
flabel metal2 s 39578 0 39634 800 0 FreeSans 224 90 0 0 la_data_out[99]
port 369 nsew signal tristate
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 la_data_out[9]
port 370 nsew signal tristate
flabel metal2 s 12346 0 12402 800 0 FreeSans 224 90 0 0 la_oenb[0]
port 371 nsew signal input
flabel metal2 s 39946 0 40002 800 0 FreeSans 224 90 0 0 la_oenb[100]
port 372 nsew signal input
flabel metal2 s 40222 0 40278 800 0 FreeSans 224 90 0 0 la_oenb[101]
port 373 nsew signal input
flabel metal2 s 40498 0 40554 800 0 FreeSans 224 90 0 0 la_oenb[102]
port 374 nsew signal input
flabel metal2 s 40774 0 40830 800 0 FreeSans 224 90 0 0 la_oenb[103]
port 375 nsew signal input
flabel metal2 s 41050 0 41106 800 0 FreeSans 224 90 0 0 la_oenb[104]
port 376 nsew signal input
flabel metal2 s 41326 0 41382 800 0 FreeSans 224 90 0 0 la_oenb[105]
port 377 nsew signal input
flabel metal2 s 41602 0 41658 800 0 FreeSans 224 90 0 0 la_oenb[106]
port 378 nsew signal input
flabel metal2 s 41878 0 41934 800 0 FreeSans 224 90 0 0 la_oenb[107]
port 379 nsew signal input
flabel metal2 s 42154 0 42210 800 0 FreeSans 224 90 0 0 la_oenb[108]
port 380 nsew signal input
flabel metal2 s 42430 0 42486 800 0 FreeSans 224 90 0 0 la_oenb[109]
port 381 nsew signal input
flabel metal2 s 15106 0 15162 800 0 FreeSans 224 90 0 0 la_oenb[10]
port 382 nsew signal input
flabel metal2 s 42706 0 42762 800 0 FreeSans 224 90 0 0 la_oenb[110]
port 383 nsew signal input
flabel metal2 s 42982 0 43038 800 0 FreeSans 224 90 0 0 la_oenb[111]
port 384 nsew signal input
flabel metal2 s 43258 0 43314 800 0 FreeSans 224 90 0 0 la_oenb[112]
port 385 nsew signal input
flabel metal2 s 43534 0 43590 800 0 FreeSans 224 90 0 0 la_oenb[113]
port 386 nsew signal input
flabel metal2 s 43810 0 43866 800 0 FreeSans 224 90 0 0 la_oenb[114]
port 387 nsew signal input
flabel metal2 s 44086 0 44142 800 0 FreeSans 224 90 0 0 la_oenb[115]
port 388 nsew signal input
flabel metal2 s 44362 0 44418 800 0 FreeSans 224 90 0 0 la_oenb[116]
port 389 nsew signal input
flabel metal2 s 44638 0 44694 800 0 FreeSans 224 90 0 0 la_oenb[117]
port 390 nsew signal input
flabel metal2 s 44914 0 44970 800 0 FreeSans 224 90 0 0 la_oenb[118]
port 391 nsew signal input
flabel metal2 s 45190 0 45246 800 0 FreeSans 224 90 0 0 la_oenb[119]
port 392 nsew signal input
flabel metal2 s 15382 0 15438 800 0 FreeSans 224 90 0 0 la_oenb[11]
port 393 nsew signal input
flabel metal2 s 45466 0 45522 800 0 FreeSans 224 90 0 0 la_oenb[120]
port 394 nsew signal input
flabel metal2 s 45742 0 45798 800 0 FreeSans 224 90 0 0 la_oenb[121]
port 395 nsew signal input
flabel metal2 s 46018 0 46074 800 0 FreeSans 224 90 0 0 la_oenb[122]
port 396 nsew signal input
flabel metal2 s 46294 0 46350 800 0 FreeSans 224 90 0 0 la_oenb[123]
port 397 nsew signal input
flabel metal2 s 46570 0 46626 800 0 FreeSans 224 90 0 0 la_oenb[124]
port 398 nsew signal input
flabel metal2 s 46846 0 46902 800 0 FreeSans 224 90 0 0 la_oenb[125]
port 399 nsew signal input
flabel metal2 s 47122 0 47178 800 0 FreeSans 224 90 0 0 la_oenb[126]
port 400 nsew signal input
flabel metal2 s 47398 0 47454 800 0 FreeSans 224 90 0 0 la_oenb[127]
port 401 nsew signal input
flabel metal2 s 15658 0 15714 800 0 FreeSans 224 90 0 0 la_oenb[12]
port 402 nsew signal input
flabel metal2 s 15934 0 15990 800 0 FreeSans 224 90 0 0 la_oenb[13]
port 403 nsew signal input
flabel metal2 s 16210 0 16266 800 0 FreeSans 224 90 0 0 la_oenb[14]
port 404 nsew signal input
flabel metal2 s 16486 0 16542 800 0 FreeSans 224 90 0 0 la_oenb[15]
port 405 nsew signal input
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 la_oenb[16]
port 406 nsew signal input
flabel metal2 s 17038 0 17094 800 0 FreeSans 224 90 0 0 la_oenb[17]
port 407 nsew signal input
flabel metal2 s 17314 0 17370 800 0 FreeSans 224 90 0 0 la_oenb[18]
port 408 nsew signal input
flabel metal2 s 17590 0 17646 800 0 FreeSans 224 90 0 0 la_oenb[19]
port 409 nsew signal input
flabel metal2 s 12622 0 12678 800 0 FreeSans 224 90 0 0 la_oenb[1]
port 410 nsew signal input
flabel metal2 s 17866 0 17922 800 0 FreeSans 224 90 0 0 la_oenb[20]
port 411 nsew signal input
flabel metal2 s 18142 0 18198 800 0 FreeSans 224 90 0 0 la_oenb[21]
port 412 nsew signal input
flabel metal2 s 18418 0 18474 800 0 FreeSans 224 90 0 0 la_oenb[22]
port 413 nsew signal input
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 la_oenb[23]
port 414 nsew signal input
flabel metal2 s 18970 0 19026 800 0 FreeSans 224 90 0 0 la_oenb[24]
port 415 nsew signal input
flabel metal2 s 19246 0 19302 800 0 FreeSans 224 90 0 0 la_oenb[25]
port 416 nsew signal input
flabel metal2 s 19522 0 19578 800 0 FreeSans 224 90 0 0 la_oenb[26]
port 417 nsew signal input
flabel metal2 s 19798 0 19854 800 0 FreeSans 224 90 0 0 la_oenb[27]
port 418 nsew signal input
flabel metal2 s 20074 0 20130 800 0 FreeSans 224 90 0 0 la_oenb[28]
port 419 nsew signal input
flabel metal2 s 20350 0 20406 800 0 FreeSans 224 90 0 0 la_oenb[29]
port 420 nsew signal input
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 la_oenb[2]
port 421 nsew signal input
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 la_oenb[30]
port 422 nsew signal input
flabel metal2 s 20902 0 20958 800 0 FreeSans 224 90 0 0 la_oenb[31]
port 423 nsew signal input
flabel metal2 s 21178 0 21234 800 0 FreeSans 224 90 0 0 la_oenb[32]
port 424 nsew signal input
flabel metal2 s 21454 0 21510 800 0 FreeSans 224 90 0 0 la_oenb[33]
port 425 nsew signal input
flabel metal2 s 21730 0 21786 800 0 FreeSans 224 90 0 0 la_oenb[34]
port 426 nsew signal input
flabel metal2 s 22006 0 22062 800 0 FreeSans 224 90 0 0 la_oenb[35]
port 427 nsew signal input
flabel metal2 s 22282 0 22338 800 0 FreeSans 224 90 0 0 la_oenb[36]
port 428 nsew signal input
flabel metal2 s 22558 0 22614 800 0 FreeSans 224 90 0 0 la_oenb[37]
port 429 nsew signal input
flabel metal2 s 22834 0 22890 800 0 FreeSans 224 90 0 0 la_oenb[38]
port 430 nsew signal input
flabel metal2 s 23110 0 23166 800 0 FreeSans 224 90 0 0 la_oenb[39]
port 431 nsew signal input
flabel metal2 s 13174 0 13230 800 0 FreeSans 224 90 0 0 la_oenb[3]
port 432 nsew signal input
flabel metal2 s 23386 0 23442 800 0 FreeSans 224 90 0 0 la_oenb[40]
port 433 nsew signal input
flabel metal2 s 23662 0 23718 800 0 FreeSans 224 90 0 0 la_oenb[41]
port 434 nsew signal input
flabel metal2 s 23938 0 23994 800 0 FreeSans 224 90 0 0 la_oenb[42]
port 435 nsew signal input
flabel metal2 s 24214 0 24270 800 0 FreeSans 224 90 0 0 la_oenb[43]
port 436 nsew signal input
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 la_oenb[44]
port 437 nsew signal input
flabel metal2 s 24766 0 24822 800 0 FreeSans 224 90 0 0 la_oenb[45]
port 438 nsew signal input
flabel metal2 s 25042 0 25098 800 0 FreeSans 224 90 0 0 la_oenb[46]
port 439 nsew signal input
flabel metal2 s 25318 0 25374 800 0 FreeSans 224 90 0 0 la_oenb[47]
port 440 nsew signal input
flabel metal2 s 25594 0 25650 800 0 FreeSans 224 90 0 0 la_oenb[48]
port 441 nsew signal input
flabel metal2 s 25870 0 25926 800 0 FreeSans 224 90 0 0 la_oenb[49]
port 442 nsew signal input
flabel metal2 s 13450 0 13506 800 0 FreeSans 224 90 0 0 la_oenb[4]
port 443 nsew signal input
flabel metal2 s 26146 0 26202 800 0 FreeSans 224 90 0 0 la_oenb[50]
port 444 nsew signal input
flabel metal2 s 26422 0 26478 800 0 FreeSans 224 90 0 0 la_oenb[51]
port 445 nsew signal input
flabel metal2 s 26698 0 26754 800 0 FreeSans 224 90 0 0 la_oenb[52]
port 446 nsew signal input
flabel metal2 s 26974 0 27030 800 0 FreeSans 224 90 0 0 la_oenb[53]
port 447 nsew signal input
flabel metal2 s 27250 0 27306 800 0 FreeSans 224 90 0 0 la_oenb[54]
port 448 nsew signal input
flabel metal2 s 27526 0 27582 800 0 FreeSans 224 90 0 0 la_oenb[55]
port 449 nsew signal input
flabel metal2 s 27802 0 27858 800 0 FreeSans 224 90 0 0 la_oenb[56]
port 450 nsew signal input
flabel metal2 s 28078 0 28134 800 0 FreeSans 224 90 0 0 la_oenb[57]
port 451 nsew signal input
flabel metal2 s 28354 0 28410 800 0 FreeSans 224 90 0 0 la_oenb[58]
port 452 nsew signal input
flabel metal2 s 28630 0 28686 800 0 FreeSans 224 90 0 0 la_oenb[59]
port 453 nsew signal input
flabel metal2 s 13726 0 13782 800 0 FreeSans 224 90 0 0 la_oenb[5]
port 454 nsew signal input
flabel metal2 s 28906 0 28962 800 0 FreeSans 224 90 0 0 la_oenb[60]
port 455 nsew signal input
flabel metal2 s 29182 0 29238 800 0 FreeSans 224 90 0 0 la_oenb[61]
port 456 nsew signal input
flabel metal2 s 29458 0 29514 800 0 FreeSans 224 90 0 0 la_oenb[62]
port 457 nsew signal input
flabel metal2 s 29734 0 29790 800 0 FreeSans 224 90 0 0 la_oenb[63]
port 458 nsew signal input
flabel metal2 s 30010 0 30066 800 0 FreeSans 224 90 0 0 la_oenb[64]
port 459 nsew signal input
flabel metal2 s 30286 0 30342 800 0 FreeSans 224 90 0 0 la_oenb[65]
port 460 nsew signal input
flabel metal2 s 30562 0 30618 800 0 FreeSans 224 90 0 0 la_oenb[66]
port 461 nsew signal input
flabel metal2 s 30838 0 30894 800 0 FreeSans 224 90 0 0 la_oenb[67]
port 462 nsew signal input
flabel metal2 s 31114 0 31170 800 0 FreeSans 224 90 0 0 la_oenb[68]
port 463 nsew signal input
flabel metal2 s 31390 0 31446 800 0 FreeSans 224 90 0 0 la_oenb[69]
port 464 nsew signal input
flabel metal2 s 14002 0 14058 800 0 FreeSans 224 90 0 0 la_oenb[6]
port 465 nsew signal input
flabel metal2 s 31666 0 31722 800 0 FreeSans 224 90 0 0 la_oenb[70]
port 466 nsew signal input
flabel metal2 s 31942 0 31998 800 0 FreeSans 224 90 0 0 la_oenb[71]
port 467 nsew signal input
flabel metal2 s 32218 0 32274 800 0 FreeSans 224 90 0 0 la_oenb[72]
port 468 nsew signal input
flabel metal2 s 32494 0 32550 800 0 FreeSans 224 90 0 0 la_oenb[73]
port 469 nsew signal input
flabel metal2 s 32770 0 32826 800 0 FreeSans 224 90 0 0 la_oenb[74]
port 470 nsew signal input
flabel metal2 s 33046 0 33102 800 0 FreeSans 224 90 0 0 la_oenb[75]
port 471 nsew signal input
flabel metal2 s 33322 0 33378 800 0 FreeSans 224 90 0 0 la_oenb[76]
port 472 nsew signal input
flabel metal2 s 33598 0 33654 800 0 FreeSans 224 90 0 0 la_oenb[77]
port 473 nsew signal input
flabel metal2 s 33874 0 33930 800 0 FreeSans 224 90 0 0 la_oenb[78]
port 474 nsew signal input
flabel metal2 s 34150 0 34206 800 0 FreeSans 224 90 0 0 la_oenb[79]
port 475 nsew signal input
flabel metal2 s 14278 0 14334 800 0 FreeSans 224 90 0 0 la_oenb[7]
port 476 nsew signal input
flabel metal2 s 34426 0 34482 800 0 FreeSans 224 90 0 0 la_oenb[80]
port 477 nsew signal input
flabel metal2 s 34702 0 34758 800 0 FreeSans 224 90 0 0 la_oenb[81]
port 478 nsew signal input
flabel metal2 s 34978 0 35034 800 0 FreeSans 224 90 0 0 la_oenb[82]
port 479 nsew signal input
flabel metal2 s 35254 0 35310 800 0 FreeSans 224 90 0 0 la_oenb[83]
port 480 nsew signal input
flabel metal2 s 35530 0 35586 800 0 FreeSans 224 90 0 0 la_oenb[84]
port 481 nsew signal input
flabel metal2 s 35806 0 35862 800 0 FreeSans 224 90 0 0 la_oenb[85]
port 482 nsew signal input
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 la_oenb[86]
port 483 nsew signal input
flabel metal2 s 36358 0 36414 800 0 FreeSans 224 90 0 0 la_oenb[87]
port 484 nsew signal input
flabel metal2 s 36634 0 36690 800 0 FreeSans 224 90 0 0 la_oenb[88]
port 485 nsew signal input
flabel metal2 s 36910 0 36966 800 0 FreeSans 224 90 0 0 la_oenb[89]
port 486 nsew signal input
flabel metal2 s 14554 0 14610 800 0 FreeSans 224 90 0 0 la_oenb[8]
port 487 nsew signal input
flabel metal2 s 37186 0 37242 800 0 FreeSans 224 90 0 0 la_oenb[90]
port 488 nsew signal input
flabel metal2 s 37462 0 37518 800 0 FreeSans 224 90 0 0 la_oenb[91]
port 489 nsew signal input
flabel metal2 s 37738 0 37794 800 0 FreeSans 224 90 0 0 la_oenb[92]
port 490 nsew signal input
flabel metal2 s 38014 0 38070 800 0 FreeSans 224 90 0 0 la_oenb[93]
port 491 nsew signal input
flabel metal2 s 38290 0 38346 800 0 FreeSans 224 90 0 0 la_oenb[94]
port 492 nsew signal input
flabel metal2 s 38566 0 38622 800 0 FreeSans 224 90 0 0 la_oenb[95]
port 493 nsew signal input
flabel metal2 s 38842 0 38898 800 0 FreeSans 224 90 0 0 la_oenb[96]
port 494 nsew signal input
flabel metal2 s 39118 0 39174 800 0 FreeSans 224 90 0 0 la_oenb[97]
port 495 nsew signal input
flabel metal2 s 39394 0 39450 800 0 FreeSans 224 90 0 0 la_oenb[98]
port 496 nsew signal input
flabel metal2 s 39670 0 39726 800 0 FreeSans 224 90 0 0 la_oenb[99]
port 497 nsew signal input
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 la_oenb[9]
port 498 nsew signal input
flabel metal4 s 4208 2128 4528 47376 0 FreeSans 1920 90 0 0 vccd1
port 499 nsew power bidirectional
flabel metal4 s 34928 2128 35248 47376 0 FreeSans 1920 90 0 0 vccd1
port 499 nsew power bidirectional
flabel metal4 s 19568 2128 19888 47376 0 FreeSans 1920 90 0 0 vssd1
port 500 nsew ground bidirectional
flabel metal2 s 2410 0 2466 800 0 FreeSans 224 90 0 0 wb_clk_i
port 501 nsew signal input
flabel metal2 s 2502 0 2558 800 0 FreeSans 224 90 0 0 wb_rst_i
port 502 nsew signal input
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 wbs_ack_o
port 503 nsew signal tristate
flabel metal2 s 2962 0 3018 800 0 FreeSans 224 90 0 0 wbs_adr_i[0]
port 504 nsew signal input
flabel metal2 s 6090 0 6146 800 0 FreeSans 224 90 0 0 wbs_adr_i[10]
port 505 nsew signal input
flabel metal2 s 6366 0 6422 800 0 FreeSans 224 90 0 0 wbs_adr_i[11]
port 506 nsew signal input
flabel metal2 s 6642 0 6698 800 0 FreeSans 224 90 0 0 wbs_adr_i[12]
port 507 nsew signal input
flabel metal2 s 6918 0 6974 800 0 FreeSans 224 90 0 0 wbs_adr_i[13]
port 508 nsew signal input
flabel metal2 s 7194 0 7250 800 0 FreeSans 224 90 0 0 wbs_adr_i[14]
port 509 nsew signal input
flabel metal2 s 7470 0 7526 800 0 FreeSans 224 90 0 0 wbs_adr_i[15]
port 510 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 wbs_adr_i[16]
port 511 nsew signal input
flabel metal2 s 8022 0 8078 800 0 FreeSans 224 90 0 0 wbs_adr_i[17]
port 512 nsew signal input
flabel metal2 s 8298 0 8354 800 0 FreeSans 224 90 0 0 wbs_adr_i[18]
port 513 nsew signal input
flabel metal2 s 8574 0 8630 800 0 FreeSans 224 90 0 0 wbs_adr_i[19]
port 514 nsew signal input
flabel metal2 s 3330 0 3386 800 0 FreeSans 224 90 0 0 wbs_adr_i[1]
port 515 nsew signal input
flabel metal2 s 8850 0 8906 800 0 FreeSans 224 90 0 0 wbs_adr_i[20]
port 516 nsew signal input
flabel metal2 s 9126 0 9182 800 0 FreeSans 224 90 0 0 wbs_adr_i[21]
port 517 nsew signal input
flabel metal2 s 9402 0 9458 800 0 FreeSans 224 90 0 0 wbs_adr_i[22]
port 518 nsew signal input
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 wbs_adr_i[23]
port 519 nsew signal input
flabel metal2 s 9954 0 10010 800 0 FreeSans 224 90 0 0 wbs_adr_i[24]
port 520 nsew signal input
flabel metal2 s 10230 0 10286 800 0 FreeSans 224 90 0 0 wbs_adr_i[25]
port 521 nsew signal input
flabel metal2 s 10506 0 10562 800 0 FreeSans 224 90 0 0 wbs_adr_i[26]
port 522 nsew signal input
flabel metal2 s 10782 0 10838 800 0 FreeSans 224 90 0 0 wbs_adr_i[27]
port 523 nsew signal input
flabel metal2 s 11058 0 11114 800 0 FreeSans 224 90 0 0 wbs_adr_i[28]
port 524 nsew signal input
flabel metal2 s 11334 0 11390 800 0 FreeSans 224 90 0 0 wbs_adr_i[29]
port 525 nsew signal input
flabel metal2 s 3698 0 3754 800 0 FreeSans 224 90 0 0 wbs_adr_i[2]
port 526 nsew signal input
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 wbs_adr_i[30]
port 527 nsew signal input
flabel metal2 s 11886 0 11942 800 0 FreeSans 224 90 0 0 wbs_adr_i[31]
port 528 nsew signal input
flabel metal2 s 4066 0 4122 800 0 FreeSans 224 90 0 0 wbs_adr_i[3]
port 529 nsew signal input
flabel metal2 s 4434 0 4490 800 0 FreeSans 224 90 0 0 wbs_adr_i[4]
port 530 nsew signal input
flabel metal2 s 4710 0 4766 800 0 FreeSans 224 90 0 0 wbs_adr_i[5]
port 531 nsew signal input
flabel metal2 s 4986 0 5042 800 0 FreeSans 224 90 0 0 wbs_adr_i[6]
port 532 nsew signal input
flabel metal2 s 5262 0 5318 800 0 FreeSans 224 90 0 0 wbs_adr_i[7]
port 533 nsew signal input
flabel metal2 s 5538 0 5594 800 0 FreeSans 224 90 0 0 wbs_adr_i[8]
port 534 nsew signal input
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 wbs_adr_i[9]
port 535 nsew signal input
flabel metal2 s 2686 0 2742 800 0 FreeSans 224 90 0 0 wbs_cyc_i
port 536 nsew signal input
flabel metal2 s 3054 0 3110 800 0 FreeSans 224 90 0 0 wbs_dat_i[0]
port 537 nsew signal input
flabel metal2 s 6182 0 6238 800 0 FreeSans 224 90 0 0 wbs_dat_i[10]
port 538 nsew signal input
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 wbs_dat_i[11]
port 539 nsew signal input
flabel metal2 s 6734 0 6790 800 0 FreeSans 224 90 0 0 wbs_dat_i[12]
port 540 nsew signal input
flabel metal2 s 7010 0 7066 800 0 FreeSans 224 90 0 0 wbs_dat_i[13]
port 541 nsew signal input
flabel metal2 s 7286 0 7342 800 0 FreeSans 224 90 0 0 wbs_dat_i[14]
port 542 nsew signal input
flabel metal2 s 7562 0 7618 800 0 FreeSans 224 90 0 0 wbs_dat_i[15]
port 543 nsew signal input
flabel metal2 s 7838 0 7894 800 0 FreeSans 224 90 0 0 wbs_dat_i[16]
port 544 nsew signal input
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 wbs_dat_i[17]
port 545 nsew signal input
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 wbs_dat_i[18]
port 546 nsew signal input
flabel metal2 s 8666 0 8722 800 0 FreeSans 224 90 0 0 wbs_dat_i[19]
port 547 nsew signal input
flabel metal2 s 3422 0 3478 800 0 FreeSans 224 90 0 0 wbs_dat_i[1]
port 548 nsew signal input
flabel metal2 s 8942 0 8998 800 0 FreeSans 224 90 0 0 wbs_dat_i[20]
port 549 nsew signal input
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 wbs_dat_i[21]
port 550 nsew signal input
flabel metal2 s 9494 0 9550 800 0 FreeSans 224 90 0 0 wbs_dat_i[22]
port 551 nsew signal input
flabel metal2 s 9770 0 9826 800 0 FreeSans 224 90 0 0 wbs_dat_i[23]
port 552 nsew signal input
flabel metal2 s 10046 0 10102 800 0 FreeSans 224 90 0 0 wbs_dat_i[24]
port 553 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 wbs_dat_i[25]
port 554 nsew signal input
flabel metal2 s 10598 0 10654 800 0 FreeSans 224 90 0 0 wbs_dat_i[26]
port 555 nsew signal input
flabel metal2 s 10874 0 10930 800 0 FreeSans 224 90 0 0 wbs_dat_i[27]
port 556 nsew signal input
flabel metal2 s 11150 0 11206 800 0 FreeSans 224 90 0 0 wbs_dat_i[28]
port 557 nsew signal input
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 wbs_dat_i[29]
port 558 nsew signal input
flabel metal2 s 3790 0 3846 800 0 FreeSans 224 90 0 0 wbs_dat_i[2]
port 559 nsew signal input
flabel metal2 s 11702 0 11758 800 0 FreeSans 224 90 0 0 wbs_dat_i[30]
port 560 nsew signal input
flabel metal2 s 11978 0 12034 800 0 FreeSans 224 90 0 0 wbs_dat_i[31]
port 561 nsew signal input
flabel metal2 s 4158 0 4214 800 0 FreeSans 224 90 0 0 wbs_dat_i[3]
port 562 nsew signal input
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 wbs_dat_i[4]
port 563 nsew signal input
flabel metal2 s 4802 0 4858 800 0 FreeSans 224 90 0 0 wbs_dat_i[5]
port 564 nsew signal input
flabel metal2 s 5078 0 5134 800 0 FreeSans 224 90 0 0 wbs_dat_i[6]
port 565 nsew signal input
flabel metal2 s 5354 0 5410 800 0 FreeSans 224 90 0 0 wbs_dat_i[7]
port 566 nsew signal input
flabel metal2 s 5630 0 5686 800 0 FreeSans 224 90 0 0 wbs_dat_i[8]
port 567 nsew signal input
flabel metal2 s 5906 0 5962 800 0 FreeSans 224 90 0 0 wbs_dat_i[9]
port 568 nsew signal input
flabel metal2 s 3146 0 3202 800 0 FreeSans 224 90 0 0 wbs_dat_o[0]
port 569 nsew signal tristate
flabel metal2 s 6274 0 6330 800 0 FreeSans 224 90 0 0 wbs_dat_o[10]
port 570 nsew signal tristate
flabel metal2 s 6550 0 6606 800 0 FreeSans 224 90 0 0 wbs_dat_o[11]
port 571 nsew signal tristate
flabel metal2 s 6826 0 6882 800 0 FreeSans 224 90 0 0 wbs_dat_o[12]
port 572 nsew signal tristate
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 wbs_dat_o[13]
port 573 nsew signal tristate
flabel metal2 s 7378 0 7434 800 0 FreeSans 224 90 0 0 wbs_dat_o[14]
port 574 nsew signal tristate
flabel metal2 s 7654 0 7710 800 0 FreeSans 224 90 0 0 wbs_dat_o[15]
port 575 nsew signal tristate
flabel metal2 s 7930 0 7986 800 0 FreeSans 224 90 0 0 wbs_dat_o[16]
port 576 nsew signal tristate
flabel metal2 s 8206 0 8262 800 0 FreeSans 224 90 0 0 wbs_dat_o[17]
port 577 nsew signal tristate
flabel metal2 s 8482 0 8538 800 0 FreeSans 224 90 0 0 wbs_dat_o[18]
port 578 nsew signal tristate
flabel metal2 s 8758 0 8814 800 0 FreeSans 224 90 0 0 wbs_dat_o[19]
port 579 nsew signal tristate
flabel metal2 s 3514 0 3570 800 0 FreeSans 224 90 0 0 wbs_dat_o[1]
port 580 nsew signal tristate
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 wbs_dat_o[20]
port 581 nsew signal tristate
flabel metal2 s 9310 0 9366 800 0 FreeSans 224 90 0 0 wbs_dat_o[21]
port 582 nsew signal tristate
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 wbs_dat_o[22]
port 583 nsew signal tristate
flabel metal2 s 9862 0 9918 800 0 FreeSans 224 90 0 0 wbs_dat_o[23]
port 584 nsew signal tristate
flabel metal2 s 10138 0 10194 800 0 FreeSans 224 90 0 0 wbs_dat_o[24]
port 585 nsew signal tristate
flabel metal2 s 10414 0 10470 800 0 FreeSans 224 90 0 0 wbs_dat_o[25]
port 586 nsew signal tristate
flabel metal2 s 10690 0 10746 800 0 FreeSans 224 90 0 0 wbs_dat_o[26]
port 587 nsew signal tristate
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 wbs_dat_o[27]
port 588 nsew signal tristate
flabel metal2 s 11242 0 11298 800 0 FreeSans 224 90 0 0 wbs_dat_o[28]
port 589 nsew signal tristate
flabel metal2 s 11518 0 11574 800 0 FreeSans 224 90 0 0 wbs_dat_o[29]
port 590 nsew signal tristate
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 wbs_dat_o[2]
port 591 nsew signal tristate
flabel metal2 s 11794 0 11850 800 0 FreeSans 224 90 0 0 wbs_dat_o[30]
port 592 nsew signal tristate
flabel metal2 s 12070 0 12126 800 0 FreeSans 224 90 0 0 wbs_dat_o[31]
port 593 nsew signal tristate
flabel metal2 s 4250 0 4306 800 0 FreeSans 224 90 0 0 wbs_dat_o[3]
port 594 nsew signal tristate
flabel metal2 s 4618 0 4674 800 0 FreeSans 224 90 0 0 wbs_dat_o[4]
port 595 nsew signal tristate
flabel metal2 s 4894 0 4950 800 0 FreeSans 224 90 0 0 wbs_dat_o[5]
port 596 nsew signal tristate
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 wbs_dat_o[6]
port 597 nsew signal tristate
flabel metal2 s 5446 0 5502 800 0 FreeSans 224 90 0 0 wbs_dat_o[7]
port 598 nsew signal tristate
flabel metal2 s 5722 0 5778 800 0 FreeSans 224 90 0 0 wbs_dat_o[8]
port 599 nsew signal tristate
flabel metal2 s 5998 0 6054 800 0 FreeSans 224 90 0 0 wbs_dat_o[9]
port 600 nsew signal tristate
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 wbs_sel_i[0]
port 601 nsew signal input
flabel metal2 s 3606 0 3662 800 0 FreeSans 224 90 0 0 wbs_sel_i[1]
port 602 nsew signal input
flabel metal2 s 3974 0 4030 800 0 FreeSans 224 90 0 0 wbs_sel_i[2]
port 603 nsew signal input
flabel metal2 s 4342 0 4398 800 0 FreeSans 224 90 0 0 wbs_sel_i[3]
port 604 nsew signal input
flabel metal2 s 2778 0 2834 800 0 FreeSans 224 90 0 0 wbs_stb_i
port 605 nsew signal input
flabel metal2 s 2870 0 2926 800 0 FreeSans 224 90 0 0 wbs_we_i
port 606 nsew signal input
rlabel metal1 24978 47328 24978 47328 0 vccd1
rlabel metal1 24978 46784 24978 46784 0 vssd1
rlabel metal1 27646 44914 27646 44914 0 _000_
rlabel metal1 28520 45934 28520 45934 0 _001_
rlabel metal1 25484 46546 25484 46546 0 _002_
rlabel metal2 23690 46104 23690 46104 0 _003_
rlabel metal1 29762 43962 29762 43962 0 _004_
rlabel metal2 25530 44132 25530 44132 0 _005_
rlabel metal1 24748 42874 24748 42874 0 _006_
rlabel metal2 28198 44744 28198 44744 0 _007_
rlabel metal1 28658 44778 28658 44778 0 _008_
rlabel metal2 28106 44098 28106 44098 0 _009_
rlabel metal2 26634 44098 26634 44098 0 _010_
rlabel metal1 26404 44370 26404 44370 0 _011_
rlabel metal1 25484 44302 25484 44302 0 _012_
rlabel metal2 24702 45900 24702 45900 0 _013_
rlabel metal2 24610 44132 24610 44132 0 _014_
rlabel metal1 23046 45356 23046 45356 0 _015_
rlabel metal1 23920 45798 23920 45798 0 _016_
rlabel metal1 20746 45968 20746 45968 0 _017_
rlabel metal1 22494 45900 22494 45900 0 _018_
rlabel metal2 22862 46308 22862 46308 0 _019_
rlabel metal1 39054 45526 39054 45526 0 _020_
rlabel metal2 37950 46070 37950 46070 0 _021_
rlabel metal2 31786 45934 31786 45934 0 _022_
rlabel metal2 32522 46342 32522 46342 0 _023_
rlabel metal2 37582 44710 37582 44710 0 _024_
rlabel metal1 33449 44846 33449 44846 0 _025_
rlabel metal2 32614 44710 32614 44710 0 _026_
rlabel metal1 36294 44506 36294 44506 0 _027_
rlabel metal1 36064 44438 36064 44438 0 _028_
rlabel metal2 35466 44098 35466 44098 0 _029_
rlabel metal2 34638 44812 34638 44812 0 _030_
rlabel metal2 35374 44132 35374 44132 0 _031_
rlabel metal1 33074 45934 33074 45934 0 _032_
rlabel metal1 32430 45492 32430 45492 0 _033_
rlabel metal2 32338 45254 32338 45254 0 _034_
rlabel metal2 32338 46036 32338 46036 0 _035_
rlabel metal2 32890 46393 32890 46393 0 _036_
rlabel metal1 31004 47022 31004 47022 0 _037_
rlabel metal1 31004 46954 31004 46954 0 _038_
rlabel metal1 22862 46410 22862 46410 0 _039_
rlabel metal1 27830 45968 27830 45968 0 _040_
rlabel metal1 25944 46682 25944 46682 0 _041_
rlabel metal1 25392 45526 25392 45526 0 _042_
rlabel metal1 20102 46614 20102 46614 0 _043_
rlabel metal1 33580 46478 33580 46478 0 _044_
rlabel metal1 34960 46682 34960 46682 0 _045_
rlabel viali 33903 47022 33903 47022 0 _046_
rlabel metal2 19918 47192 19918 47192 0 _047_
rlabel metal1 18906 46138 18906 46138 0 _048_
rlabel metal1 19366 45458 19366 45458 0 _049_
rlabel metal2 27278 43588 27278 43588 0 _050_
rlabel metal2 27554 45118 27554 45118 0 _051_
rlabel metal2 28566 46784 28566 46784 0 _052_
rlabel metal2 27370 46308 27370 46308 0 _053_
rlabel metal1 21572 45934 21572 45934 0 _054_
rlabel metal1 34914 43962 34914 43962 0 _055_
rlabel metal1 35926 44370 35926 44370 0 _056_
rlabel metal2 36110 46444 36110 46444 0 _057_
rlabel metal1 36156 46138 36156 46138 0 _058_
rlabel metal2 37582 46053 37582 46053 0 _059_
rlabel metal2 20470 46376 20470 46376 0 _060_
rlabel metal1 20700 46070 20700 46070 0 _061_
rlabel metal1 26312 45594 26312 45594 0 _062_
rlabel metal1 27186 45390 27186 45390 0 _063_
rlabel metal1 25668 44370 25668 44370 0 _064_
rlabel metal1 26165 45390 26165 45390 0 _065_
rlabel metal2 25438 44982 25438 44982 0 _066_
rlabel metal1 22310 45492 22310 45492 0 _067_
rlabel metal2 34086 46240 34086 46240 0 _068_
rlabel metal2 34546 44370 34546 44370 0 _069_
rlabel metal1 33856 44914 33856 44914 0 _070_
rlabel metal2 33718 44676 33718 44676 0 _071_
rlabel metal2 33626 45662 33626 45662 0 _072_
rlabel metal2 33442 45118 33442 45118 0 _073_
rlabel metal2 20838 44540 20838 44540 0 _074_
rlabel metal2 22034 45050 22034 45050 0 _075_
rlabel metal2 23966 44132 23966 44132 0 _076_
rlabel metal2 23414 44540 23414 44540 0 _077_
rlabel metal1 21735 47022 21735 47022 0 _078_
rlabel metal1 22540 47090 22540 47090 0 _079_
rlabel via1 24426 46546 24426 46546 0 _080_
rlabel metal2 24334 46393 24334 46393 0 _081_
rlabel metal2 22770 45866 22770 45866 0 _082_
rlabel metal2 31878 45662 31878 45662 0 _083_
rlabel metal2 32890 45594 32890 45594 0 _084_
rlabel metal2 31326 45696 31326 45696 0 _085_
rlabel metal1 35834 46580 35834 46580 0 _086_
rlabel metal1 32062 46036 32062 46036 0 _087_
rlabel metal2 30866 46682 30866 46682 0 _088_
rlabel metal2 20562 6562 20562 6562 0 _089_
rlabel metal1 30728 2414 30728 2414 0 _090_
rlabel metal1 20148 3026 20148 3026 0 _091_
rlabel metal2 21114 5984 21114 5984 0 _092_
rlabel metal2 20378 4760 20378 4760 0 _093_
rlabel metal1 20056 3434 20056 3434 0 _094_
rlabel metal1 19596 3094 19596 3094 0 _095_
rlabel metal1 20930 2312 20930 2312 0 _096_
rlabel metal2 21758 5032 21758 5032 0 _097_
rlabel metal1 21206 4148 21206 4148 0 _098_
rlabel metal1 22586 2312 22586 2312 0 _099_
rlabel metal2 22586 5848 22586 5848 0 _100_
rlabel metal2 23138 5678 23138 5678 0 _101_
rlabel metal2 23230 5576 23230 5576 0 _102_
rlabel metal2 23046 3230 23046 3230 0 _103_
rlabel metal1 24794 2312 24794 2312 0 _104_
rlabel metal1 24242 3128 24242 3128 0 _105_
rlabel metal1 24150 2618 24150 2618 0 _106_
rlabel metal1 24150 6358 24150 6358 0 _107_
rlabel metal1 24104 4250 24104 4250 0 _108_
rlabel via1 25350 3434 25350 3434 0 _109_
rlabel metal1 25392 3094 25392 3094 0 _110_
rlabel metal1 25668 4250 25668 4250 0 _111_
rlabel metal1 26174 5576 26174 5576 0 _112_
rlabel metal2 25070 6120 25070 6120 0 _113_
rlabel metal1 27370 3128 27370 3128 0 _114_
rlabel metal1 28428 2346 28428 2346 0 _115_
rlabel metal1 27324 3706 27324 3706 0 _116_
rlabel metal2 27370 5406 27370 5406 0 _117_
rlabel metal2 28566 5406 28566 5406 0 _118_
rlabel metal1 30406 2618 30406 2618 0 _119_
rlabel metal2 28934 3230 28934 3230 0 _120_
rlabel metal2 29072 4522 29072 4522 0 _121_
rlabel metal1 29394 4182 29394 4182 0 _122_
rlabel metal1 30820 3094 30820 3094 0 _123_
rlabel metal2 29026 46291 29026 46291 0 _124_
rlabel metal2 20286 5168 20286 5168 0 _125_
rlabel metal1 20056 3570 20056 3570 0 _126_
rlabel metal1 19274 2958 19274 2958 0 _127_
rlabel metal1 19228 2482 19228 2482 0 _128_
rlabel metal1 21666 4692 21666 4692 0 _129_
rlabel metal1 20884 4046 20884 4046 0 _130_
rlabel metal1 22402 2482 22402 2482 0 _131_
rlabel metal1 22218 5746 22218 5746 0 _132_
rlabel metal1 22264 5134 22264 5134 0 _133_
rlabel metal1 21390 3910 21390 3910 0 _134_
rlabel metal2 18906 2244 18906 2244 0 _135_
rlabel metal1 23966 2346 23966 2346 0 _136_
rlabel metal2 24150 3366 24150 3366 0 _137_
rlabel metal1 24242 4012 24242 4012 0 _138_
rlabel metal2 24058 6052 24058 6052 0 _139_
rlabel metal1 23000 5066 23000 5066 0 _140_
rlabel metal1 25254 3604 25254 3604 0 _141_
rlabel metal1 27922 2822 27922 2822 0 _142_
rlabel metal1 25346 4658 25346 4658 0 _143_
rlabel metal1 26358 5202 26358 5202 0 _144_
rlabel metal1 25852 5202 25852 5202 0 _145_
rlabel metal1 26818 2618 26818 2618 0 _146_
rlabel metal1 28106 2482 28106 2482 0 _147_
rlabel metal2 28934 3876 28934 3876 0 _148_
rlabel metal2 27370 4964 27370 4964 0 _149_
rlabel metal1 27554 3978 27554 3978 0 _150_
rlabel metal1 29578 2890 29578 2890 0 _151_
rlabel metal1 30038 3162 30038 3162 0 _152_
rlabel metal1 29072 4658 29072 4658 0 _153_
rlabel metal2 29762 3876 29762 3876 0 _154_
rlabel metal1 32016 2618 32016 2618 0 _155_
rlabel metal1 31142 44302 31142 44302 0 _156_
rlabel metal2 3397 49300 3397 49300 0 io_active
rlabel metal1 24196 45526 24196 45526 0 io_in[18]
rlabel metal1 29716 47022 29716 47022 0 io_in[19]
rlabel metal1 26772 45934 26772 45934 0 io_in[20]
rlabel metal1 25530 46036 25530 46036 0 io_in[21]
rlabel metal1 32154 45900 32154 45900 0 io_in[22]
rlabel metal1 30314 47056 30314 47056 0 io_in[23]
rlabel metal1 29302 44438 29302 44438 0 io_in[24]
rlabel metal1 29164 41242 29164 41242 0 io_in[25]
rlabel metal1 33396 46954 33396 46954 0 io_in[26]
rlabel metal2 37766 47260 37766 47260 0 io_in[27]
rlabel metal2 35466 48127 35466 48127 0 io_in[28]
rlabel metal1 38732 46546 38732 46546 0 io_in[29]
rlabel metal2 40250 45764 40250 45764 0 io_in[30]
rlabel metal1 42320 45254 42320 45254 0 io_in[31]
rlabel metal1 40204 45050 40204 45050 0 io_in[32]
rlabel metal2 39698 42908 39698 42908 0 io_in[33]
rlabel metal2 41906 47984 41906 47984 0 io_in[34]
rlabel metal2 43010 47593 43010 47593 0 io_in[35]
rlabel metal2 43838 47719 43838 47719 0 io_in[36]
rlabel metal1 43010 45050 43010 45050 0 io_in[37]
rlabel metal2 4738 48256 4738 48256 0 io_oeb[0]
rlabel metal2 15686 48263 15686 48263 0 io_oeb[10]
rlabel metal1 16606 47226 16606 47226 0 io_oeb[11]
rlabel metal1 17710 46546 17710 46546 0 io_oeb[12]
rlabel metal1 18676 46070 18676 46070 0 io_oeb[13]
rlabel metal1 18906 47090 18906 47090 0 io_oeb[14]
rlabel metal1 18814 47158 18814 47158 0 io_oeb[15]
rlabel metal1 19780 46478 19780 46478 0 io_oeb[16]
rlabel metal2 18906 47328 18906 47328 0 io_oeb[17]
rlabel metal1 23644 44234 23644 44234 0 io_oeb[18]
rlabel metal1 25254 46138 25254 46138 0 io_oeb[19]
rlabel metal1 5612 47226 5612 47226 0 io_oeb[1]
rlabel metal1 28888 47158 28888 47158 0 io_oeb[20]
rlabel metal1 28060 43214 28060 43214 0 io_oeb[21]
rlabel metal1 33166 46342 33166 46342 0 io_oeb[22]
rlabel metal1 30498 43962 30498 43962 0 io_oeb[23]
rlabel metal2 31418 46631 31418 46631 0 io_oeb[24]
rlabel metal2 34178 45832 34178 45832 0 io_oeb[25]
rlabel metal2 39146 46801 39146 46801 0 io_oeb[26]
rlabel metal1 38778 46342 38778 46342 0 io_oeb[27]
rlabel metal2 40710 46937 40710 46937 0 io_oeb[28]
rlabel metal1 38548 46070 38548 46070 0 io_oeb[29]
rlabel metal2 6946 47916 6946 47916 0 io_oeb[2]
rlabel metal1 38134 45050 38134 45050 0 io_oeb[30]
rlabel metal1 40020 46478 40020 46478 0 io_oeb[31]
rlabel metal2 40066 47916 40066 47916 0 io_oeb[32]
rlabel metal2 41354 47719 41354 47719 0 io_oeb[33]
rlabel metal1 42458 46546 42458 46546 0 io_oeb[34]
rlabel metal1 43654 47226 43654 47226 0 io_oeb[35]
rlabel metal2 44482 47916 44482 47916 0 io_oeb[36]
rlabel metal2 45862 48263 45862 48263 0 io_oeb[37]
rlabel metal2 7774 48263 7774 48263 0 io_oeb[3]
rlabel metal2 9154 48256 9154 48256 0 io_oeb[4]
rlabel metal2 10258 48256 10258 48256 0 io_oeb[5]
rlabel metal2 11178 48263 11178 48263 0 io_oeb[6]
rlabel metal2 12466 48256 12466 48256 0 io_oeb[7]
rlabel metal2 13570 48256 13570 48256 0 io_oeb[8]
rlabel metal2 14674 48256 14674 48256 0 io_oeb[9]
rlabel metal2 5106 47865 5106 47865 0 io_out[0]
rlabel metal1 17020 46682 17020 46682 0 io_out[10]
rlabel metal1 18722 45832 18722 45832 0 io_out[11]
rlabel metal1 20930 45390 20930 45390 0 io_out[12]
rlabel metal2 20286 47090 20286 47090 0 io_out[13]
rlabel metal1 20056 47158 20056 47158 0 io_out[14]
rlabel metal1 21206 46410 21206 46410 0 io_out[15]
rlabel metal2 22586 47311 22586 47311 0 io_out[16]
rlabel metal2 23874 48188 23874 48188 0 io_out[17]
rlabel metal1 25254 43282 25254 43282 0 io_out[18]
rlabel metal1 26726 47226 26726 47226 0 io_out[19]
rlabel metal2 6026 48263 6026 48263 0 io_out[1]
rlabel metal2 27186 47168 27186 47168 0 io_out[20]
rlabel metal1 30176 45050 30176 45050 0 io_out[21]
rlabel metal2 29210 46631 29210 46631 0 io_out[22]
rlabel metal1 32706 46478 32706 46478 0 io_out[23]
rlabel metal2 31602 46284 31602 46284 0 io_out[24]
rlabel metal1 35604 47226 35604 47226 0 io_out[25]
rlabel metal2 33810 46284 33810 46284 0 io_out[26]
rlabel metal1 40112 47022 40112 47022 0 io_out[27]
rlabel metal1 39652 46410 39652 46410 0 io_out[28]
rlabel metal1 39238 47158 39238 47158 0 io_out[29]
rlabel metal2 7130 48263 7130 48263 0 io_out[2]
rlabel metal1 39606 45526 39606 45526 0 io_out[30]
rlabel metal1 40020 46138 40020 46138 0 io_out[31]
rlabel metal2 40710 48263 40710 48263 0 io_out[32]
rlabel metal1 41768 46138 41768 46138 0 io_out[33]
rlabel metal1 43056 47226 43056 47226 0 io_out[34]
rlabel metal2 43746 47916 43746 47916 0 io_out[35]
rlabel metal1 45034 47226 45034 47226 0 io_out[36]
rlabel metal1 46230 47226 46230 47226 0 io_out[37]
rlabel metal2 8418 48256 8418 48256 0 io_out[3]
rlabel metal2 9522 47933 9522 47933 0 io_out[4]
rlabel metal2 10626 47593 10626 47593 0 io_out[5]
rlabel metal2 11730 47610 11730 47610 0 io_out[6]
rlabel metal2 12834 47950 12834 47950 0 io_out[7]
rlabel metal1 17296 45594 17296 45594 0 io_out[8]
rlabel metal2 15042 47797 15042 47797 0 io_out[9]
rlabel metal2 12282 1588 12282 1588 0 la_data_out[0]
rlabel metal2 39882 1588 39882 1588 0 la_data_out[100]
rlabel metal2 40158 1792 40158 1792 0 la_data_out[101]
rlabel metal2 40434 2132 40434 2132 0 la_data_out[102]
rlabel metal2 40710 1860 40710 1860 0 la_data_out[103]
rlabel metal2 40986 2132 40986 2132 0 la_data_out[104]
rlabel metal2 41262 1622 41262 1622 0 la_data_out[105]
rlabel metal2 41538 2132 41538 2132 0 la_data_out[106]
rlabel metal2 41814 1588 41814 1588 0 la_data_out[107]
rlabel metal2 42090 1792 42090 1792 0 la_data_out[108]
rlabel metal2 42366 1656 42366 1656 0 la_data_out[109]
rlabel metal2 15042 2336 15042 2336 0 la_data_out[10]
rlabel metal2 42642 1860 42642 1860 0 la_data_out[110]
rlabel metal2 42918 2132 42918 2132 0 la_data_out[111]
rlabel metal2 43194 2132 43194 2132 0 la_data_out[112]
rlabel metal2 43470 1792 43470 1792 0 la_data_out[113]
rlabel metal2 43746 1622 43746 1622 0 la_data_out[114]
rlabel metal2 44022 1792 44022 1792 0 la_data_out[115]
rlabel metal2 44298 1554 44298 1554 0 la_data_out[116]
rlabel metal2 44574 1860 44574 1860 0 la_data_out[117]
rlabel metal2 44850 2132 44850 2132 0 la_data_out[118]
rlabel metal2 45126 1656 45126 1656 0 la_data_out[119]
rlabel metal2 15318 1792 15318 1792 0 la_data_out[11]
rlabel metal2 45402 1792 45402 1792 0 la_data_out[120]
rlabel metal2 45678 2132 45678 2132 0 la_data_out[121]
rlabel metal2 45954 1792 45954 1792 0 la_data_out[122]
rlabel metal2 46230 1588 46230 1588 0 la_data_out[123]
rlabel metal2 46506 2132 46506 2132 0 la_data_out[124]
rlabel metal2 46782 2132 46782 2132 0 la_data_out[125]
rlabel metal2 47058 1792 47058 1792 0 la_data_out[126]
rlabel metal2 47334 2132 47334 2132 0 la_data_out[127]
rlabel metal2 15594 1588 15594 1588 0 la_data_out[12]
rlabel metal2 15870 2166 15870 2166 0 la_data_out[13]
rlabel metal2 16146 2336 16146 2336 0 la_data_out[14]
rlabel metal2 16422 2132 16422 2132 0 la_data_out[15]
rlabel metal2 16698 1894 16698 1894 0 la_data_out[16]
rlabel metal2 16974 2676 16974 2676 0 la_data_out[17]
rlabel metal2 17250 2200 17250 2200 0 la_data_out[18]
rlabel metal2 17526 1826 17526 1826 0 la_data_out[19]
rlabel metal2 12558 2132 12558 2132 0 la_data_out[1]
rlabel metal2 17802 1792 17802 1792 0 la_data_out[20]
rlabel metal2 18078 2336 18078 2336 0 la_data_out[21]
rlabel metal2 18354 1656 18354 1656 0 la_data_out[22]
rlabel metal2 18630 2166 18630 2166 0 la_data_out[23]
rlabel metal2 18906 1163 18906 1163 0 la_data_out[24]
rlabel metal2 19182 2370 19182 2370 0 la_data_out[25]
rlabel metal2 19458 2880 19458 2880 0 la_data_out[26]
rlabel metal2 19734 1418 19734 1418 0 la_data_out[27]
rlabel metal2 20010 1350 20010 1350 0 la_data_out[28]
rlabel metal2 20286 2200 20286 2200 0 la_data_out[29]
rlabel metal2 12834 1622 12834 1622 0 la_data_out[2]
rlabel metal2 20562 1792 20562 1792 0 la_data_out[30]
rlabel metal2 20838 2234 20838 2234 0 la_data_out[31]
rlabel metal2 21114 2642 21114 2642 0 la_data_out[32]
rlabel metal2 21390 2166 21390 2166 0 la_data_out[33]
rlabel metal2 21666 1860 21666 1860 0 la_data_out[34]
rlabel metal2 21942 1554 21942 1554 0 la_data_out[35]
rlabel metal2 22218 2744 22218 2744 0 la_data_out[36]
rlabel metal2 22494 2404 22494 2404 0 la_data_out[37]
rlabel metal2 22770 1622 22770 1622 0 la_data_out[38]
rlabel metal2 23046 1761 23046 1761 0 la_data_out[39]
rlabel metal2 13110 2132 13110 2132 0 la_data_out[3]
rlabel metal2 23322 1761 23322 1761 0 la_data_out[40]
rlabel metal2 23598 2710 23598 2710 0 la_data_out[41]
rlabel metal1 23736 2958 23736 2958 0 la_data_out[42]
rlabel metal2 24150 1622 24150 1622 0 la_data_out[43]
rlabel metal2 24426 1860 24426 1860 0 la_data_out[44]
rlabel metal2 24702 2404 24702 2404 0 la_data_out[45]
rlabel metal2 24978 3458 24978 3458 0 la_data_out[46]
rlabel metal1 25208 5134 25208 5134 0 la_data_out[47]
rlabel metal2 25530 2166 25530 2166 0 la_data_out[48]
rlabel metal2 25806 1860 25806 1860 0 la_data_out[49]
rlabel metal2 13386 1826 13386 1826 0 la_data_out[4]
rlabel metal2 26082 2710 26082 2710 0 la_data_out[50]
rlabel metal2 26312 5780 26312 5780 0 la_data_out[51]
rlabel metal1 26588 6222 26588 6222 0 la_data_out[52]
rlabel metal1 27232 2890 27232 2890 0 la_data_out[53]
rlabel metal2 27186 1554 27186 1554 0 la_data_out[54]
rlabel metal2 27462 2404 27462 2404 0 la_data_out[55]
rlabel metal2 27738 1639 27738 1639 0 la_data_out[56]
rlabel metal1 28612 3638 28612 3638 0 la_data_out[57]
rlabel metal1 28198 3570 28198 3570 0 la_data_out[58]
rlabel metal2 28566 1860 28566 1860 0 la_data_out[59]
rlabel metal2 13662 2132 13662 2132 0 la_data_out[5]
rlabel metal2 28842 2710 28842 2710 0 la_data_out[60]
rlabel metal1 29118 3944 29118 3944 0 la_data_out[61]
rlabel metal1 29486 2958 29486 2958 0 la_data_out[62]
rlabel metal2 29900 12420 29900 12420 0 la_data_out[63]
rlabel metal1 30130 3910 30130 3910 0 la_data_out[64]
rlabel metal1 30636 3570 30636 3570 0 la_data_out[65]
rlabel metal2 30498 1554 30498 1554 0 la_data_out[66]
rlabel metal2 30820 2890 30820 2890 0 la_data_out[67]
rlabel metal2 31050 1299 31050 1299 0 la_data_out[68]
rlabel metal2 31326 1622 31326 1622 0 la_data_out[69]
rlabel metal2 13938 1792 13938 1792 0 la_data_out[6]
rlabel metal2 31602 1826 31602 1826 0 la_data_out[70]
rlabel metal2 31878 2132 31878 2132 0 la_data_out[71]
rlabel metal2 32154 1860 32154 1860 0 la_data_out[72]
rlabel metal2 32430 2132 32430 2132 0 la_data_out[73]
rlabel metal2 32706 1894 32706 1894 0 la_data_out[74]
rlabel metal2 32982 2200 32982 2200 0 la_data_out[75]
rlabel metal2 33258 1656 33258 1656 0 la_data_out[76]
rlabel metal2 33534 1826 33534 1826 0 la_data_out[77]
rlabel metal2 33810 1588 33810 1588 0 la_data_out[78]
rlabel metal2 34086 1860 34086 1860 0 la_data_out[79]
rlabel metal2 14214 1656 14214 1656 0 la_data_out[7]
rlabel metal2 34362 2132 34362 2132 0 la_data_out[80]
rlabel metal2 34638 1622 34638 1622 0 la_data_out[81]
rlabel metal2 34914 1299 34914 1299 0 la_data_out[82]
rlabel metal2 35190 1095 35190 1095 0 la_data_out[83]
rlabel metal2 35466 1656 35466 1656 0 la_data_out[84]
rlabel metal2 35742 2132 35742 2132 0 la_data_out[85]
rlabel metal2 36018 1792 36018 1792 0 la_data_out[86]
rlabel metal2 36294 2132 36294 2132 0 la_data_out[87]
rlabel metal2 36570 1588 36570 1588 0 la_data_out[88]
rlabel metal2 36846 2200 36846 2200 0 la_data_out[89]
rlabel metal2 14490 1826 14490 1826 0 la_data_out[8]
rlabel metal2 37122 1860 37122 1860 0 la_data_out[90]
rlabel metal2 37398 1622 37398 1622 0 la_data_out[91]
rlabel metal2 37674 2132 37674 2132 0 la_data_out[92]
rlabel metal2 37950 1826 37950 1826 0 la_data_out[93]
rlabel metal2 38226 2132 38226 2132 0 la_data_out[94]
rlabel metal2 38502 1656 38502 1656 0 la_data_out[95]
rlabel metal2 38778 1860 38778 1860 0 la_data_out[96]
rlabel metal2 39054 1792 39054 1792 0 la_data_out[97]
rlabel metal2 39330 1622 39330 1622 0 la_data_out[98]
rlabel metal2 39606 2132 39606 2132 0 la_data_out[99]
rlabel metal2 14766 1622 14766 1622 0 la_data_out[9]
rlabel metal2 2622 1588 2622 1588 0 wbs_ack_o
rlabel metal2 3174 1792 3174 1792 0 wbs_dat_o[0]
rlabel metal2 6302 1826 6302 1826 0 wbs_dat_o[10]
rlabel metal2 6578 1792 6578 1792 0 wbs_dat_o[11]
rlabel metal2 6854 2132 6854 2132 0 wbs_dat_o[12]
rlabel metal2 7130 1656 7130 1656 0 wbs_dat_o[13]
rlabel metal1 6463 2414 6463 2414 0 wbs_dat_o[14]
rlabel metal2 7682 2132 7682 2132 0 wbs_dat_o[15]
rlabel metal2 7958 1860 7958 1860 0 wbs_dat_o[16]
rlabel metal2 8234 1622 8234 1622 0 wbs_dat_o[17]
rlabel metal2 8510 2132 8510 2132 0 wbs_dat_o[18]
rlabel metal2 8786 1826 8786 1826 0 wbs_dat_o[19]
rlabel metal2 3542 1622 3542 1622 0 wbs_dat_o[1]
rlabel metal2 9062 1792 9062 1792 0 wbs_dat_o[20]
rlabel metal2 9338 2132 9338 2132 0 wbs_dat_o[21]
rlabel metal2 9614 1656 9614 1656 0 wbs_dat_o[22]
rlabel metal2 9890 1860 9890 1860 0 wbs_dat_o[23]
rlabel metal2 10166 2132 10166 2132 0 wbs_dat_o[24]
rlabel metal2 10442 1622 10442 1622 0 wbs_dat_o[25]
rlabel metal2 10718 1792 10718 1792 0 wbs_dat_o[26]
rlabel metal2 10994 2132 10994 2132 0 wbs_dat_o[27]
rlabel metal2 11270 1826 11270 1826 0 wbs_dat_o[28]
rlabel metal2 11546 1656 11546 1656 0 wbs_dat_o[29]
rlabel metal2 3910 1792 3910 1792 0 wbs_dat_o[2]
rlabel metal2 11822 2132 11822 2132 0 wbs_dat_o[30]
rlabel metal2 12098 1792 12098 1792 0 wbs_dat_o[31]
rlabel metal2 4278 1656 4278 1656 0 wbs_dat_o[3]
rlabel metal2 4646 1588 4646 1588 0 wbs_dat_o[4]
rlabel metal2 4922 1826 4922 1826 0 wbs_dat_o[5]
rlabel metal2 5198 2132 5198 2132 0 wbs_dat_o[6]
rlabel metal2 5474 1860 5474 1860 0 wbs_dat_o[7]
rlabel metal2 5750 1588 5750 1588 0 wbs_dat_o[8]
rlabel metal2 6026 2132 6026 2132 0 wbs_dat_o[9]
<< properties >>
string FIXED_BBOX 0 0 50000 50000
<< end >>
