magic
tech sky130A
magscale 1 2
timestamp 1666199351
<< nwell >>
rect -126 0 4006 338
rect 4048 0 8180 338
rect 8222 0 11354 338
rect 11396 0 14528 338
rect 14570 0 18702 338
rect 18744 0 22876 338
<< mvpmos >>
rect -60 119 3940 219
rect 4114 119 8114 219
rect 8288 119 11288 219
rect 11462 119 14462 219
rect 14636 119 18636 219
rect 18810 119 22810 219
<< mvpdiff >>
rect -60 264 3940 272
rect -60 230 18 264
rect 52 230 86 264
rect 120 230 154 264
rect 188 230 222 264
rect 256 230 290 264
rect 324 230 358 264
rect 392 230 426 264
rect 460 230 494 264
rect 528 230 562 264
rect 596 230 630 264
rect 664 230 698 264
rect 732 230 766 264
rect 800 230 834 264
rect 868 230 902 264
rect 936 230 970 264
rect 1004 230 1038 264
rect 1072 230 1106 264
rect 1140 230 1174 264
rect 1208 230 1242 264
rect 1276 230 1310 264
rect 1344 230 1378 264
rect 1412 230 1446 264
rect 1480 230 1514 264
rect 1548 230 1582 264
rect 1616 230 1650 264
rect 1684 230 1718 264
rect 1752 230 1786 264
rect 1820 230 1854 264
rect 1888 230 1922 264
rect 1956 230 1990 264
rect 2024 230 2058 264
rect 2092 230 2126 264
rect 2160 230 2194 264
rect 2228 230 2262 264
rect 2296 230 2330 264
rect 2364 230 2398 264
rect 2432 230 2466 264
rect 2500 230 2534 264
rect 2568 230 2602 264
rect 2636 230 2670 264
rect 2704 230 2738 264
rect 2772 230 2806 264
rect 2840 230 2874 264
rect 2908 230 2942 264
rect 2976 230 3010 264
rect 3044 230 3078 264
rect 3112 230 3146 264
rect 3180 230 3214 264
rect 3248 230 3282 264
rect 3316 230 3350 264
rect 3384 230 3418 264
rect 3452 230 3486 264
rect 3520 230 3554 264
rect 3588 230 3622 264
rect 3656 230 3690 264
rect 3724 230 3758 264
rect 3792 230 3826 264
rect 3860 230 3894 264
rect 3928 230 3940 264
rect -60 219 3940 230
rect 4114 264 8114 272
rect 4114 230 4192 264
rect 4226 230 4260 264
rect 4294 230 4328 264
rect 4362 230 4396 264
rect 4430 230 4464 264
rect 4498 230 4532 264
rect 4566 230 4600 264
rect 4634 230 4668 264
rect 4702 230 4736 264
rect 4770 230 4804 264
rect 4838 230 4872 264
rect 4906 230 4940 264
rect 4974 230 5008 264
rect 5042 230 5076 264
rect 5110 230 5144 264
rect 5178 230 5212 264
rect 5246 230 5280 264
rect 5314 230 5348 264
rect 5382 230 5416 264
rect 5450 230 5484 264
rect 5518 230 5552 264
rect 5586 230 5620 264
rect 5654 230 5688 264
rect 5722 230 5756 264
rect 5790 230 5824 264
rect 5858 230 5892 264
rect 5926 230 5960 264
rect 5994 230 6028 264
rect 6062 230 6096 264
rect 6130 230 6164 264
rect 6198 230 6232 264
rect 6266 230 6300 264
rect 6334 230 6368 264
rect 6402 230 6436 264
rect 6470 230 6504 264
rect 6538 230 6572 264
rect 6606 230 6640 264
rect 6674 230 6708 264
rect 6742 230 6776 264
rect 6810 230 6844 264
rect 6878 230 6912 264
rect 6946 230 6980 264
rect 7014 230 7048 264
rect 7082 230 7116 264
rect 7150 230 7184 264
rect 7218 230 7252 264
rect 7286 230 7320 264
rect 7354 230 7388 264
rect 7422 230 7456 264
rect 7490 230 7524 264
rect 7558 230 7592 264
rect 7626 230 7660 264
rect 7694 230 7728 264
rect 7762 230 7796 264
rect 7830 230 7864 264
rect 7898 230 7932 264
rect 7966 230 8000 264
rect 8034 230 8068 264
rect 8102 230 8114 264
rect 4114 219 8114 230
rect 8288 264 11288 272
rect 8288 230 8318 264
rect 8352 230 8386 264
rect 8420 230 8454 264
rect 8488 230 8522 264
rect 8556 230 8590 264
rect 8624 230 8658 264
rect 8692 230 8726 264
rect 8760 230 8794 264
rect 8828 230 8862 264
rect 8896 230 8930 264
rect 8964 230 8998 264
rect 9032 230 9066 264
rect 9100 230 9134 264
rect 9168 230 9202 264
rect 9236 230 9270 264
rect 9304 230 9338 264
rect 9372 230 9406 264
rect 9440 230 9474 264
rect 9508 230 9542 264
rect 9576 230 9610 264
rect 9644 230 9678 264
rect 9712 230 9746 264
rect 9780 230 9814 264
rect 9848 230 9882 264
rect 9916 230 9950 264
rect 9984 230 10018 264
rect 10052 230 10086 264
rect 10120 230 10154 264
rect 10188 230 10222 264
rect 10256 230 10290 264
rect 10324 230 10358 264
rect 10392 230 10426 264
rect 10460 230 10494 264
rect 10528 230 10562 264
rect 10596 230 10630 264
rect 10664 230 10698 264
rect 10732 230 10766 264
rect 10800 230 10834 264
rect 10868 230 10902 264
rect 10936 230 10970 264
rect 11004 230 11038 264
rect 11072 230 11106 264
rect 11140 230 11174 264
rect 11208 230 11242 264
rect 11276 230 11288 264
rect 8288 219 11288 230
rect 11462 264 14462 272
rect 11462 230 11474 264
rect 11508 230 11542 264
rect 11576 230 11610 264
rect 11644 230 11678 264
rect 11712 230 11746 264
rect 11780 230 11814 264
rect 11848 230 11882 264
rect 11916 230 11950 264
rect 11984 230 12018 264
rect 12052 230 12086 264
rect 12120 230 12154 264
rect 12188 230 12222 264
rect 12256 230 12290 264
rect 12324 230 12358 264
rect 12392 230 12426 264
rect 12460 230 12494 264
rect 12528 230 12562 264
rect 12596 230 12630 264
rect 12664 230 12698 264
rect 12732 230 12766 264
rect 12800 230 12834 264
rect 12868 230 12902 264
rect 12936 230 12970 264
rect 13004 230 13038 264
rect 13072 230 13106 264
rect 13140 230 13174 264
rect 13208 230 13242 264
rect 13276 230 13310 264
rect 13344 230 13378 264
rect 13412 230 13446 264
rect 13480 230 13514 264
rect 13548 230 13582 264
rect 13616 230 13650 264
rect 13684 230 13718 264
rect 13752 230 13786 264
rect 13820 230 13854 264
rect 13888 230 13922 264
rect 13956 230 13990 264
rect 14024 230 14058 264
rect 14092 230 14126 264
rect 14160 230 14194 264
rect 14228 230 14262 264
rect 14296 230 14330 264
rect 14364 230 14398 264
rect 14432 230 14462 264
rect 11462 219 14462 230
rect 14636 264 18636 272
rect 14636 230 14648 264
rect 14682 230 14716 264
rect 14750 230 14784 264
rect 14818 230 14852 264
rect 14886 230 14920 264
rect 14954 230 14988 264
rect 15022 230 15056 264
rect 15090 230 15124 264
rect 15158 230 15192 264
rect 15226 230 15260 264
rect 15294 230 15328 264
rect 15362 230 15396 264
rect 15430 230 15464 264
rect 15498 230 15532 264
rect 15566 230 15600 264
rect 15634 230 15668 264
rect 15702 230 15736 264
rect 15770 230 15804 264
rect 15838 230 15872 264
rect 15906 230 15940 264
rect 15974 230 16008 264
rect 16042 230 16076 264
rect 16110 230 16144 264
rect 16178 230 16212 264
rect 16246 230 16280 264
rect 16314 230 16348 264
rect 16382 230 16416 264
rect 16450 230 16484 264
rect 16518 230 16552 264
rect 16586 230 16620 264
rect 16654 230 16688 264
rect 16722 230 16756 264
rect 16790 230 16824 264
rect 16858 230 16892 264
rect 16926 230 16960 264
rect 16994 230 17028 264
rect 17062 230 17096 264
rect 17130 230 17164 264
rect 17198 230 17232 264
rect 17266 230 17300 264
rect 17334 230 17368 264
rect 17402 230 17436 264
rect 17470 230 17504 264
rect 17538 230 17572 264
rect 17606 230 17640 264
rect 17674 230 17708 264
rect 17742 230 17776 264
rect 17810 230 17844 264
rect 17878 230 17912 264
rect 17946 230 17980 264
rect 18014 230 18048 264
rect 18082 230 18116 264
rect 18150 230 18184 264
rect 18218 230 18252 264
rect 18286 230 18320 264
rect 18354 230 18388 264
rect 18422 230 18456 264
rect 18490 230 18524 264
rect 18558 230 18636 264
rect 14636 219 18636 230
rect 18810 264 22810 272
rect 18810 230 18822 264
rect 18856 230 18890 264
rect 18924 230 18958 264
rect 18992 230 19026 264
rect 19060 230 19094 264
rect 19128 230 19162 264
rect 19196 230 19230 264
rect 19264 230 19298 264
rect 19332 230 19366 264
rect 19400 230 19434 264
rect 19468 230 19502 264
rect 19536 230 19570 264
rect 19604 230 19638 264
rect 19672 230 19706 264
rect 19740 230 19774 264
rect 19808 230 19842 264
rect 19876 230 19910 264
rect 19944 230 19978 264
rect 20012 230 20046 264
rect 20080 230 20114 264
rect 20148 230 20182 264
rect 20216 230 20250 264
rect 20284 230 20318 264
rect 20352 230 20386 264
rect 20420 230 20454 264
rect 20488 230 20522 264
rect 20556 230 20590 264
rect 20624 230 20658 264
rect 20692 230 20726 264
rect 20760 230 20794 264
rect 20828 230 20862 264
rect 20896 230 20930 264
rect 20964 230 20998 264
rect 21032 230 21066 264
rect 21100 230 21134 264
rect 21168 230 21202 264
rect 21236 230 21270 264
rect 21304 230 21338 264
rect 21372 230 21406 264
rect 21440 230 21474 264
rect 21508 230 21542 264
rect 21576 230 21610 264
rect 21644 230 21678 264
rect 21712 230 21746 264
rect 21780 230 21814 264
rect 21848 230 21882 264
rect 21916 230 21950 264
rect 21984 230 22018 264
rect 22052 230 22086 264
rect 22120 230 22154 264
rect 22188 230 22222 264
rect 22256 230 22290 264
rect 22324 230 22358 264
rect 22392 230 22426 264
rect 22460 230 22494 264
rect 22528 230 22562 264
rect 22596 230 22630 264
rect 22664 230 22698 264
rect 22732 230 22810 264
rect 18810 219 22810 230
rect -60 108 3940 119
rect -60 74 18 108
rect 52 74 86 108
rect 120 74 154 108
rect 188 74 222 108
rect 256 74 290 108
rect 324 74 358 108
rect 392 74 426 108
rect 460 74 494 108
rect 528 74 562 108
rect 596 74 630 108
rect 664 74 698 108
rect 732 74 766 108
rect 800 74 834 108
rect 868 74 902 108
rect 936 74 970 108
rect 1004 74 1038 108
rect 1072 74 1106 108
rect 1140 74 1174 108
rect 1208 74 1242 108
rect 1276 74 1310 108
rect 1344 74 1378 108
rect 1412 74 1446 108
rect 1480 74 1514 108
rect 1548 74 1582 108
rect 1616 74 1650 108
rect 1684 74 1718 108
rect 1752 74 1786 108
rect 1820 74 1854 108
rect 1888 74 1922 108
rect 1956 74 1990 108
rect 2024 74 2058 108
rect 2092 74 2126 108
rect 2160 74 2194 108
rect 2228 74 2262 108
rect 2296 74 2330 108
rect 2364 74 2398 108
rect 2432 74 2466 108
rect 2500 74 2534 108
rect 2568 74 2602 108
rect 2636 74 2670 108
rect 2704 74 2738 108
rect 2772 74 2806 108
rect 2840 74 2874 108
rect 2908 74 2942 108
rect 2976 74 3010 108
rect 3044 74 3078 108
rect 3112 74 3146 108
rect 3180 74 3214 108
rect 3248 74 3282 108
rect 3316 74 3350 108
rect 3384 74 3418 108
rect 3452 74 3486 108
rect 3520 74 3554 108
rect 3588 74 3622 108
rect 3656 74 3690 108
rect 3724 74 3758 108
rect 3792 74 3826 108
rect 3860 74 3894 108
rect 3928 74 3940 108
rect -60 66 3940 74
rect 4114 108 8114 119
rect 4114 74 4192 108
rect 4226 74 4260 108
rect 4294 74 4328 108
rect 4362 74 4396 108
rect 4430 74 4464 108
rect 4498 74 4532 108
rect 4566 74 4600 108
rect 4634 74 4668 108
rect 4702 74 4736 108
rect 4770 74 4804 108
rect 4838 74 4872 108
rect 4906 74 4940 108
rect 4974 74 5008 108
rect 5042 74 5076 108
rect 5110 74 5144 108
rect 5178 74 5212 108
rect 5246 74 5280 108
rect 5314 74 5348 108
rect 5382 74 5416 108
rect 5450 74 5484 108
rect 5518 74 5552 108
rect 5586 74 5620 108
rect 5654 74 5688 108
rect 5722 74 5756 108
rect 5790 74 5824 108
rect 5858 74 5892 108
rect 5926 74 5960 108
rect 5994 74 6028 108
rect 6062 74 6096 108
rect 6130 74 6164 108
rect 6198 74 6232 108
rect 6266 74 6300 108
rect 6334 74 6368 108
rect 6402 74 6436 108
rect 6470 74 6504 108
rect 6538 74 6572 108
rect 6606 74 6640 108
rect 6674 74 6708 108
rect 6742 74 6776 108
rect 6810 74 6844 108
rect 6878 74 6912 108
rect 6946 74 6980 108
rect 7014 74 7048 108
rect 7082 74 7116 108
rect 7150 74 7184 108
rect 7218 74 7252 108
rect 7286 74 7320 108
rect 7354 74 7388 108
rect 7422 74 7456 108
rect 7490 74 7524 108
rect 7558 74 7592 108
rect 7626 74 7660 108
rect 7694 74 7728 108
rect 7762 74 7796 108
rect 7830 74 7864 108
rect 7898 74 7932 108
rect 7966 74 8000 108
rect 8034 74 8068 108
rect 8102 74 8114 108
rect 4114 66 8114 74
rect 8288 108 11288 119
rect 8288 74 8318 108
rect 8352 74 8386 108
rect 8420 74 8454 108
rect 8488 74 8522 108
rect 8556 74 8590 108
rect 8624 74 8658 108
rect 8692 74 8726 108
rect 8760 74 8794 108
rect 8828 74 8862 108
rect 8896 74 8930 108
rect 8964 74 8998 108
rect 9032 74 9066 108
rect 9100 74 9134 108
rect 9168 74 9202 108
rect 9236 74 9270 108
rect 9304 74 9338 108
rect 9372 74 9406 108
rect 9440 74 9474 108
rect 9508 74 9542 108
rect 9576 74 9610 108
rect 9644 74 9678 108
rect 9712 74 9746 108
rect 9780 74 9814 108
rect 9848 74 9882 108
rect 9916 74 9950 108
rect 9984 74 10018 108
rect 10052 74 10086 108
rect 10120 74 10154 108
rect 10188 74 10222 108
rect 10256 74 10290 108
rect 10324 74 10358 108
rect 10392 74 10426 108
rect 10460 74 10494 108
rect 10528 74 10562 108
rect 10596 74 10630 108
rect 10664 74 10698 108
rect 10732 74 10766 108
rect 10800 74 10834 108
rect 10868 74 10902 108
rect 10936 74 10970 108
rect 11004 74 11038 108
rect 11072 74 11106 108
rect 11140 74 11174 108
rect 11208 74 11242 108
rect 11276 74 11288 108
rect 8288 66 11288 74
rect 11462 108 14462 119
rect 11462 74 11474 108
rect 11508 74 11542 108
rect 11576 74 11610 108
rect 11644 74 11678 108
rect 11712 74 11746 108
rect 11780 74 11814 108
rect 11848 74 11882 108
rect 11916 74 11950 108
rect 11984 74 12018 108
rect 12052 74 12086 108
rect 12120 74 12154 108
rect 12188 74 12222 108
rect 12256 74 12290 108
rect 12324 74 12358 108
rect 12392 74 12426 108
rect 12460 74 12494 108
rect 12528 74 12562 108
rect 12596 74 12630 108
rect 12664 74 12698 108
rect 12732 74 12766 108
rect 12800 74 12834 108
rect 12868 74 12902 108
rect 12936 74 12970 108
rect 13004 74 13038 108
rect 13072 74 13106 108
rect 13140 74 13174 108
rect 13208 74 13242 108
rect 13276 74 13310 108
rect 13344 74 13378 108
rect 13412 74 13446 108
rect 13480 74 13514 108
rect 13548 74 13582 108
rect 13616 74 13650 108
rect 13684 74 13718 108
rect 13752 74 13786 108
rect 13820 74 13854 108
rect 13888 74 13922 108
rect 13956 74 13990 108
rect 14024 74 14058 108
rect 14092 74 14126 108
rect 14160 74 14194 108
rect 14228 74 14262 108
rect 14296 74 14330 108
rect 14364 74 14398 108
rect 14432 74 14462 108
rect 11462 66 14462 74
rect 14636 108 18636 119
rect 14636 74 14648 108
rect 14682 74 14716 108
rect 14750 74 14784 108
rect 14818 74 14852 108
rect 14886 74 14920 108
rect 14954 74 14988 108
rect 15022 74 15056 108
rect 15090 74 15124 108
rect 15158 74 15192 108
rect 15226 74 15260 108
rect 15294 74 15328 108
rect 15362 74 15396 108
rect 15430 74 15464 108
rect 15498 74 15532 108
rect 15566 74 15600 108
rect 15634 74 15668 108
rect 15702 74 15736 108
rect 15770 74 15804 108
rect 15838 74 15872 108
rect 15906 74 15940 108
rect 15974 74 16008 108
rect 16042 74 16076 108
rect 16110 74 16144 108
rect 16178 74 16212 108
rect 16246 74 16280 108
rect 16314 74 16348 108
rect 16382 74 16416 108
rect 16450 74 16484 108
rect 16518 74 16552 108
rect 16586 74 16620 108
rect 16654 74 16688 108
rect 16722 74 16756 108
rect 16790 74 16824 108
rect 16858 74 16892 108
rect 16926 74 16960 108
rect 16994 74 17028 108
rect 17062 74 17096 108
rect 17130 74 17164 108
rect 17198 74 17232 108
rect 17266 74 17300 108
rect 17334 74 17368 108
rect 17402 74 17436 108
rect 17470 74 17504 108
rect 17538 74 17572 108
rect 17606 74 17640 108
rect 17674 74 17708 108
rect 17742 74 17776 108
rect 17810 74 17844 108
rect 17878 74 17912 108
rect 17946 74 17980 108
rect 18014 74 18048 108
rect 18082 74 18116 108
rect 18150 74 18184 108
rect 18218 74 18252 108
rect 18286 74 18320 108
rect 18354 74 18388 108
rect 18422 74 18456 108
rect 18490 74 18524 108
rect 18558 74 18636 108
rect 14636 66 18636 74
rect 18810 108 22810 119
rect 18810 74 18822 108
rect 18856 74 18890 108
rect 18924 74 18958 108
rect 18992 74 19026 108
rect 19060 74 19094 108
rect 19128 74 19162 108
rect 19196 74 19230 108
rect 19264 74 19298 108
rect 19332 74 19366 108
rect 19400 74 19434 108
rect 19468 74 19502 108
rect 19536 74 19570 108
rect 19604 74 19638 108
rect 19672 74 19706 108
rect 19740 74 19774 108
rect 19808 74 19842 108
rect 19876 74 19910 108
rect 19944 74 19978 108
rect 20012 74 20046 108
rect 20080 74 20114 108
rect 20148 74 20182 108
rect 20216 74 20250 108
rect 20284 74 20318 108
rect 20352 74 20386 108
rect 20420 74 20454 108
rect 20488 74 20522 108
rect 20556 74 20590 108
rect 20624 74 20658 108
rect 20692 74 20726 108
rect 20760 74 20794 108
rect 20828 74 20862 108
rect 20896 74 20930 108
rect 20964 74 20998 108
rect 21032 74 21066 108
rect 21100 74 21134 108
rect 21168 74 21202 108
rect 21236 74 21270 108
rect 21304 74 21338 108
rect 21372 74 21406 108
rect 21440 74 21474 108
rect 21508 74 21542 108
rect 21576 74 21610 108
rect 21644 74 21678 108
rect 21712 74 21746 108
rect 21780 74 21814 108
rect 21848 74 21882 108
rect 21916 74 21950 108
rect 21984 74 22018 108
rect 22052 74 22086 108
rect 22120 74 22154 108
rect 22188 74 22222 108
rect 22256 74 22290 108
rect 22324 74 22358 108
rect 22392 74 22426 108
rect 22460 74 22494 108
rect 22528 74 22562 108
rect 22596 74 22630 108
rect 22664 74 22698 108
rect 22732 74 22810 108
rect 18810 66 22810 74
<< mvpdiffc >>
rect 18 230 52 264
rect 86 230 120 264
rect 154 230 188 264
rect 222 230 256 264
rect 290 230 324 264
rect 358 230 392 264
rect 426 230 460 264
rect 494 230 528 264
rect 562 230 596 264
rect 630 230 664 264
rect 698 230 732 264
rect 766 230 800 264
rect 834 230 868 264
rect 902 230 936 264
rect 970 230 1004 264
rect 1038 230 1072 264
rect 1106 230 1140 264
rect 1174 230 1208 264
rect 1242 230 1276 264
rect 1310 230 1344 264
rect 1378 230 1412 264
rect 1446 230 1480 264
rect 1514 230 1548 264
rect 1582 230 1616 264
rect 1650 230 1684 264
rect 1718 230 1752 264
rect 1786 230 1820 264
rect 1854 230 1888 264
rect 1922 230 1956 264
rect 1990 230 2024 264
rect 2058 230 2092 264
rect 2126 230 2160 264
rect 2194 230 2228 264
rect 2262 230 2296 264
rect 2330 230 2364 264
rect 2398 230 2432 264
rect 2466 230 2500 264
rect 2534 230 2568 264
rect 2602 230 2636 264
rect 2670 230 2704 264
rect 2738 230 2772 264
rect 2806 230 2840 264
rect 2874 230 2908 264
rect 2942 230 2976 264
rect 3010 230 3044 264
rect 3078 230 3112 264
rect 3146 230 3180 264
rect 3214 230 3248 264
rect 3282 230 3316 264
rect 3350 230 3384 264
rect 3418 230 3452 264
rect 3486 230 3520 264
rect 3554 230 3588 264
rect 3622 230 3656 264
rect 3690 230 3724 264
rect 3758 230 3792 264
rect 3826 230 3860 264
rect 3894 230 3928 264
rect 4192 230 4226 264
rect 4260 230 4294 264
rect 4328 230 4362 264
rect 4396 230 4430 264
rect 4464 230 4498 264
rect 4532 230 4566 264
rect 4600 230 4634 264
rect 4668 230 4702 264
rect 4736 230 4770 264
rect 4804 230 4838 264
rect 4872 230 4906 264
rect 4940 230 4974 264
rect 5008 230 5042 264
rect 5076 230 5110 264
rect 5144 230 5178 264
rect 5212 230 5246 264
rect 5280 230 5314 264
rect 5348 230 5382 264
rect 5416 230 5450 264
rect 5484 230 5518 264
rect 5552 230 5586 264
rect 5620 230 5654 264
rect 5688 230 5722 264
rect 5756 230 5790 264
rect 5824 230 5858 264
rect 5892 230 5926 264
rect 5960 230 5994 264
rect 6028 230 6062 264
rect 6096 230 6130 264
rect 6164 230 6198 264
rect 6232 230 6266 264
rect 6300 230 6334 264
rect 6368 230 6402 264
rect 6436 230 6470 264
rect 6504 230 6538 264
rect 6572 230 6606 264
rect 6640 230 6674 264
rect 6708 230 6742 264
rect 6776 230 6810 264
rect 6844 230 6878 264
rect 6912 230 6946 264
rect 6980 230 7014 264
rect 7048 230 7082 264
rect 7116 230 7150 264
rect 7184 230 7218 264
rect 7252 230 7286 264
rect 7320 230 7354 264
rect 7388 230 7422 264
rect 7456 230 7490 264
rect 7524 230 7558 264
rect 7592 230 7626 264
rect 7660 230 7694 264
rect 7728 230 7762 264
rect 7796 230 7830 264
rect 7864 230 7898 264
rect 7932 230 7966 264
rect 8000 230 8034 264
rect 8068 230 8102 264
rect 8318 230 8352 264
rect 8386 230 8420 264
rect 8454 230 8488 264
rect 8522 230 8556 264
rect 8590 230 8624 264
rect 8658 230 8692 264
rect 8726 230 8760 264
rect 8794 230 8828 264
rect 8862 230 8896 264
rect 8930 230 8964 264
rect 8998 230 9032 264
rect 9066 230 9100 264
rect 9134 230 9168 264
rect 9202 230 9236 264
rect 9270 230 9304 264
rect 9338 230 9372 264
rect 9406 230 9440 264
rect 9474 230 9508 264
rect 9542 230 9576 264
rect 9610 230 9644 264
rect 9678 230 9712 264
rect 9746 230 9780 264
rect 9814 230 9848 264
rect 9882 230 9916 264
rect 9950 230 9984 264
rect 10018 230 10052 264
rect 10086 230 10120 264
rect 10154 230 10188 264
rect 10222 230 10256 264
rect 10290 230 10324 264
rect 10358 230 10392 264
rect 10426 230 10460 264
rect 10494 230 10528 264
rect 10562 230 10596 264
rect 10630 230 10664 264
rect 10698 230 10732 264
rect 10766 230 10800 264
rect 10834 230 10868 264
rect 10902 230 10936 264
rect 10970 230 11004 264
rect 11038 230 11072 264
rect 11106 230 11140 264
rect 11174 230 11208 264
rect 11242 230 11276 264
rect 11474 230 11508 264
rect 11542 230 11576 264
rect 11610 230 11644 264
rect 11678 230 11712 264
rect 11746 230 11780 264
rect 11814 230 11848 264
rect 11882 230 11916 264
rect 11950 230 11984 264
rect 12018 230 12052 264
rect 12086 230 12120 264
rect 12154 230 12188 264
rect 12222 230 12256 264
rect 12290 230 12324 264
rect 12358 230 12392 264
rect 12426 230 12460 264
rect 12494 230 12528 264
rect 12562 230 12596 264
rect 12630 230 12664 264
rect 12698 230 12732 264
rect 12766 230 12800 264
rect 12834 230 12868 264
rect 12902 230 12936 264
rect 12970 230 13004 264
rect 13038 230 13072 264
rect 13106 230 13140 264
rect 13174 230 13208 264
rect 13242 230 13276 264
rect 13310 230 13344 264
rect 13378 230 13412 264
rect 13446 230 13480 264
rect 13514 230 13548 264
rect 13582 230 13616 264
rect 13650 230 13684 264
rect 13718 230 13752 264
rect 13786 230 13820 264
rect 13854 230 13888 264
rect 13922 230 13956 264
rect 13990 230 14024 264
rect 14058 230 14092 264
rect 14126 230 14160 264
rect 14194 230 14228 264
rect 14262 230 14296 264
rect 14330 230 14364 264
rect 14398 230 14432 264
rect 14648 230 14682 264
rect 14716 230 14750 264
rect 14784 230 14818 264
rect 14852 230 14886 264
rect 14920 230 14954 264
rect 14988 230 15022 264
rect 15056 230 15090 264
rect 15124 230 15158 264
rect 15192 230 15226 264
rect 15260 230 15294 264
rect 15328 230 15362 264
rect 15396 230 15430 264
rect 15464 230 15498 264
rect 15532 230 15566 264
rect 15600 230 15634 264
rect 15668 230 15702 264
rect 15736 230 15770 264
rect 15804 230 15838 264
rect 15872 230 15906 264
rect 15940 230 15974 264
rect 16008 230 16042 264
rect 16076 230 16110 264
rect 16144 230 16178 264
rect 16212 230 16246 264
rect 16280 230 16314 264
rect 16348 230 16382 264
rect 16416 230 16450 264
rect 16484 230 16518 264
rect 16552 230 16586 264
rect 16620 230 16654 264
rect 16688 230 16722 264
rect 16756 230 16790 264
rect 16824 230 16858 264
rect 16892 230 16926 264
rect 16960 230 16994 264
rect 17028 230 17062 264
rect 17096 230 17130 264
rect 17164 230 17198 264
rect 17232 230 17266 264
rect 17300 230 17334 264
rect 17368 230 17402 264
rect 17436 230 17470 264
rect 17504 230 17538 264
rect 17572 230 17606 264
rect 17640 230 17674 264
rect 17708 230 17742 264
rect 17776 230 17810 264
rect 17844 230 17878 264
rect 17912 230 17946 264
rect 17980 230 18014 264
rect 18048 230 18082 264
rect 18116 230 18150 264
rect 18184 230 18218 264
rect 18252 230 18286 264
rect 18320 230 18354 264
rect 18388 230 18422 264
rect 18456 230 18490 264
rect 18524 230 18558 264
rect 18822 230 18856 264
rect 18890 230 18924 264
rect 18958 230 18992 264
rect 19026 230 19060 264
rect 19094 230 19128 264
rect 19162 230 19196 264
rect 19230 230 19264 264
rect 19298 230 19332 264
rect 19366 230 19400 264
rect 19434 230 19468 264
rect 19502 230 19536 264
rect 19570 230 19604 264
rect 19638 230 19672 264
rect 19706 230 19740 264
rect 19774 230 19808 264
rect 19842 230 19876 264
rect 19910 230 19944 264
rect 19978 230 20012 264
rect 20046 230 20080 264
rect 20114 230 20148 264
rect 20182 230 20216 264
rect 20250 230 20284 264
rect 20318 230 20352 264
rect 20386 230 20420 264
rect 20454 230 20488 264
rect 20522 230 20556 264
rect 20590 230 20624 264
rect 20658 230 20692 264
rect 20726 230 20760 264
rect 20794 230 20828 264
rect 20862 230 20896 264
rect 20930 230 20964 264
rect 20998 230 21032 264
rect 21066 230 21100 264
rect 21134 230 21168 264
rect 21202 230 21236 264
rect 21270 230 21304 264
rect 21338 230 21372 264
rect 21406 230 21440 264
rect 21474 230 21508 264
rect 21542 230 21576 264
rect 21610 230 21644 264
rect 21678 230 21712 264
rect 21746 230 21780 264
rect 21814 230 21848 264
rect 21882 230 21916 264
rect 21950 230 21984 264
rect 22018 230 22052 264
rect 22086 230 22120 264
rect 22154 230 22188 264
rect 22222 230 22256 264
rect 22290 230 22324 264
rect 22358 230 22392 264
rect 22426 230 22460 264
rect 22494 230 22528 264
rect 22562 230 22596 264
rect 22630 230 22664 264
rect 22698 230 22732 264
rect 18 74 52 108
rect 86 74 120 108
rect 154 74 188 108
rect 222 74 256 108
rect 290 74 324 108
rect 358 74 392 108
rect 426 74 460 108
rect 494 74 528 108
rect 562 74 596 108
rect 630 74 664 108
rect 698 74 732 108
rect 766 74 800 108
rect 834 74 868 108
rect 902 74 936 108
rect 970 74 1004 108
rect 1038 74 1072 108
rect 1106 74 1140 108
rect 1174 74 1208 108
rect 1242 74 1276 108
rect 1310 74 1344 108
rect 1378 74 1412 108
rect 1446 74 1480 108
rect 1514 74 1548 108
rect 1582 74 1616 108
rect 1650 74 1684 108
rect 1718 74 1752 108
rect 1786 74 1820 108
rect 1854 74 1888 108
rect 1922 74 1956 108
rect 1990 74 2024 108
rect 2058 74 2092 108
rect 2126 74 2160 108
rect 2194 74 2228 108
rect 2262 74 2296 108
rect 2330 74 2364 108
rect 2398 74 2432 108
rect 2466 74 2500 108
rect 2534 74 2568 108
rect 2602 74 2636 108
rect 2670 74 2704 108
rect 2738 74 2772 108
rect 2806 74 2840 108
rect 2874 74 2908 108
rect 2942 74 2976 108
rect 3010 74 3044 108
rect 3078 74 3112 108
rect 3146 74 3180 108
rect 3214 74 3248 108
rect 3282 74 3316 108
rect 3350 74 3384 108
rect 3418 74 3452 108
rect 3486 74 3520 108
rect 3554 74 3588 108
rect 3622 74 3656 108
rect 3690 74 3724 108
rect 3758 74 3792 108
rect 3826 74 3860 108
rect 3894 74 3928 108
rect 4192 74 4226 108
rect 4260 74 4294 108
rect 4328 74 4362 108
rect 4396 74 4430 108
rect 4464 74 4498 108
rect 4532 74 4566 108
rect 4600 74 4634 108
rect 4668 74 4702 108
rect 4736 74 4770 108
rect 4804 74 4838 108
rect 4872 74 4906 108
rect 4940 74 4974 108
rect 5008 74 5042 108
rect 5076 74 5110 108
rect 5144 74 5178 108
rect 5212 74 5246 108
rect 5280 74 5314 108
rect 5348 74 5382 108
rect 5416 74 5450 108
rect 5484 74 5518 108
rect 5552 74 5586 108
rect 5620 74 5654 108
rect 5688 74 5722 108
rect 5756 74 5790 108
rect 5824 74 5858 108
rect 5892 74 5926 108
rect 5960 74 5994 108
rect 6028 74 6062 108
rect 6096 74 6130 108
rect 6164 74 6198 108
rect 6232 74 6266 108
rect 6300 74 6334 108
rect 6368 74 6402 108
rect 6436 74 6470 108
rect 6504 74 6538 108
rect 6572 74 6606 108
rect 6640 74 6674 108
rect 6708 74 6742 108
rect 6776 74 6810 108
rect 6844 74 6878 108
rect 6912 74 6946 108
rect 6980 74 7014 108
rect 7048 74 7082 108
rect 7116 74 7150 108
rect 7184 74 7218 108
rect 7252 74 7286 108
rect 7320 74 7354 108
rect 7388 74 7422 108
rect 7456 74 7490 108
rect 7524 74 7558 108
rect 7592 74 7626 108
rect 7660 74 7694 108
rect 7728 74 7762 108
rect 7796 74 7830 108
rect 7864 74 7898 108
rect 7932 74 7966 108
rect 8000 74 8034 108
rect 8068 74 8102 108
rect 8318 74 8352 108
rect 8386 74 8420 108
rect 8454 74 8488 108
rect 8522 74 8556 108
rect 8590 74 8624 108
rect 8658 74 8692 108
rect 8726 74 8760 108
rect 8794 74 8828 108
rect 8862 74 8896 108
rect 8930 74 8964 108
rect 8998 74 9032 108
rect 9066 74 9100 108
rect 9134 74 9168 108
rect 9202 74 9236 108
rect 9270 74 9304 108
rect 9338 74 9372 108
rect 9406 74 9440 108
rect 9474 74 9508 108
rect 9542 74 9576 108
rect 9610 74 9644 108
rect 9678 74 9712 108
rect 9746 74 9780 108
rect 9814 74 9848 108
rect 9882 74 9916 108
rect 9950 74 9984 108
rect 10018 74 10052 108
rect 10086 74 10120 108
rect 10154 74 10188 108
rect 10222 74 10256 108
rect 10290 74 10324 108
rect 10358 74 10392 108
rect 10426 74 10460 108
rect 10494 74 10528 108
rect 10562 74 10596 108
rect 10630 74 10664 108
rect 10698 74 10732 108
rect 10766 74 10800 108
rect 10834 74 10868 108
rect 10902 74 10936 108
rect 10970 74 11004 108
rect 11038 74 11072 108
rect 11106 74 11140 108
rect 11174 74 11208 108
rect 11242 74 11276 108
rect 11474 74 11508 108
rect 11542 74 11576 108
rect 11610 74 11644 108
rect 11678 74 11712 108
rect 11746 74 11780 108
rect 11814 74 11848 108
rect 11882 74 11916 108
rect 11950 74 11984 108
rect 12018 74 12052 108
rect 12086 74 12120 108
rect 12154 74 12188 108
rect 12222 74 12256 108
rect 12290 74 12324 108
rect 12358 74 12392 108
rect 12426 74 12460 108
rect 12494 74 12528 108
rect 12562 74 12596 108
rect 12630 74 12664 108
rect 12698 74 12732 108
rect 12766 74 12800 108
rect 12834 74 12868 108
rect 12902 74 12936 108
rect 12970 74 13004 108
rect 13038 74 13072 108
rect 13106 74 13140 108
rect 13174 74 13208 108
rect 13242 74 13276 108
rect 13310 74 13344 108
rect 13378 74 13412 108
rect 13446 74 13480 108
rect 13514 74 13548 108
rect 13582 74 13616 108
rect 13650 74 13684 108
rect 13718 74 13752 108
rect 13786 74 13820 108
rect 13854 74 13888 108
rect 13922 74 13956 108
rect 13990 74 14024 108
rect 14058 74 14092 108
rect 14126 74 14160 108
rect 14194 74 14228 108
rect 14262 74 14296 108
rect 14330 74 14364 108
rect 14398 74 14432 108
rect 14648 74 14682 108
rect 14716 74 14750 108
rect 14784 74 14818 108
rect 14852 74 14886 108
rect 14920 74 14954 108
rect 14988 74 15022 108
rect 15056 74 15090 108
rect 15124 74 15158 108
rect 15192 74 15226 108
rect 15260 74 15294 108
rect 15328 74 15362 108
rect 15396 74 15430 108
rect 15464 74 15498 108
rect 15532 74 15566 108
rect 15600 74 15634 108
rect 15668 74 15702 108
rect 15736 74 15770 108
rect 15804 74 15838 108
rect 15872 74 15906 108
rect 15940 74 15974 108
rect 16008 74 16042 108
rect 16076 74 16110 108
rect 16144 74 16178 108
rect 16212 74 16246 108
rect 16280 74 16314 108
rect 16348 74 16382 108
rect 16416 74 16450 108
rect 16484 74 16518 108
rect 16552 74 16586 108
rect 16620 74 16654 108
rect 16688 74 16722 108
rect 16756 74 16790 108
rect 16824 74 16858 108
rect 16892 74 16926 108
rect 16960 74 16994 108
rect 17028 74 17062 108
rect 17096 74 17130 108
rect 17164 74 17198 108
rect 17232 74 17266 108
rect 17300 74 17334 108
rect 17368 74 17402 108
rect 17436 74 17470 108
rect 17504 74 17538 108
rect 17572 74 17606 108
rect 17640 74 17674 108
rect 17708 74 17742 108
rect 17776 74 17810 108
rect 17844 74 17878 108
rect 17912 74 17946 108
rect 17980 74 18014 108
rect 18048 74 18082 108
rect 18116 74 18150 108
rect 18184 74 18218 108
rect 18252 74 18286 108
rect 18320 74 18354 108
rect 18388 74 18422 108
rect 18456 74 18490 108
rect 18524 74 18558 108
rect 18822 74 18856 108
rect 18890 74 18924 108
rect 18958 74 18992 108
rect 19026 74 19060 108
rect 19094 74 19128 108
rect 19162 74 19196 108
rect 19230 74 19264 108
rect 19298 74 19332 108
rect 19366 74 19400 108
rect 19434 74 19468 108
rect 19502 74 19536 108
rect 19570 74 19604 108
rect 19638 74 19672 108
rect 19706 74 19740 108
rect 19774 74 19808 108
rect 19842 74 19876 108
rect 19910 74 19944 108
rect 19978 74 20012 108
rect 20046 74 20080 108
rect 20114 74 20148 108
rect 20182 74 20216 108
rect 20250 74 20284 108
rect 20318 74 20352 108
rect 20386 74 20420 108
rect 20454 74 20488 108
rect 20522 74 20556 108
rect 20590 74 20624 108
rect 20658 74 20692 108
rect 20726 74 20760 108
rect 20794 74 20828 108
rect 20862 74 20896 108
rect 20930 74 20964 108
rect 20998 74 21032 108
rect 21066 74 21100 108
rect 21134 74 21168 108
rect 21202 74 21236 108
rect 21270 74 21304 108
rect 21338 74 21372 108
rect 21406 74 21440 108
rect 21474 74 21508 108
rect 21542 74 21576 108
rect 21610 74 21644 108
rect 21678 74 21712 108
rect 21746 74 21780 108
rect 21814 74 21848 108
rect 21882 74 21916 108
rect 21950 74 21984 108
rect 22018 74 22052 108
rect 22086 74 22120 108
rect 22154 74 22188 108
rect 22222 74 22256 108
rect 22290 74 22324 108
rect 22358 74 22392 108
rect 22426 74 22460 108
rect 22494 74 22528 108
rect 22562 74 22596 108
rect 22630 74 22664 108
rect 22698 74 22732 108
<< poly >>
rect -86 119 -60 219
rect 3940 187 4046 219
rect 3940 153 3989 187
rect 4023 153 4046 187
rect 3940 119 4046 153
rect 4088 119 4114 219
rect 8114 187 8220 219
rect 8114 153 8163 187
rect 8197 153 8220 187
rect 8114 119 8220 153
rect 8262 119 8288 219
rect 11288 187 11394 219
rect 11288 153 11337 187
rect 11371 153 11394 187
rect 11288 119 11394 153
rect 11436 119 11462 219
rect 14462 187 14568 219
rect 14462 153 14511 187
rect 14545 153 14568 187
rect 14462 119 14568 153
rect 14610 119 14636 219
rect 18636 187 18742 219
rect 18636 153 18685 187
rect 18719 153 18742 187
rect 18636 119 18742 153
rect 18784 119 18810 219
rect 22810 187 22916 219
rect 22810 153 22859 187
rect 22893 153 22916 187
rect 22810 119 22916 153
rect 3966 85 3989 119
rect 4023 85 4046 119
rect 3966 69 4046 85
rect 8140 85 8163 119
rect 8197 85 8220 119
rect 8140 69 8220 85
rect 11314 85 11337 119
rect 11371 85 11394 119
rect 11314 69 11394 85
rect 14488 85 14511 119
rect 14545 85 14568 119
rect 14488 69 14568 85
rect 18662 85 18685 119
rect 18719 85 18742 119
rect 18662 69 18742 85
rect 22836 85 22859 119
rect 22893 85 22916 119
rect 22836 69 22916 85
<< polycont >>
rect 3989 153 4023 187
rect 8163 153 8197 187
rect 11337 153 11371 187
rect 14511 153 14545 187
rect 18685 153 18719 187
rect 22859 153 22893 187
rect 3989 85 4023 119
rect 8163 85 8197 119
rect 11337 85 11371 119
rect 14511 85 14545 119
rect 18685 85 18719 119
rect 22859 85 22893 119
<< locali >>
rect -16 230 18 264
rect 56 230 86 264
rect 128 230 154 264
rect 200 230 222 264
rect 272 230 290 264
rect 344 230 358 264
rect 416 230 426 264
rect 488 230 494 264
rect 560 230 562 264
rect 596 230 598 264
rect 664 230 670 264
rect 732 230 742 264
rect 800 230 814 264
rect 868 230 886 264
rect 936 230 958 264
rect 1004 230 1030 264
rect 1072 230 1102 264
rect 1140 230 1174 264
rect 1208 230 1242 264
rect 1280 230 1310 264
rect 1352 230 1378 264
rect 1424 230 1446 264
rect 1496 230 1514 264
rect 1568 230 1582 264
rect 1640 230 1650 264
rect 1712 230 1718 264
rect 1784 230 1786 264
rect 1820 230 1822 264
rect 1888 230 1894 264
rect 1956 230 1966 264
rect 2024 230 2038 264
rect 2092 230 2110 264
rect 2160 230 2182 264
rect 2228 230 2254 264
rect 2296 230 2326 264
rect 2364 230 2398 264
rect 2432 230 2466 264
rect 2504 230 2534 264
rect 2576 230 2602 264
rect 2648 230 2670 264
rect 2720 230 2738 264
rect 2792 230 2806 264
rect 2864 230 2874 264
rect 2936 230 2942 264
rect 3008 230 3010 264
rect 3044 230 3046 264
rect 3112 230 3118 264
rect 3180 230 3190 264
rect 3248 230 3262 264
rect 3316 230 3334 264
rect 3384 230 3406 264
rect 3452 230 3478 264
rect 3520 230 3550 264
rect 3588 230 3622 264
rect 3656 230 3690 264
rect 3728 230 3758 264
rect 3800 230 3826 264
rect 3872 230 3894 264
rect 4158 230 4192 264
rect 4230 230 4260 264
rect 4302 230 4328 264
rect 4374 230 4396 264
rect 4446 230 4464 264
rect 4518 230 4532 264
rect 4590 230 4600 264
rect 4662 230 4668 264
rect 4734 230 4736 264
rect 4770 230 4772 264
rect 4838 230 4844 264
rect 4906 230 4916 264
rect 4974 230 4988 264
rect 5042 230 5060 264
rect 5110 230 5132 264
rect 5178 230 5204 264
rect 5246 230 5276 264
rect 5314 230 5348 264
rect 5382 230 5416 264
rect 5454 230 5484 264
rect 5526 230 5552 264
rect 5598 230 5620 264
rect 5670 230 5688 264
rect 5742 230 5756 264
rect 5814 230 5824 264
rect 5886 230 5892 264
rect 5958 230 5960 264
rect 5994 230 5996 264
rect 6062 230 6068 264
rect 6130 230 6140 264
rect 6198 230 6212 264
rect 6266 230 6284 264
rect 6334 230 6356 264
rect 6402 230 6428 264
rect 6470 230 6500 264
rect 6538 230 6572 264
rect 6606 230 6640 264
rect 6678 230 6708 264
rect 6750 230 6776 264
rect 6822 230 6844 264
rect 6894 230 6912 264
rect 6966 230 6980 264
rect 7038 230 7048 264
rect 7110 230 7116 264
rect 7182 230 7184 264
rect 7218 230 7220 264
rect 7286 230 7292 264
rect 7354 230 7364 264
rect 7422 230 7436 264
rect 7490 230 7508 264
rect 7558 230 7580 264
rect 7626 230 7652 264
rect 7694 230 7724 264
rect 7762 230 7796 264
rect 7830 230 7864 264
rect 7902 230 7932 264
rect 7974 230 8000 264
rect 8046 230 8068 264
rect 8302 230 8306 264
rect 8352 230 8378 264
rect 8420 230 8450 264
rect 8488 230 8522 264
rect 8556 230 8590 264
rect 8628 230 8658 264
rect 8700 230 8726 264
rect 8772 230 8794 264
rect 8844 230 8862 264
rect 8916 230 8930 264
rect 8988 230 8998 264
rect 9060 230 9066 264
rect 9132 230 9134 264
rect 9168 230 9170 264
rect 9236 230 9242 264
rect 9304 230 9314 264
rect 9372 230 9386 264
rect 9440 230 9458 264
rect 9508 230 9530 264
rect 9576 230 9602 264
rect 9644 230 9674 264
rect 9712 230 9746 264
rect 9780 230 9814 264
rect 9852 230 9882 264
rect 9924 230 9950 264
rect 9996 230 10018 264
rect 10068 230 10086 264
rect 10140 230 10154 264
rect 10212 230 10222 264
rect 10284 230 10290 264
rect 10356 230 10358 264
rect 10392 230 10394 264
rect 10460 230 10466 264
rect 10528 230 10538 264
rect 10596 230 10610 264
rect 10664 230 10682 264
rect 10732 230 10754 264
rect 10800 230 10826 264
rect 10868 230 10898 264
rect 10936 230 10970 264
rect 11004 230 11038 264
rect 11076 230 11106 264
rect 11148 230 11174 264
rect 11220 230 11242 264
rect 11508 230 11530 264
rect 11576 230 11602 264
rect 11644 230 11674 264
rect 11712 230 11746 264
rect 11780 230 11814 264
rect 11852 230 11882 264
rect 11924 230 11950 264
rect 11996 230 12018 264
rect 12068 230 12086 264
rect 12140 230 12154 264
rect 12212 230 12222 264
rect 12284 230 12290 264
rect 12356 230 12358 264
rect 12392 230 12394 264
rect 12460 230 12466 264
rect 12528 230 12538 264
rect 12596 230 12610 264
rect 12664 230 12682 264
rect 12732 230 12754 264
rect 12800 230 12826 264
rect 12868 230 12898 264
rect 12936 230 12970 264
rect 13004 230 13038 264
rect 13076 230 13106 264
rect 13148 230 13174 264
rect 13220 230 13242 264
rect 13292 230 13310 264
rect 13364 230 13378 264
rect 13436 230 13446 264
rect 13508 230 13514 264
rect 13580 230 13582 264
rect 13616 230 13618 264
rect 13684 230 13690 264
rect 13752 230 13762 264
rect 13820 230 13834 264
rect 13888 230 13906 264
rect 13956 230 13978 264
rect 14024 230 14050 264
rect 14092 230 14122 264
rect 14160 230 14194 264
rect 14228 230 14262 264
rect 14300 230 14330 264
rect 14372 230 14398 264
rect 14444 230 14448 264
rect 14682 230 14704 264
rect 14750 230 14776 264
rect 14818 230 14848 264
rect 14886 230 14920 264
rect 14954 230 14988 264
rect 15026 230 15056 264
rect 15098 230 15124 264
rect 15170 230 15192 264
rect 15242 230 15260 264
rect 15314 230 15328 264
rect 15386 230 15396 264
rect 15458 230 15464 264
rect 15530 230 15532 264
rect 15566 230 15568 264
rect 15634 230 15640 264
rect 15702 230 15712 264
rect 15770 230 15784 264
rect 15838 230 15856 264
rect 15906 230 15928 264
rect 15974 230 16000 264
rect 16042 230 16072 264
rect 16110 230 16144 264
rect 16178 230 16212 264
rect 16250 230 16280 264
rect 16322 230 16348 264
rect 16394 230 16416 264
rect 16466 230 16484 264
rect 16538 230 16552 264
rect 16610 230 16620 264
rect 16682 230 16688 264
rect 16754 230 16756 264
rect 16790 230 16792 264
rect 16858 230 16864 264
rect 16926 230 16936 264
rect 16994 230 17008 264
rect 17062 230 17080 264
rect 17130 230 17152 264
rect 17198 230 17224 264
rect 17266 230 17296 264
rect 17334 230 17368 264
rect 17402 230 17436 264
rect 17474 230 17504 264
rect 17546 230 17572 264
rect 17618 230 17640 264
rect 17690 230 17708 264
rect 17762 230 17776 264
rect 17834 230 17844 264
rect 17906 230 17912 264
rect 17978 230 17980 264
rect 18014 230 18016 264
rect 18082 230 18088 264
rect 18150 230 18160 264
rect 18218 230 18232 264
rect 18286 230 18304 264
rect 18354 230 18376 264
rect 18422 230 18448 264
rect 18490 230 18520 264
rect 18558 230 18592 264
rect 18856 230 18878 264
rect 18924 230 18950 264
rect 18992 230 19022 264
rect 19060 230 19094 264
rect 19128 230 19162 264
rect 19200 230 19230 264
rect 19272 230 19298 264
rect 19344 230 19366 264
rect 19416 230 19434 264
rect 19488 230 19502 264
rect 19560 230 19570 264
rect 19632 230 19638 264
rect 19704 230 19706 264
rect 19740 230 19742 264
rect 19808 230 19814 264
rect 19876 230 19886 264
rect 19944 230 19958 264
rect 20012 230 20030 264
rect 20080 230 20102 264
rect 20148 230 20174 264
rect 20216 230 20246 264
rect 20284 230 20318 264
rect 20352 230 20386 264
rect 20424 230 20454 264
rect 20496 230 20522 264
rect 20568 230 20590 264
rect 20640 230 20658 264
rect 20712 230 20726 264
rect 20784 230 20794 264
rect 20856 230 20862 264
rect 20928 230 20930 264
rect 20964 230 20966 264
rect 21032 230 21038 264
rect 21100 230 21110 264
rect 21168 230 21182 264
rect 21236 230 21254 264
rect 21304 230 21326 264
rect 21372 230 21398 264
rect 21440 230 21470 264
rect 21508 230 21542 264
rect 21576 230 21610 264
rect 21648 230 21678 264
rect 21720 230 21746 264
rect 21792 230 21814 264
rect 21864 230 21882 264
rect 21936 230 21950 264
rect 22008 230 22018 264
rect 22080 230 22086 264
rect 22152 230 22154 264
rect 22188 230 22190 264
rect 22256 230 22262 264
rect 22324 230 22334 264
rect 22392 230 22406 264
rect 22460 230 22478 264
rect 22528 230 22550 264
rect 22596 230 22622 264
rect 22664 230 22694 264
rect 22732 230 22766 264
rect 3982 189 4030 203
rect 8156 189 8204 203
rect 11330 189 11378 203
rect 14504 189 14552 203
rect 18678 189 18726 203
rect 22852 189 22900 203
rect 4016 187 4054 189
rect 4023 155 4054 187
rect 8190 187 8228 189
rect 8197 155 8228 187
rect 11364 187 11402 189
rect 11371 155 11402 187
rect 14509 187 14547 189
rect 14509 155 14511 187
rect 3982 153 3989 155
rect 4023 153 4030 155
rect 3982 119 4030 153
rect -16 74 18 108
rect 56 74 86 108
rect 128 74 154 108
rect 200 74 222 108
rect 272 74 290 108
rect 344 74 358 108
rect 416 74 426 108
rect 488 74 494 108
rect 560 74 562 108
rect 596 74 598 108
rect 664 74 670 108
rect 732 74 742 108
rect 800 74 814 108
rect 868 74 886 108
rect 936 74 958 108
rect 1004 74 1030 108
rect 1072 74 1102 108
rect 1140 74 1174 108
rect 1208 74 1242 108
rect 1280 74 1310 108
rect 1352 74 1378 108
rect 1424 74 1446 108
rect 1496 74 1514 108
rect 1568 74 1582 108
rect 1640 74 1650 108
rect 1712 74 1718 108
rect 1784 74 1786 108
rect 1820 74 1822 108
rect 1888 74 1894 108
rect 1956 74 1966 108
rect 2024 74 2038 108
rect 2092 74 2110 108
rect 2160 74 2182 108
rect 2228 74 2254 108
rect 2296 74 2326 108
rect 2364 74 2398 108
rect 2432 74 2466 108
rect 2504 74 2534 108
rect 2576 74 2602 108
rect 2648 74 2670 108
rect 2720 74 2738 108
rect 2792 74 2806 108
rect 2864 74 2874 108
rect 2936 74 2942 108
rect 3008 74 3010 108
rect 3044 74 3046 108
rect 3112 74 3118 108
rect 3180 74 3190 108
rect 3248 74 3262 108
rect 3316 74 3334 108
rect 3384 74 3406 108
rect 3452 74 3478 108
rect 3520 74 3550 108
rect 3588 74 3622 108
rect 3656 74 3690 108
rect 3728 74 3758 108
rect 3800 74 3826 108
rect 3872 74 3894 108
rect 3982 85 3989 119
rect 4023 85 4030 119
rect 8156 153 8163 155
rect 8197 153 8204 155
rect 8156 119 8204 153
rect 3982 69 4030 85
rect 4158 74 4192 108
rect 4230 74 4260 108
rect 4302 74 4328 108
rect 4374 74 4396 108
rect 4446 74 4464 108
rect 4518 74 4532 108
rect 4590 74 4600 108
rect 4662 74 4668 108
rect 4734 74 4736 108
rect 4770 74 4772 108
rect 4838 74 4844 108
rect 4906 74 4916 108
rect 4974 74 4988 108
rect 5042 74 5060 108
rect 5110 74 5132 108
rect 5178 74 5204 108
rect 5246 74 5276 108
rect 5314 74 5348 108
rect 5382 74 5416 108
rect 5454 74 5484 108
rect 5526 74 5552 108
rect 5598 74 5620 108
rect 5670 74 5688 108
rect 5742 74 5756 108
rect 5814 74 5824 108
rect 5886 74 5892 108
rect 5958 74 5960 108
rect 5994 74 5996 108
rect 6062 74 6068 108
rect 6130 74 6140 108
rect 6198 74 6212 108
rect 6266 74 6284 108
rect 6334 74 6356 108
rect 6402 74 6428 108
rect 6470 74 6500 108
rect 6538 74 6572 108
rect 6606 74 6640 108
rect 6678 74 6708 108
rect 6750 74 6776 108
rect 6822 74 6844 108
rect 6894 74 6912 108
rect 6966 74 6980 108
rect 7038 74 7048 108
rect 7110 74 7116 108
rect 7182 74 7184 108
rect 7218 74 7220 108
rect 7286 74 7292 108
rect 7354 74 7364 108
rect 7422 74 7436 108
rect 7490 74 7508 108
rect 7558 74 7580 108
rect 7626 74 7652 108
rect 7694 74 7724 108
rect 7762 74 7796 108
rect 7830 74 7864 108
rect 7902 74 7932 108
rect 7974 74 8000 108
rect 8046 74 8068 108
rect 8156 85 8163 119
rect 8197 85 8204 119
rect 11330 153 11337 155
rect 11371 153 11378 155
rect 11330 119 11378 153
rect 8156 69 8204 85
rect 8302 74 8306 108
rect 8352 74 8378 108
rect 8420 74 8450 108
rect 8488 74 8522 108
rect 8556 74 8590 108
rect 8628 74 8658 108
rect 8700 74 8726 108
rect 8772 74 8794 108
rect 8844 74 8862 108
rect 8916 74 8930 108
rect 8988 74 8998 108
rect 9060 74 9066 108
rect 9132 74 9134 108
rect 9168 74 9170 108
rect 9236 74 9242 108
rect 9304 74 9314 108
rect 9372 74 9386 108
rect 9440 74 9458 108
rect 9508 74 9530 108
rect 9576 74 9602 108
rect 9644 74 9674 108
rect 9712 74 9746 108
rect 9780 74 9814 108
rect 9852 74 9882 108
rect 9924 74 9950 108
rect 9996 74 10018 108
rect 10068 74 10086 108
rect 10140 74 10154 108
rect 10212 74 10222 108
rect 10284 74 10290 108
rect 10356 74 10358 108
rect 10392 74 10394 108
rect 10460 74 10466 108
rect 10528 74 10538 108
rect 10596 74 10610 108
rect 10664 74 10682 108
rect 10732 74 10754 108
rect 10800 74 10826 108
rect 10868 74 10898 108
rect 10936 74 10970 108
rect 11004 74 11038 108
rect 11076 74 11106 108
rect 11148 74 11174 108
rect 11220 74 11242 108
rect 11330 85 11337 119
rect 11371 85 11378 119
rect 14504 153 14511 155
rect 14545 155 14547 187
rect 18651 187 18691 189
rect 18651 155 18685 187
rect 18725 155 18726 189
rect 22828 187 22866 189
rect 22828 155 22859 187
rect 14545 153 14552 155
rect 14504 119 14552 153
rect 11330 69 11378 85
rect 11508 74 11530 108
rect 11576 74 11602 108
rect 11644 74 11674 108
rect 11712 74 11746 108
rect 11780 74 11814 108
rect 11852 74 11882 108
rect 11924 74 11950 108
rect 11996 74 12018 108
rect 12068 74 12086 108
rect 12140 74 12154 108
rect 12212 74 12222 108
rect 12284 74 12290 108
rect 12356 74 12358 108
rect 12392 74 12394 108
rect 12460 74 12466 108
rect 12528 74 12538 108
rect 12596 74 12610 108
rect 12664 74 12682 108
rect 12732 74 12754 108
rect 12800 74 12826 108
rect 12868 74 12898 108
rect 12936 74 12970 108
rect 13004 74 13038 108
rect 13076 74 13106 108
rect 13148 74 13174 108
rect 13220 74 13242 108
rect 13292 74 13310 108
rect 13364 74 13378 108
rect 13436 74 13446 108
rect 13508 74 13514 108
rect 13580 74 13582 108
rect 13616 74 13618 108
rect 13684 74 13690 108
rect 13752 74 13762 108
rect 13820 74 13834 108
rect 13888 74 13906 108
rect 13956 74 13978 108
rect 14024 74 14050 108
rect 14092 74 14122 108
rect 14160 74 14194 108
rect 14228 74 14262 108
rect 14300 74 14330 108
rect 14372 74 14398 108
rect 14444 74 14448 108
rect 14504 85 14511 119
rect 14545 85 14552 119
rect 18678 153 18685 155
rect 18719 153 18726 155
rect 18678 119 18726 153
rect 14504 69 14552 85
rect 14682 74 14704 108
rect 14750 74 14776 108
rect 14818 74 14848 108
rect 14886 74 14920 108
rect 14954 74 14988 108
rect 15026 74 15056 108
rect 15098 74 15124 108
rect 15170 74 15192 108
rect 15242 74 15260 108
rect 15314 74 15328 108
rect 15386 74 15396 108
rect 15458 74 15464 108
rect 15530 74 15532 108
rect 15566 74 15568 108
rect 15634 74 15640 108
rect 15702 74 15712 108
rect 15770 74 15784 108
rect 15838 74 15856 108
rect 15906 74 15928 108
rect 15974 74 16000 108
rect 16042 74 16072 108
rect 16110 74 16144 108
rect 16178 74 16212 108
rect 16250 74 16280 108
rect 16322 74 16348 108
rect 16394 74 16416 108
rect 16466 74 16484 108
rect 16538 74 16552 108
rect 16610 74 16620 108
rect 16682 74 16688 108
rect 16754 74 16756 108
rect 16790 74 16792 108
rect 16858 74 16864 108
rect 16926 74 16936 108
rect 16994 74 17008 108
rect 17062 74 17080 108
rect 17130 74 17152 108
rect 17198 74 17224 108
rect 17266 74 17296 108
rect 17334 74 17368 108
rect 17402 74 17436 108
rect 17474 74 17504 108
rect 17546 74 17572 108
rect 17618 74 17640 108
rect 17690 74 17708 108
rect 17762 74 17776 108
rect 17834 74 17844 108
rect 17906 74 17912 108
rect 17978 74 17980 108
rect 18014 74 18016 108
rect 18082 74 18088 108
rect 18150 74 18160 108
rect 18218 74 18232 108
rect 18286 74 18304 108
rect 18354 74 18376 108
rect 18422 74 18448 108
rect 18490 74 18520 108
rect 18558 74 18592 108
rect 18678 85 18685 119
rect 18719 85 18726 119
rect 22852 153 22859 155
rect 22893 153 22900 155
rect 22852 119 22900 153
rect 18678 69 18726 85
rect 18856 74 18878 108
rect 18924 74 18950 108
rect 18992 74 19022 108
rect 19060 74 19094 108
rect 19128 74 19162 108
rect 19200 74 19230 108
rect 19272 74 19298 108
rect 19344 74 19366 108
rect 19416 74 19434 108
rect 19488 74 19502 108
rect 19560 74 19570 108
rect 19632 74 19638 108
rect 19704 74 19706 108
rect 19740 74 19742 108
rect 19808 74 19814 108
rect 19876 74 19886 108
rect 19944 74 19958 108
rect 20012 74 20030 108
rect 20080 74 20102 108
rect 20148 74 20174 108
rect 20216 74 20246 108
rect 20284 74 20318 108
rect 20352 74 20386 108
rect 20424 74 20454 108
rect 20496 74 20522 108
rect 20568 74 20590 108
rect 20640 74 20658 108
rect 20712 74 20726 108
rect 20784 74 20794 108
rect 20856 74 20862 108
rect 20928 74 20930 108
rect 20964 74 20966 108
rect 21032 74 21038 108
rect 21100 74 21110 108
rect 21168 74 21182 108
rect 21236 74 21254 108
rect 21304 74 21326 108
rect 21372 74 21398 108
rect 21440 74 21470 108
rect 21508 74 21542 108
rect 21576 74 21610 108
rect 21648 74 21678 108
rect 21720 74 21746 108
rect 21792 74 21814 108
rect 21864 74 21882 108
rect 21936 74 21950 108
rect 22008 74 22018 108
rect 22080 74 22086 108
rect 22152 74 22154 108
rect 22188 74 22190 108
rect 22256 74 22262 108
rect 22324 74 22334 108
rect 22392 74 22406 108
rect 22460 74 22478 108
rect 22528 74 22550 108
rect 22596 74 22622 108
rect 22664 74 22694 108
rect 22732 74 22766 108
rect 22852 85 22859 119
rect 22893 85 22900 119
rect 22852 69 22900 85
<< viali >>
rect -50 230 -16 264
rect 22 230 52 264
rect 52 230 56 264
rect 94 230 120 264
rect 120 230 128 264
rect 166 230 188 264
rect 188 230 200 264
rect 238 230 256 264
rect 256 230 272 264
rect 310 230 324 264
rect 324 230 344 264
rect 382 230 392 264
rect 392 230 416 264
rect 454 230 460 264
rect 460 230 488 264
rect 526 230 528 264
rect 528 230 560 264
rect 598 230 630 264
rect 630 230 632 264
rect 670 230 698 264
rect 698 230 704 264
rect 742 230 766 264
rect 766 230 776 264
rect 814 230 834 264
rect 834 230 848 264
rect 886 230 902 264
rect 902 230 920 264
rect 958 230 970 264
rect 970 230 992 264
rect 1030 230 1038 264
rect 1038 230 1064 264
rect 1102 230 1106 264
rect 1106 230 1136 264
rect 1174 230 1208 264
rect 1246 230 1276 264
rect 1276 230 1280 264
rect 1318 230 1344 264
rect 1344 230 1352 264
rect 1390 230 1412 264
rect 1412 230 1424 264
rect 1462 230 1480 264
rect 1480 230 1496 264
rect 1534 230 1548 264
rect 1548 230 1568 264
rect 1606 230 1616 264
rect 1616 230 1640 264
rect 1678 230 1684 264
rect 1684 230 1712 264
rect 1750 230 1752 264
rect 1752 230 1784 264
rect 1822 230 1854 264
rect 1854 230 1856 264
rect 1894 230 1922 264
rect 1922 230 1928 264
rect 1966 230 1990 264
rect 1990 230 2000 264
rect 2038 230 2058 264
rect 2058 230 2072 264
rect 2110 230 2126 264
rect 2126 230 2144 264
rect 2182 230 2194 264
rect 2194 230 2216 264
rect 2254 230 2262 264
rect 2262 230 2288 264
rect 2326 230 2330 264
rect 2330 230 2360 264
rect 2398 230 2432 264
rect 2470 230 2500 264
rect 2500 230 2504 264
rect 2542 230 2568 264
rect 2568 230 2576 264
rect 2614 230 2636 264
rect 2636 230 2648 264
rect 2686 230 2704 264
rect 2704 230 2720 264
rect 2758 230 2772 264
rect 2772 230 2792 264
rect 2830 230 2840 264
rect 2840 230 2864 264
rect 2902 230 2908 264
rect 2908 230 2936 264
rect 2974 230 2976 264
rect 2976 230 3008 264
rect 3046 230 3078 264
rect 3078 230 3080 264
rect 3118 230 3146 264
rect 3146 230 3152 264
rect 3190 230 3214 264
rect 3214 230 3224 264
rect 3262 230 3282 264
rect 3282 230 3296 264
rect 3334 230 3350 264
rect 3350 230 3368 264
rect 3406 230 3418 264
rect 3418 230 3440 264
rect 3478 230 3486 264
rect 3486 230 3512 264
rect 3550 230 3554 264
rect 3554 230 3584 264
rect 3622 230 3656 264
rect 3694 230 3724 264
rect 3724 230 3728 264
rect 3766 230 3792 264
rect 3792 230 3800 264
rect 3838 230 3860 264
rect 3860 230 3872 264
rect 3910 230 3928 264
rect 3928 230 3944 264
rect 4124 230 4158 264
rect 4196 230 4226 264
rect 4226 230 4230 264
rect 4268 230 4294 264
rect 4294 230 4302 264
rect 4340 230 4362 264
rect 4362 230 4374 264
rect 4412 230 4430 264
rect 4430 230 4446 264
rect 4484 230 4498 264
rect 4498 230 4518 264
rect 4556 230 4566 264
rect 4566 230 4590 264
rect 4628 230 4634 264
rect 4634 230 4662 264
rect 4700 230 4702 264
rect 4702 230 4734 264
rect 4772 230 4804 264
rect 4804 230 4806 264
rect 4844 230 4872 264
rect 4872 230 4878 264
rect 4916 230 4940 264
rect 4940 230 4950 264
rect 4988 230 5008 264
rect 5008 230 5022 264
rect 5060 230 5076 264
rect 5076 230 5094 264
rect 5132 230 5144 264
rect 5144 230 5166 264
rect 5204 230 5212 264
rect 5212 230 5238 264
rect 5276 230 5280 264
rect 5280 230 5310 264
rect 5348 230 5382 264
rect 5420 230 5450 264
rect 5450 230 5454 264
rect 5492 230 5518 264
rect 5518 230 5526 264
rect 5564 230 5586 264
rect 5586 230 5598 264
rect 5636 230 5654 264
rect 5654 230 5670 264
rect 5708 230 5722 264
rect 5722 230 5742 264
rect 5780 230 5790 264
rect 5790 230 5814 264
rect 5852 230 5858 264
rect 5858 230 5886 264
rect 5924 230 5926 264
rect 5926 230 5958 264
rect 5996 230 6028 264
rect 6028 230 6030 264
rect 6068 230 6096 264
rect 6096 230 6102 264
rect 6140 230 6164 264
rect 6164 230 6174 264
rect 6212 230 6232 264
rect 6232 230 6246 264
rect 6284 230 6300 264
rect 6300 230 6318 264
rect 6356 230 6368 264
rect 6368 230 6390 264
rect 6428 230 6436 264
rect 6436 230 6462 264
rect 6500 230 6504 264
rect 6504 230 6534 264
rect 6572 230 6606 264
rect 6644 230 6674 264
rect 6674 230 6678 264
rect 6716 230 6742 264
rect 6742 230 6750 264
rect 6788 230 6810 264
rect 6810 230 6822 264
rect 6860 230 6878 264
rect 6878 230 6894 264
rect 6932 230 6946 264
rect 6946 230 6966 264
rect 7004 230 7014 264
rect 7014 230 7038 264
rect 7076 230 7082 264
rect 7082 230 7110 264
rect 7148 230 7150 264
rect 7150 230 7182 264
rect 7220 230 7252 264
rect 7252 230 7254 264
rect 7292 230 7320 264
rect 7320 230 7326 264
rect 7364 230 7388 264
rect 7388 230 7398 264
rect 7436 230 7456 264
rect 7456 230 7470 264
rect 7508 230 7524 264
rect 7524 230 7542 264
rect 7580 230 7592 264
rect 7592 230 7614 264
rect 7652 230 7660 264
rect 7660 230 7686 264
rect 7724 230 7728 264
rect 7728 230 7758 264
rect 7796 230 7830 264
rect 7868 230 7898 264
rect 7898 230 7902 264
rect 7940 230 7966 264
rect 7966 230 7974 264
rect 8012 230 8034 264
rect 8034 230 8046 264
rect 8084 230 8102 264
rect 8102 230 8118 264
rect 8306 230 8318 264
rect 8318 230 8340 264
rect 8378 230 8386 264
rect 8386 230 8412 264
rect 8450 230 8454 264
rect 8454 230 8484 264
rect 8522 230 8556 264
rect 8594 230 8624 264
rect 8624 230 8628 264
rect 8666 230 8692 264
rect 8692 230 8700 264
rect 8738 230 8760 264
rect 8760 230 8772 264
rect 8810 230 8828 264
rect 8828 230 8844 264
rect 8882 230 8896 264
rect 8896 230 8916 264
rect 8954 230 8964 264
rect 8964 230 8988 264
rect 9026 230 9032 264
rect 9032 230 9060 264
rect 9098 230 9100 264
rect 9100 230 9132 264
rect 9170 230 9202 264
rect 9202 230 9204 264
rect 9242 230 9270 264
rect 9270 230 9276 264
rect 9314 230 9338 264
rect 9338 230 9348 264
rect 9386 230 9406 264
rect 9406 230 9420 264
rect 9458 230 9474 264
rect 9474 230 9492 264
rect 9530 230 9542 264
rect 9542 230 9564 264
rect 9602 230 9610 264
rect 9610 230 9636 264
rect 9674 230 9678 264
rect 9678 230 9708 264
rect 9746 230 9780 264
rect 9818 230 9848 264
rect 9848 230 9852 264
rect 9890 230 9916 264
rect 9916 230 9924 264
rect 9962 230 9984 264
rect 9984 230 9996 264
rect 10034 230 10052 264
rect 10052 230 10068 264
rect 10106 230 10120 264
rect 10120 230 10140 264
rect 10178 230 10188 264
rect 10188 230 10212 264
rect 10250 230 10256 264
rect 10256 230 10284 264
rect 10322 230 10324 264
rect 10324 230 10356 264
rect 10394 230 10426 264
rect 10426 230 10428 264
rect 10466 230 10494 264
rect 10494 230 10500 264
rect 10538 230 10562 264
rect 10562 230 10572 264
rect 10610 230 10630 264
rect 10630 230 10644 264
rect 10682 230 10698 264
rect 10698 230 10716 264
rect 10754 230 10766 264
rect 10766 230 10788 264
rect 10826 230 10834 264
rect 10834 230 10860 264
rect 10898 230 10902 264
rect 10902 230 10932 264
rect 10970 230 11004 264
rect 11042 230 11072 264
rect 11072 230 11076 264
rect 11114 230 11140 264
rect 11140 230 11148 264
rect 11186 230 11208 264
rect 11208 230 11220 264
rect 11258 230 11276 264
rect 11276 230 11292 264
rect 11458 230 11474 264
rect 11474 230 11492 264
rect 11530 230 11542 264
rect 11542 230 11564 264
rect 11602 230 11610 264
rect 11610 230 11636 264
rect 11674 230 11678 264
rect 11678 230 11708 264
rect 11746 230 11780 264
rect 11818 230 11848 264
rect 11848 230 11852 264
rect 11890 230 11916 264
rect 11916 230 11924 264
rect 11962 230 11984 264
rect 11984 230 11996 264
rect 12034 230 12052 264
rect 12052 230 12068 264
rect 12106 230 12120 264
rect 12120 230 12140 264
rect 12178 230 12188 264
rect 12188 230 12212 264
rect 12250 230 12256 264
rect 12256 230 12284 264
rect 12322 230 12324 264
rect 12324 230 12356 264
rect 12394 230 12426 264
rect 12426 230 12428 264
rect 12466 230 12494 264
rect 12494 230 12500 264
rect 12538 230 12562 264
rect 12562 230 12572 264
rect 12610 230 12630 264
rect 12630 230 12644 264
rect 12682 230 12698 264
rect 12698 230 12716 264
rect 12754 230 12766 264
rect 12766 230 12788 264
rect 12826 230 12834 264
rect 12834 230 12860 264
rect 12898 230 12902 264
rect 12902 230 12932 264
rect 12970 230 13004 264
rect 13042 230 13072 264
rect 13072 230 13076 264
rect 13114 230 13140 264
rect 13140 230 13148 264
rect 13186 230 13208 264
rect 13208 230 13220 264
rect 13258 230 13276 264
rect 13276 230 13292 264
rect 13330 230 13344 264
rect 13344 230 13364 264
rect 13402 230 13412 264
rect 13412 230 13436 264
rect 13474 230 13480 264
rect 13480 230 13508 264
rect 13546 230 13548 264
rect 13548 230 13580 264
rect 13618 230 13650 264
rect 13650 230 13652 264
rect 13690 230 13718 264
rect 13718 230 13724 264
rect 13762 230 13786 264
rect 13786 230 13796 264
rect 13834 230 13854 264
rect 13854 230 13868 264
rect 13906 230 13922 264
rect 13922 230 13940 264
rect 13978 230 13990 264
rect 13990 230 14012 264
rect 14050 230 14058 264
rect 14058 230 14084 264
rect 14122 230 14126 264
rect 14126 230 14156 264
rect 14194 230 14228 264
rect 14266 230 14296 264
rect 14296 230 14300 264
rect 14338 230 14364 264
rect 14364 230 14372 264
rect 14410 230 14432 264
rect 14432 230 14444 264
rect 14632 230 14648 264
rect 14648 230 14666 264
rect 14704 230 14716 264
rect 14716 230 14738 264
rect 14776 230 14784 264
rect 14784 230 14810 264
rect 14848 230 14852 264
rect 14852 230 14882 264
rect 14920 230 14954 264
rect 14992 230 15022 264
rect 15022 230 15026 264
rect 15064 230 15090 264
rect 15090 230 15098 264
rect 15136 230 15158 264
rect 15158 230 15170 264
rect 15208 230 15226 264
rect 15226 230 15242 264
rect 15280 230 15294 264
rect 15294 230 15314 264
rect 15352 230 15362 264
rect 15362 230 15386 264
rect 15424 230 15430 264
rect 15430 230 15458 264
rect 15496 230 15498 264
rect 15498 230 15530 264
rect 15568 230 15600 264
rect 15600 230 15602 264
rect 15640 230 15668 264
rect 15668 230 15674 264
rect 15712 230 15736 264
rect 15736 230 15746 264
rect 15784 230 15804 264
rect 15804 230 15818 264
rect 15856 230 15872 264
rect 15872 230 15890 264
rect 15928 230 15940 264
rect 15940 230 15962 264
rect 16000 230 16008 264
rect 16008 230 16034 264
rect 16072 230 16076 264
rect 16076 230 16106 264
rect 16144 230 16178 264
rect 16216 230 16246 264
rect 16246 230 16250 264
rect 16288 230 16314 264
rect 16314 230 16322 264
rect 16360 230 16382 264
rect 16382 230 16394 264
rect 16432 230 16450 264
rect 16450 230 16466 264
rect 16504 230 16518 264
rect 16518 230 16538 264
rect 16576 230 16586 264
rect 16586 230 16610 264
rect 16648 230 16654 264
rect 16654 230 16682 264
rect 16720 230 16722 264
rect 16722 230 16754 264
rect 16792 230 16824 264
rect 16824 230 16826 264
rect 16864 230 16892 264
rect 16892 230 16898 264
rect 16936 230 16960 264
rect 16960 230 16970 264
rect 17008 230 17028 264
rect 17028 230 17042 264
rect 17080 230 17096 264
rect 17096 230 17114 264
rect 17152 230 17164 264
rect 17164 230 17186 264
rect 17224 230 17232 264
rect 17232 230 17258 264
rect 17296 230 17300 264
rect 17300 230 17330 264
rect 17368 230 17402 264
rect 17440 230 17470 264
rect 17470 230 17474 264
rect 17512 230 17538 264
rect 17538 230 17546 264
rect 17584 230 17606 264
rect 17606 230 17618 264
rect 17656 230 17674 264
rect 17674 230 17690 264
rect 17728 230 17742 264
rect 17742 230 17762 264
rect 17800 230 17810 264
rect 17810 230 17834 264
rect 17872 230 17878 264
rect 17878 230 17906 264
rect 17944 230 17946 264
rect 17946 230 17978 264
rect 18016 230 18048 264
rect 18048 230 18050 264
rect 18088 230 18116 264
rect 18116 230 18122 264
rect 18160 230 18184 264
rect 18184 230 18194 264
rect 18232 230 18252 264
rect 18252 230 18266 264
rect 18304 230 18320 264
rect 18320 230 18338 264
rect 18376 230 18388 264
rect 18388 230 18410 264
rect 18448 230 18456 264
rect 18456 230 18482 264
rect 18520 230 18524 264
rect 18524 230 18554 264
rect 18592 230 18626 264
rect 18806 230 18822 264
rect 18822 230 18840 264
rect 18878 230 18890 264
rect 18890 230 18912 264
rect 18950 230 18958 264
rect 18958 230 18984 264
rect 19022 230 19026 264
rect 19026 230 19056 264
rect 19094 230 19128 264
rect 19166 230 19196 264
rect 19196 230 19200 264
rect 19238 230 19264 264
rect 19264 230 19272 264
rect 19310 230 19332 264
rect 19332 230 19344 264
rect 19382 230 19400 264
rect 19400 230 19416 264
rect 19454 230 19468 264
rect 19468 230 19488 264
rect 19526 230 19536 264
rect 19536 230 19560 264
rect 19598 230 19604 264
rect 19604 230 19632 264
rect 19670 230 19672 264
rect 19672 230 19704 264
rect 19742 230 19774 264
rect 19774 230 19776 264
rect 19814 230 19842 264
rect 19842 230 19848 264
rect 19886 230 19910 264
rect 19910 230 19920 264
rect 19958 230 19978 264
rect 19978 230 19992 264
rect 20030 230 20046 264
rect 20046 230 20064 264
rect 20102 230 20114 264
rect 20114 230 20136 264
rect 20174 230 20182 264
rect 20182 230 20208 264
rect 20246 230 20250 264
rect 20250 230 20280 264
rect 20318 230 20352 264
rect 20390 230 20420 264
rect 20420 230 20424 264
rect 20462 230 20488 264
rect 20488 230 20496 264
rect 20534 230 20556 264
rect 20556 230 20568 264
rect 20606 230 20624 264
rect 20624 230 20640 264
rect 20678 230 20692 264
rect 20692 230 20712 264
rect 20750 230 20760 264
rect 20760 230 20784 264
rect 20822 230 20828 264
rect 20828 230 20856 264
rect 20894 230 20896 264
rect 20896 230 20928 264
rect 20966 230 20998 264
rect 20998 230 21000 264
rect 21038 230 21066 264
rect 21066 230 21072 264
rect 21110 230 21134 264
rect 21134 230 21144 264
rect 21182 230 21202 264
rect 21202 230 21216 264
rect 21254 230 21270 264
rect 21270 230 21288 264
rect 21326 230 21338 264
rect 21338 230 21360 264
rect 21398 230 21406 264
rect 21406 230 21432 264
rect 21470 230 21474 264
rect 21474 230 21504 264
rect 21542 230 21576 264
rect 21614 230 21644 264
rect 21644 230 21648 264
rect 21686 230 21712 264
rect 21712 230 21720 264
rect 21758 230 21780 264
rect 21780 230 21792 264
rect 21830 230 21848 264
rect 21848 230 21864 264
rect 21902 230 21916 264
rect 21916 230 21936 264
rect 21974 230 21984 264
rect 21984 230 22008 264
rect 22046 230 22052 264
rect 22052 230 22080 264
rect 22118 230 22120 264
rect 22120 230 22152 264
rect 22190 230 22222 264
rect 22222 230 22224 264
rect 22262 230 22290 264
rect 22290 230 22296 264
rect 22334 230 22358 264
rect 22358 230 22368 264
rect 22406 230 22426 264
rect 22426 230 22440 264
rect 22478 230 22494 264
rect 22494 230 22512 264
rect 22550 230 22562 264
rect 22562 230 22584 264
rect 22622 230 22630 264
rect 22630 230 22656 264
rect 22694 230 22698 264
rect 22698 230 22728 264
rect 22766 230 22800 264
rect 3982 187 4016 189
rect 3982 155 3989 187
rect 3989 155 4016 187
rect 4054 155 4088 189
rect 8156 187 8190 189
rect 8156 155 8163 187
rect 8163 155 8190 187
rect 8228 155 8262 189
rect 11330 187 11364 189
rect 11330 155 11337 187
rect 11337 155 11364 187
rect 11402 155 11436 189
rect 14475 155 14509 189
rect -50 74 -16 108
rect 22 74 52 108
rect 52 74 56 108
rect 94 74 120 108
rect 120 74 128 108
rect 166 74 188 108
rect 188 74 200 108
rect 238 74 256 108
rect 256 74 272 108
rect 310 74 324 108
rect 324 74 344 108
rect 382 74 392 108
rect 392 74 416 108
rect 454 74 460 108
rect 460 74 488 108
rect 526 74 528 108
rect 528 74 560 108
rect 598 74 630 108
rect 630 74 632 108
rect 670 74 698 108
rect 698 74 704 108
rect 742 74 766 108
rect 766 74 776 108
rect 814 74 834 108
rect 834 74 848 108
rect 886 74 902 108
rect 902 74 920 108
rect 958 74 970 108
rect 970 74 992 108
rect 1030 74 1038 108
rect 1038 74 1064 108
rect 1102 74 1106 108
rect 1106 74 1136 108
rect 1174 74 1208 108
rect 1246 74 1276 108
rect 1276 74 1280 108
rect 1318 74 1344 108
rect 1344 74 1352 108
rect 1390 74 1412 108
rect 1412 74 1424 108
rect 1462 74 1480 108
rect 1480 74 1496 108
rect 1534 74 1548 108
rect 1548 74 1568 108
rect 1606 74 1616 108
rect 1616 74 1640 108
rect 1678 74 1684 108
rect 1684 74 1712 108
rect 1750 74 1752 108
rect 1752 74 1784 108
rect 1822 74 1854 108
rect 1854 74 1856 108
rect 1894 74 1922 108
rect 1922 74 1928 108
rect 1966 74 1990 108
rect 1990 74 2000 108
rect 2038 74 2058 108
rect 2058 74 2072 108
rect 2110 74 2126 108
rect 2126 74 2144 108
rect 2182 74 2194 108
rect 2194 74 2216 108
rect 2254 74 2262 108
rect 2262 74 2288 108
rect 2326 74 2330 108
rect 2330 74 2360 108
rect 2398 74 2432 108
rect 2470 74 2500 108
rect 2500 74 2504 108
rect 2542 74 2568 108
rect 2568 74 2576 108
rect 2614 74 2636 108
rect 2636 74 2648 108
rect 2686 74 2704 108
rect 2704 74 2720 108
rect 2758 74 2772 108
rect 2772 74 2792 108
rect 2830 74 2840 108
rect 2840 74 2864 108
rect 2902 74 2908 108
rect 2908 74 2936 108
rect 2974 74 2976 108
rect 2976 74 3008 108
rect 3046 74 3078 108
rect 3078 74 3080 108
rect 3118 74 3146 108
rect 3146 74 3152 108
rect 3190 74 3214 108
rect 3214 74 3224 108
rect 3262 74 3282 108
rect 3282 74 3296 108
rect 3334 74 3350 108
rect 3350 74 3368 108
rect 3406 74 3418 108
rect 3418 74 3440 108
rect 3478 74 3486 108
rect 3486 74 3512 108
rect 3550 74 3554 108
rect 3554 74 3584 108
rect 3622 74 3656 108
rect 3694 74 3724 108
rect 3724 74 3728 108
rect 3766 74 3792 108
rect 3792 74 3800 108
rect 3838 74 3860 108
rect 3860 74 3872 108
rect 3910 74 3928 108
rect 3928 74 3944 108
rect 4124 74 4158 108
rect 4196 74 4226 108
rect 4226 74 4230 108
rect 4268 74 4294 108
rect 4294 74 4302 108
rect 4340 74 4362 108
rect 4362 74 4374 108
rect 4412 74 4430 108
rect 4430 74 4446 108
rect 4484 74 4498 108
rect 4498 74 4518 108
rect 4556 74 4566 108
rect 4566 74 4590 108
rect 4628 74 4634 108
rect 4634 74 4662 108
rect 4700 74 4702 108
rect 4702 74 4734 108
rect 4772 74 4804 108
rect 4804 74 4806 108
rect 4844 74 4872 108
rect 4872 74 4878 108
rect 4916 74 4940 108
rect 4940 74 4950 108
rect 4988 74 5008 108
rect 5008 74 5022 108
rect 5060 74 5076 108
rect 5076 74 5094 108
rect 5132 74 5144 108
rect 5144 74 5166 108
rect 5204 74 5212 108
rect 5212 74 5238 108
rect 5276 74 5280 108
rect 5280 74 5310 108
rect 5348 74 5382 108
rect 5420 74 5450 108
rect 5450 74 5454 108
rect 5492 74 5518 108
rect 5518 74 5526 108
rect 5564 74 5586 108
rect 5586 74 5598 108
rect 5636 74 5654 108
rect 5654 74 5670 108
rect 5708 74 5722 108
rect 5722 74 5742 108
rect 5780 74 5790 108
rect 5790 74 5814 108
rect 5852 74 5858 108
rect 5858 74 5886 108
rect 5924 74 5926 108
rect 5926 74 5958 108
rect 5996 74 6028 108
rect 6028 74 6030 108
rect 6068 74 6096 108
rect 6096 74 6102 108
rect 6140 74 6164 108
rect 6164 74 6174 108
rect 6212 74 6232 108
rect 6232 74 6246 108
rect 6284 74 6300 108
rect 6300 74 6318 108
rect 6356 74 6368 108
rect 6368 74 6390 108
rect 6428 74 6436 108
rect 6436 74 6462 108
rect 6500 74 6504 108
rect 6504 74 6534 108
rect 6572 74 6606 108
rect 6644 74 6674 108
rect 6674 74 6678 108
rect 6716 74 6742 108
rect 6742 74 6750 108
rect 6788 74 6810 108
rect 6810 74 6822 108
rect 6860 74 6878 108
rect 6878 74 6894 108
rect 6932 74 6946 108
rect 6946 74 6966 108
rect 7004 74 7014 108
rect 7014 74 7038 108
rect 7076 74 7082 108
rect 7082 74 7110 108
rect 7148 74 7150 108
rect 7150 74 7182 108
rect 7220 74 7252 108
rect 7252 74 7254 108
rect 7292 74 7320 108
rect 7320 74 7326 108
rect 7364 74 7388 108
rect 7388 74 7398 108
rect 7436 74 7456 108
rect 7456 74 7470 108
rect 7508 74 7524 108
rect 7524 74 7542 108
rect 7580 74 7592 108
rect 7592 74 7614 108
rect 7652 74 7660 108
rect 7660 74 7686 108
rect 7724 74 7728 108
rect 7728 74 7758 108
rect 7796 74 7830 108
rect 7868 74 7898 108
rect 7898 74 7902 108
rect 7940 74 7966 108
rect 7966 74 7974 108
rect 8012 74 8034 108
rect 8034 74 8046 108
rect 8084 74 8102 108
rect 8102 74 8118 108
rect 8306 74 8318 108
rect 8318 74 8340 108
rect 8378 74 8386 108
rect 8386 74 8412 108
rect 8450 74 8454 108
rect 8454 74 8484 108
rect 8522 74 8556 108
rect 8594 74 8624 108
rect 8624 74 8628 108
rect 8666 74 8692 108
rect 8692 74 8700 108
rect 8738 74 8760 108
rect 8760 74 8772 108
rect 8810 74 8828 108
rect 8828 74 8844 108
rect 8882 74 8896 108
rect 8896 74 8916 108
rect 8954 74 8964 108
rect 8964 74 8988 108
rect 9026 74 9032 108
rect 9032 74 9060 108
rect 9098 74 9100 108
rect 9100 74 9132 108
rect 9170 74 9202 108
rect 9202 74 9204 108
rect 9242 74 9270 108
rect 9270 74 9276 108
rect 9314 74 9338 108
rect 9338 74 9348 108
rect 9386 74 9406 108
rect 9406 74 9420 108
rect 9458 74 9474 108
rect 9474 74 9492 108
rect 9530 74 9542 108
rect 9542 74 9564 108
rect 9602 74 9610 108
rect 9610 74 9636 108
rect 9674 74 9678 108
rect 9678 74 9708 108
rect 9746 74 9780 108
rect 9818 74 9848 108
rect 9848 74 9852 108
rect 9890 74 9916 108
rect 9916 74 9924 108
rect 9962 74 9984 108
rect 9984 74 9996 108
rect 10034 74 10052 108
rect 10052 74 10068 108
rect 10106 74 10120 108
rect 10120 74 10140 108
rect 10178 74 10188 108
rect 10188 74 10212 108
rect 10250 74 10256 108
rect 10256 74 10284 108
rect 10322 74 10324 108
rect 10324 74 10356 108
rect 10394 74 10426 108
rect 10426 74 10428 108
rect 10466 74 10494 108
rect 10494 74 10500 108
rect 10538 74 10562 108
rect 10562 74 10572 108
rect 10610 74 10630 108
rect 10630 74 10644 108
rect 10682 74 10698 108
rect 10698 74 10716 108
rect 10754 74 10766 108
rect 10766 74 10788 108
rect 10826 74 10834 108
rect 10834 74 10860 108
rect 10898 74 10902 108
rect 10902 74 10932 108
rect 10970 74 11004 108
rect 11042 74 11072 108
rect 11072 74 11076 108
rect 11114 74 11140 108
rect 11140 74 11148 108
rect 11186 74 11208 108
rect 11208 74 11220 108
rect 11258 74 11276 108
rect 11276 74 11292 108
rect 14547 155 14581 189
rect 18617 155 18651 189
rect 18691 187 18725 189
rect 18691 155 18719 187
rect 18719 155 18725 187
rect 22794 155 22828 189
rect 22866 187 22900 189
rect 22866 155 22893 187
rect 22893 155 22900 187
rect 11458 74 11474 108
rect 11474 74 11492 108
rect 11530 74 11542 108
rect 11542 74 11564 108
rect 11602 74 11610 108
rect 11610 74 11636 108
rect 11674 74 11678 108
rect 11678 74 11708 108
rect 11746 74 11780 108
rect 11818 74 11848 108
rect 11848 74 11852 108
rect 11890 74 11916 108
rect 11916 74 11924 108
rect 11962 74 11984 108
rect 11984 74 11996 108
rect 12034 74 12052 108
rect 12052 74 12068 108
rect 12106 74 12120 108
rect 12120 74 12140 108
rect 12178 74 12188 108
rect 12188 74 12212 108
rect 12250 74 12256 108
rect 12256 74 12284 108
rect 12322 74 12324 108
rect 12324 74 12356 108
rect 12394 74 12426 108
rect 12426 74 12428 108
rect 12466 74 12494 108
rect 12494 74 12500 108
rect 12538 74 12562 108
rect 12562 74 12572 108
rect 12610 74 12630 108
rect 12630 74 12644 108
rect 12682 74 12698 108
rect 12698 74 12716 108
rect 12754 74 12766 108
rect 12766 74 12788 108
rect 12826 74 12834 108
rect 12834 74 12860 108
rect 12898 74 12902 108
rect 12902 74 12932 108
rect 12970 74 13004 108
rect 13042 74 13072 108
rect 13072 74 13076 108
rect 13114 74 13140 108
rect 13140 74 13148 108
rect 13186 74 13208 108
rect 13208 74 13220 108
rect 13258 74 13276 108
rect 13276 74 13292 108
rect 13330 74 13344 108
rect 13344 74 13364 108
rect 13402 74 13412 108
rect 13412 74 13436 108
rect 13474 74 13480 108
rect 13480 74 13508 108
rect 13546 74 13548 108
rect 13548 74 13580 108
rect 13618 74 13650 108
rect 13650 74 13652 108
rect 13690 74 13718 108
rect 13718 74 13724 108
rect 13762 74 13786 108
rect 13786 74 13796 108
rect 13834 74 13854 108
rect 13854 74 13868 108
rect 13906 74 13922 108
rect 13922 74 13940 108
rect 13978 74 13990 108
rect 13990 74 14012 108
rect 14050 74 14058 108
rect 14058 74 14084 108
rect 14122 74 14126 108
rect 14126 74 14156 108
rect 14194 74 14228 108
rect 14266 74 14296 108
rect 14296 74 14300 108
rect 14338 74 14364 108
rect 14364 74 14372 108
rect 14410 74 14432 108
rect 14432 74 14444 108
rect 14632 74 14648 108
rect 14648 74 14666 108
rect 14704 74 14716 108
rect 14716 74 14738 108
rect 14776 74 14784 108
rect 14784 74 14810 108
rect 14848 74 14852 108
rect 14852 74 14882 108
rect 14920 74 14954 108
rect 14992 74 15022 108
rect 15022 74 15026 108
rect 15064 74 15090 108
rect 15090 74 15098 108
rect 15136 74 15158 108
rect 15158 74 15170 108
rect 15208 74 15226 108
rect 15226 74 15242 108
rect 15280 74 15294 108
rect 15294 74 15314 108
rect 15352 74 15362 108
rect 15362 74 15386 108
rect 15424 74 15430 108
rect 15430 74 15458 108
rect 15496 74 15498 108
rect 15498 74 15530 108
rect 15568 74 15600 108
rect 15600 74 15602 108
rect 15640 74 15668 108
rect 15668 74 15674 108
rect 15712 74 15736 108
rect 15736 74 15746 108
rect 15784 74 15804 108
rect 15804 74 15818 108
rect 15856 74 15872 108
rect 15872 74 15890 108
rect 15928 74 15940 108
rect 15940 74 15962 108
rect 16000 74 16008 108
rect 16008 74 16034 108
rect 16072 74 16076 108
rect 16076 74 16106 108
rect 16144 74 16178 108
rect 16216 74 16246 108
rect 16246 74 16250 108
rect 16288 74 16314 108
rect 16314 74 16322 108
rect 16360 74 16382 108
rect 16382 74 16394 108
rect 16432 74 16450 108
rect 16450 74 16466 108
rect 16504 74 16518 108
rect 16518 74 16538 108
rect 16576 74 16586 108
rect 16586 74 16610 108
rect 16648 74 16654 108
rect 16654 74 16682 108
rect 16720 74 16722 108
rect 16722 74 16754 108
rect 16792 74 16824 108
rect 16824 74 16826 108
rect 16864 74 16892 108
rect 16892 74 16898 108
rect 16936 74 16960 108
rect 16960 74 16970 108
rect 17008 74 17028 108
rect 17028 74 17042 108
rect 17080 74 17096 108
rect 17096 74 17114 108
rect 17152 74 17164 108
rect 17164 74 17186 108
rect 17224 74 17232 108
rect 17232 74 17258 108
rect 17296 74 17300 108
rect 17300 74 17330 108
rect 17368 74 17402 108
rect 17440 74 17470 108
rect 17470 74 17474 108
rect 17512 74 17538 108
rect 17538 74 17546 108
rect 17584 74 17606 108
rect 17606 74 17618 108
rect 17656 74 17674 108
rect 17674 74 17690 108
rect 17728 74 17742 108
rect 17742 74 17762 108
rect 17800 74 17810 108
rect 17810 74 17834 108
rect 17872 74 17878 108
rect 17878 74 17906 108
rect 17944 74 17946 108
rect 17946 74 17978 108
rect 18016 74 18048 108
rect 18048 74 18050 108
rect 18088 74 18116 108
rect 18116 74 18122 108
rect 18160 74 18184 108
rect 18184 74 18194 108
rect 18232 74 18252 108
rect 18252 74 18266 108
rect 18304 74 18320 108
rect 18320 74 18338 108
rect 18376 74 18388 108
rect 18388 74 18410 108
rect 18448 74 18456 108
rect 18456 74 18482 108
rect 18520 74 18524 108
rect 18524 74 18554 108
rect 18592 74 18626 108
rect 18806 74 18822 108
rect 18822 74 18840 108
rect 18878 74 18890 108
rect 18890 74 18912 108
rect 18950 74 18958 108
rect 18958 74 18984 108
rect 19022 74 19026 108
rect 19026 74 19056 108
rect 19094 74 19128 108
rect 19166 74 19196 108
rect 19196 74 19200 108
rect 19238 74 19264 108
rect 19264 74 19272 108
rect 19310 74 19332 108
rect 19332 74 19344 108
rect 19382 74 19400 108
rect 19400 74 19416 108
rect 19454 74 19468 108
rect 19468 74 19488 108
rect 19526 74 19536 108
rect 19536 74 19560 108
rect 19598 74 19604 108
rect 19604 74 19632 108
rect 19670 74 19672 108
rect 19672 74 19704 108
rect 19742 74 19774 108
rect 19774 74 19776 108
rect 19814 74 19842 108
rect 19842 74 19848 108
rect 19886 74 19910 108
rect 19910 74 19920 108
rect 19958 74 19978 108
rect 19978 74 19992 108
rect 20030 74 20046 108
rect 20046 74 20064 108
rect 20102 74 20114 108
rect 20114 74 20136 108
rect 20174 74 20182 108
rect 20182 74 20208 108
rect 20246 74 20250 108
rect 20250 74 20280 108
rect 20318 74 20352 108
rect 20390 74 20420 108
rect 20420 74 20424 108
rect 20462 74 20488 108
rect 20488 74 20496 108
rect 20534 74 20556 108
rect 20556 74 20568 108
rect 20606 74 20624 108
rect 20624 74 20640 108
rect 20678 74 20692 108
rect 20692 74 20712 108
rect 20750 74 20760 108
rect 20760 74 20784 108
rect 20822 74 20828 108
rect 20828 74 20856 108
rect 20894 74 20896 108
rect 20896 74 20928 108
rect 20966 74 20998 108
rect 20998 74 21000 108
rect 21038 74 21066 108
rect 21066 74 21072 108
rect 21110 74 21134 108
rect 21134 74 21144 108
rect 21182 74 21202 108
rect 21202 74 21216 108
rect 21254 74 21270 108
rect 21270 74 21288 108
rect 21326 74 21338 108
rect 21338 74 21360 108
rect 21398 74 21406 108
rect 21406 74 21432 108
rect 21470 74 21474 108
rect 21474 74 21504 108
rect 21542 74 21576 108
rect 21614 74 21644 108
rect 21644 74 21648 108
rect 21686 74 21712 108
rect 21712 74 21720 108
rect 21758 74 21780 108
rect 21780 74 21792 108
rect 21830 74 21848 108
rect 21848 74 21864 108
rect 21902 74 21916 108
rect 21916 74 21936 108
rect 21974 74 21984 108
rect 21984 74 22008 108
rect 22046 74 22052 108
rect 22052 74 22080 108
rect 22118 74 22120 108
rect 22120 74 22152 108
rect 22190 74 22222 108
rect 22222 74 22224 108
rect 22262 74 22290 108
rect 22290 74 22296 108
rect 22334 74 22358 108
rect 22358 74 22368 108
rect 22406 74 22426 108
rect 22426 74 22440 108
rect 22478 74 22494 108
rect 22494 74 22512 108
rect 22550 74 22562 108
rect 22562 74 22584 108
rect 22622 74 22630 108
rect 22630 74 22656 108
rect 22694 74 22698 108
rect 22698 74 22728 108
rect 22766 74 22800 108
<< metal1 >>
rect -73 264 23503 308
rect -73 230 -50 264
rect -16 230 22 264
rect 56 230 94 264
rect 128 230 166 264
rect 200 230 238 264
rect 272 230 310 264
rect 344 230 382 264
rect 416 230 454 264
rect 488 230 526 264
rect 560 230 598 264
rect 632 230 670 264
rect 704 230 742 264
rect 776 230 814 264
rect 848 230 886 264
rect 920 230 958 264
rect 992 230 1030 264
rect 1064 230 1102 264
rect 1136 230 1174 264
rect 1208 230 1246 264
rect 1280 230 1318 264
rect 1352 230 1390 264
rect 1424 230 1462 264
rect 1496 230 1534 264
rect 1568 230 1606 264
rect 1640 230 1678 264
rect 1712 230 1750 264
rect 1784 230 1822 264
rect 1856 230 1894 264
rect 1928 230 1966 264
rect 2000 230 2038 264
rect 2072 230 2110 264
rect 2144 230 2182 264
rect 2216 230 2254 264
rect 2288 230 2326 264
rect 2360 230 2398 264
rect 2432 230 2470 264
rect 2504 230 2542 264
rect 2576 230 2614 264
rect 2648 230 2686 264
rect 2720 230 2758 264
rect 2792 230 2830 264
rect 2864 230 2902 264
rect 2936 230 2974 264
rect 3008 230 3046 264
rect 3080 230 3118 264
rect 3152 230 3190 264
rect 3224 230 3262 264
rect 3296 230 3334 264
rect 3368 230 3406 264
rect 3440 230 3478 264
rect 3512 230 3550 264
rect 3584 230 3622 264
rect 3656 230 3694 264
rect 3728 230 3766 264
rect 3800 230 3838 264
rect 3872 230 3910 264
rect 3944 230 4124 264
rect 4158 230 4196 264
rect 4230 230 4268 264
rect 4302 230 4340 264
rect 4374 230 4412 264
rect 4446 230 4484 264
rect 4518 230 4556 264
rect 4590 230 4628 264
rect 4662 230 4700 264
rect 4734 230 4772 264
rect 4806 230 4844 264
rect 4878 230 4916 264
rect 4950 230 4988 264
rect 5022 230 5060 264
rect 5094 230 5132 264
rect 5166 230 5204 264
rect 5238 230 5276 264
rect 5310 230 5348 264
rect 5382 230 5420 264
rect 5454 230 5492 264
rect 5526 230 5564 264
rect 5598 230 5636 264
rect 5670 230 5708 264
rect 5742 230 5780 264
rect 5814 230 5852 264
rect 5886 230 5924 264
rect 5958 230 5996 264
rect 6030 230 6068 264
rect 6102 230 6140 264
rect 6174 230 6212 264
rect 6246 230 6284 264
rect 6318 230 6356 264
rect 6390 230 6428 264
rect 6462 230 6500 264
rect 6534 230 6572 264
rect 6606 230 6644 264
rect 6678 230 6716 264
rect 6750 230 6788 264
rect 6822 230 6860 264
rect 6894 230 6932 264
rect 6966 230 7004 264
rect 7038 230 7076 264
rect 7110 230 7148 264
rect 7182 230 7220 264
rect 7254 230 7292 264
rect 7326 230 7364 264
rect 7398 230 7436 264
rect 7470 230 7508 264
rect 7542 230 7580 264
rect 7614 230 7652 264
rect 7686 230 7724 264
rect 7758 230 7796 264
rect 7830 230 7868 264
rect 7902 230 7940 264
rect 7974 230 8012 264
rect 8046 230 8084 264
rect 8118 230 8306 264
rect 8340 230 8378 264
rect 8412 230 8450 264
rect 8484 230 8522 264
rect 8556 230 8594 264
rect 8628 230 8666 264
rect 8700 230 8738 264
rect 8772 230 8810 264
rect 8844 230 8882 264
rect 8916 230 8954 264
rect 8988 230 9026 264
rect 9060 230 9098 264
rect 9132 230 9170 264
rect 9204 230 9242 264
rect 9276 230 9314 264
rect 9348 230 9386 264
rect 9420 230 9458 264
rect 9492 230 9530 264
rect 9564 230 9602 264
rect 9636 230 9674 264
rect 9708 230 9746 264
rect 9780 230 9818 264
rect 9852 230 9890 264
rect 9924 230 9962 264
rect 9996 230 10034 264
rect 10068 230 10106 264
rect 10140 230 10178 264
rect 10212 230 10250 264
rect 10284 230 10322 264
rect 10356 230 10394 264
rect 10428 230 10466 264
rect 10500 230 10538 264
rect 10572 230 10610 264
rect 10644 230 10682 264
rect 10716 230 10754 264
rect 10788 230 10826 264
rect 10860 230 10898 264
rect 10932 230 10970 264
rect 11004 230 11042 264
rect 11076 230 11114 264
rect 11148 230 11186 264
rect 11220 230 11258 264
rect 11292 230 11458 264
rect 11492 230 11530 264
rect 11564 230 11602 264
rect 11636 230 11674 264
rect 11708 230 11746 264
rect 11780 230 11818 264
rect 11852 230 11890 264
rect 11924 230 11962 264
rect 11996 230 12034 264
rect 12068 230 12106 264
rect 12140 230 12178 264
rect 12212 230 12250 264
rect 12284 230 12322 264
rect 12356 230 12394 264
rect 12428 230 12466 264
rect 12500 230 12538 264
rect 12572 230 12610 264
rect 12644 230 12682 264
rect 12716 230 12754 264
rect 12788 230 12826 264
rect 12860 230 12898 264
rect 12932 230 12970 264
rect 13004 230 13042 264
rect 13076 230 13114 264
rect 13148 230 13186 264
rect 13220 230 13258 264
rect 13292 230 13330 264
rect 13364 230 13402 264
rect 13436 230 13474 264
rect 13508 230 13546 264
rect 13580 230 13618 264
rect 13652 230 13690 264
rect 13724 230 13762 264
rect 13796 230 13834 264
rect 13868 230 13906 264
rect 13940 230 13978 264
rect 14012 230 14050 264
rect 14084 230 14122 264
rect 14156 230 14194 264
rect 14228 230 14266 264
rect 14300 230 14338 264
rect 14372 230 14410 264
rect 14444 230 14632 264
rect 14666 230 14704 264
rect 14738 230 14776 264
rect 14810 230 14848 264
rect 14882 230 14920 264
rect 14954 230 14992 264
rect 15026 230 15064 264
rect 15098 230 15136 264
rect 15170 230 15208 264
rect 15242 230 15280 264
rect 15314 230 15352 264
rect 15386 230 15424 264
rect 15458 230 15496 264
rect 15530 230 15568 264
rect 15602 230 15640 264
rect 15674 230 15712 264
rect 15746 230 15784 264
rect 15818 230 15856 264
rect 15890 230 15928 264
rect 15962 230 16000 264
rect 16034 230 16072 264
rect 16106 230 16144 264
rect 16178 230 16216 264
rect 16250 230 16288 264
rect 16322 230 16360 264
rect 16394 230 16432 264
rect 16466 230 16504 264
rect 16538 230 16576 264
rect 16610 230 16648 264
rect 16682 230 16720 264
rect 16754 230 16792 264
rect 16826 230 16864 264
rect 16898 230 16936 264
rect 16970 230 17008 264
rect 17042 230 17080 264
rect 17114 230 17152 264
rect 17186 230 17224 264
rect 17258 230 17296 264
rect 17330 230 17368 264
rect 17402 230 17440 264
rect 17474 230 17512 264
rect 17546 230 17584 264
rect 17618 230 17656 264
rect 17690 230 17728 264
rect 17762 230 17800 264
rect 17834 230 17872 264
rect 17906 230 17944 264
rect 17978 230 18016 264
rect 18050 230 18088 264
rect 18122 230 18160 264
rect 18194 230 18232 264
rect 18266 230 18304 264
rect 18338 230 18376 264
rect 18410 230 18448 264
rect 18482 230 18520 264
rect 18554 230 18592 264
rect 18626 230 18806 264
rect 18840 230 18878 264
rect 18912 230 18950 264
rect 18984 230 19022 264
rect 19056 230 19094 264
rect 19128 230 19166 264
rect 19200 230 19238 264
rect 19272 230 19310 264
rect 19344 230 19382 264
rect 19416 230 19454 264
rect 19488 230 19526 264
rect 19560 230 19598 264
rect 19632 230 19670 264
rect 19704 230 19742 264
rect 19776 230 19814 264
rect 19848 230 19886 264
rect 19920 230 19958 264
rect 19992 230 20030 264
rect 20064 230 20102 264
rect 20136 230 20174 264
rect 20208 230 20246 264
rect 20280 230 20318 264
rect 20352 230 20390 264
rect 20424 230 20462 264
rect 20496 230 20534 264
rect 20568 230 20606 264
rect 20640 230 20678 264
rect 20712 230 20750 264
rect 20784 230 20822 264
rect 20856 230 20894 264
rect 20928 230 20966 264
rect 21000 230 21038 264
rect 21072 230 21110 264
rect 21144 230 21182 264
rect 21216 230 21254 264
rect 21288 230 21326 264
rect 21360 230 21398 264
rect 21432 230 21470 264
rect 21504 230 21542 264
rect 21576 230 21614 264
rect 21648 230 21686 264
rect 21720 230 21758 264
rect 21792 230 21830 264
rect 21864 230 21902 264
rect 21936 230 21974 264
rect 22008 230 22046 264
rect 22080 230 22118 264
rect 22152 230 22190 264
rect 22224 230 22262 264
rect 22296 230 22334 264
rect 22368 230 22406 264
rect 22440 230 22478 264
rect 22512 230 22550 264
rect 22584 230 22622 264
rect 22656 230 22694 264
rect 22728 230 22766 264
rect 22800 230 23503 264
rect -73 224 23503 230
rect -79 149 3806 195
rect 3807 150 3808 194
rect 3868 150 3869 194
rect 3870 189 4240 195
rect 4242 194 4302 195
rect 3870 155 3982 189
rect 4016 155 4054 189
rect 4088 155 4240 189
rect 3870 149 4240 155
rect 4241 150 4303 194
rect 4304 189 8404 195
rect 8406 194 8466 195
rect 4304 155 8156 189
rect 8190 155 8228 189
rect 8262 155 8404 189
rect 4242 149 4302 150
rect 4304 149 8404 155
rect 8405 150 8467 194
rect 8468 189 11544 195
rect 11546 194 11606 195
rect 8468 155 11330 189
rect 11364 155 11402 189
rect 11436 155 11544 189
rect 8406 149 8466 150
rect 8468 149 11544 155
rect 11545 150 11607 194
rect 11608 189 14687 195
rect 14689 194 14749 195
rect 11608 155 14475 189
rect 14509 155 14547 189
rect 14581 155 14687 189
rect 11546 149 11606 150
rect 11608 149 14687 155
rect 14688 150 14750 194
rect 14751 189 18789 195
rect 18791 194 18851 195
rect 14751 155 18617 189
rect 18651 155 18691 189
rect 18725 155 18789 189
rect 14689 149 14749 150
rect 14751 149 18789 155
rect 18790 150 18852 194
rect 18853 189 22928 195
rect 22930 194 22990 195
rect 18853 155 22794 189
rect 22828 155 22866 189
rect 22900 155 22928 189
rect 18791 149 18851 150
rect 18853 149 22928 155
rect 22929 150 22991 194
rect 22930 149 22990 150
rect 22992 149 23044 195
rect -62 108 4000 114
rect 4002 113 4062 114
rect -62 74 -50 108
rect -16 74 22 108
rect 56 74 94 108
rect 128 74 166 108
rect 200 74 238 108
rect 272 74 310 108
rect 344 74 382 108
rect 416 74 454 108
rect 488 74 526 108
rect 560 74 598 108
rect 632 74 670 108
rect 704 74 742 108
rect 776 74 814 108
rect 848 74 886 108
rect 920 74 958 108
rect 992 74 1030 108
rect 1064 74 1102 108
rect 1136 74 1174 108
rect 1208 74 1246 108
rect 1280 74 1318 108
rect 1352 74 1390 108
rect 1424 74 1462 108
rect 1496 74 1534 108
rect 1568 74 1606 108
rect 1640 74 1678 108
rect 1712 74 1750 108
rect 1784 74 1822 108
rect 1856 74 1894 108
rect 1928 74 1966 108
rect 2000 74 2038 108
rect 2072 74 2110 108
rect 2144 74 2182 108
rect 2216 74 2254 108
rect 2288 74 2326 108
rect 2360 74 2398 108
rect 2432 74 2470 108
rect 2504 74 2542 108
rect 2576 74 2614 108
rect 2648 74 2686 108
rect 2720 74 2758 108
rect 2792 74 2830 108
rect 2864 74 2902 108
rect 2936 74 2974 108
rect 3008 74 3046 108
rect 3080 74 3118 108
rect 3152 74 3190 108
rect 3224 74 3262 108
rect 3296 74 3334 108
rect 3368 74 3406 108
rect 3440 74 3478 108
rect 3512 74 3550 108
rect 3584 74 3622 108
rect 3656 74 3694 108
rect 3728 74 3766 108
rect 3800 74 3838 108
rect 3872 74 3910 108
rect 3944 74 4000 108
rect -62 68 4000 74
rect 4001 69 4063 113
rect 4064 108 8179 114
rect 8181 113 8241 114
rect 4064 74 4124 108
rect 4158 74 4196 108
rect 4230 74 4268 108
rect 4302 74 4340 108
rect 4374 74 4412 108
rect 4446 74 4484 108
rect 4518 74 4556 108
rect 4590 74 4628 108
rect 4662 74 4700 108
rect 4734 74 4772 108
rect 4806 74 4844 108
rect 4878 74 4916 108
rect 4950 74 4988 108
rect 5022 74 5060 108
rect 5094 74 5132 108
rect 5166 74 5204 108
rect 5238 74 5276 108
rect 5310 74 5348 108
rect 5382 74 5420 108
rect 5454 74 5492 108
rect 5526 74 5564 108
rect 5598 74 5636 108
rect 5670 74 5708 108
rect 5742 74 5780 108
rect 5814 74 5852 108
rect 5886 74 5924 108
rect 5958 74 5996 108
rect 6030 74 6068 108
rect 6102 74 6140 108
rect 6174 74 6212 108
rect 6246 74 6284 108
rect 6318 74 6356 108
rect 6390 74 6428 108
rect 6462 74 6500 108
rect 6534 74 6572 108
rect 6606 74 6644 108
rect 6678 74 6716 108
rect 6750 74 6788 108
rect 6822 74 6860 108
rect 6894 74 6932 108
rect 6966 74 7004 108
rect 7038 74 7076 108
rect 7110 74 7148 108
rect 7182 74 7220 108
rect 7254 74 7292 108
rect 7326 74 7364 108
rect 7398 74 7436 108
rect 7470 74 7508 108
rect 7542 74 7580 108
rect 7614 74 7652 108
rect 7686 74 7724 108
rect 7758 74 7796 108
rect 7830 74 7868 108
rect 7902 74 7940 108
rect 7974 74 8012 108
rect 8046 74 8084 108
rect 8118 74 8179 108
rect 4002 68 4062 69
rect 4064 68 8179 74
rect 8180 69 8242 113
rect 8243 108 11304 114
tri 11435 108 11441 114 se
rect 11441 108 14504 114
rect 14506 113 14566 114
rect 8243 74 8306 108
rect 8340 74 8378 108
rect 8412 74 8450 108
rect 8484 74 8522 108
rect 8556 74 8594 108
rect 8628 74 8666 108
rect 8700 74 8738 108
rect 8772 74 8810 108
rect 8844 74 8882 108
rect 8916 74 8954 108
rect 8988 74 9026 108
rect 9060 74 9098 108
rect 9132 74 9170 108
rect 9204 74 9242 108
rect 9276 74 9314 108
rect 9348 74 9386 108
rect 9420 74 9458 108
rect 9492 74 9530 108
rect 9564 74 9602 108
rect 9636 74 9674 108
rect 9708 74 9746 108
rect 9780 74 9818 108
rect 9852 74 9890 108
rect 9924 74 9962 108
rect 9996 74 10034 108
rect 10068 74 10106 108
rect 10140 74 10178 108
rect 10212 74 10250 108
rect 10284 74 10322 108
rect 10356 74 10394 108
rect 10428 74 10466 108
rect 10500 74 10538 108
rect 10572 74 10610 108
rect 10644 74 10682 108
rect 10716 74 10754 108
rect 10788 74 10826 108
rect 10860 74 10898 108
rect 10932 74 10970 108
rect 11004 74 11042 108
rect 11076 74 11114 108
rect 11148 74 11186 108
rect 11220 74 11258 108
rect 11292 74 11304 108
tri 11401 74 11435 108 se
rect 11435 74 11458 108
rect 11492 74 11530 108
rect 11564 74 11602 108
rect 11636 74 11674 108
rect 11708 74 11746 108
rect 11780 74 11818 108
rect 11852 74 11890 108
rect 11924 74 11962 108
rect 11996 74 12034 108
rect 12068 74 12106 108
rect 12140 74 12178 108
rect 12212 74 12250 108
rect 12284 74 12322 108
rect 12356 74 12394 108
rect 12428 74 12466 108
rect 12500 74 12538 108
rect 12572 74 12610 108
rect 12644 74 12682 108
rect 12716 74 12754 108
rect 12788 74 12826 108
rect 12860 74 12898 108
rect 12932 74 12970 108
rect 13004 74 13042 108
rect 13076 74 13114 108
rect 13148 74 13186 108
rect 13220 74 13258 108
rect 13292 74 13330 108
rect 13364 74 13402 108
rect 13436 74 13474 108
rect 13508 74 13546 108
rect 13580 74 13618 108
rect 13652 74 13690 108
rect 13724 74 13762 108
rect 13796 74 13834 108
rect 13868 74 13906 108
rect 13940 74 13978 108
rect 14012 74 14050 108
rect 14084 74 14122 108
rect 14156 74 14194 108
rect 14228 74 14266 108
rect 14300 74 14338 108
rect 14372 74 14410 108
rect 14444 74 14504 108
rect 8181 68 8241 69
rect 8243 68 11304 74
tri 11395 68 11401 74 se
rect 11401 68 14504 74
rect 14505 69 14567 113
rect 14568 108 18678 114
rect 18680 113 18740 114
rect 14568 74 14632 108
rect 14666 74 14704 108
rect 14738 74 14776 108
rect 14810 74 14848 108
rect 14882 74 14920 108
rect 14954 74 14992 108
rect 15026 74 15064 108
rect 15098 74 15136 108
rect 15170 74 15208 108
rect 15242 74 15280 108
rect 15314 74 15352 108
rect 15386 74 15424 108
rect 15458 74 15496 108
rect 15530 74 15568 108
rect 15602 74 15640 108
rect 15674 74 15712 108
rect 15746 74 15784 108
rect 15818 74 15856 108
rect 15890 74 15928 108
rect 15962 74 16000 108
rect 16034 74 16072 108
rect 16106 74 16144 108
rect 16178 74 16216 108
rect 16250 74 16288 108
rect 16322 74 16360 108
rect 16394 74 16432 108
rect 16466 74 16504 108
rect 16538 74 16576 108
rect 16610 74 16648 108
rect 16682 74 16720 108
rect 16754 74 16792 108
rect 16826 74 16864 108
rect 16898 74 16936 108
rect 16970 74 17008 108
rect 17042 74 17080 108
rect 17114 74 17152 108
rect 17186 74 17224 108
rect 17258 74 17296 108
rect 17330 74 17368 108
rect 17402 74 17440 108
rect 17474 74 17512 108
rect 17546 74 17584 108
rect 17618 74 17656 108
rect 17690 74 17728 108
rect 17762 74 17800 108
rect 17834 74 17872 108
rect 17906 74 17944 108
rect 17978 74 18016 108
rect 18050 74 18088 108
rect 18122 74 18160 108
rect 18194 74 18232 108
rect 18266 74 18304 108
rect 18338 74 18376 108
rect 18410 74 18448 108
rect 18482 74 18520 108
rect 18554 74 18592 108
rect 18626 74 18678 108
rect 14506 68 14566 69
rect 14568 68 18678 74
rect 18679 69 18741 113
rect 18742 108 22812 114
rect 18742 74 18806 108
rect 18840 74 18878 108
rect 18912 74 18950 108
rect 18984 74 19022 108
rect 19056 74 19094 108
rect 19128 74 19166 108
rect 19200 74 19238 108
rect 19272 74 19310 108
rect 19344 74 19382 108
rect 19416 74 19454 108
rect 19488 74 19526 108
rect 19560 74 19598 108
rect 19632 74 19670 108
rect 19704 74 19742 108
rect 19776 74 19814 108
rect 19848 74 19886 108
rect 19920 74 19958 108
rect 19992 74 20030 108
rect 20064 74 20102 108
rect 20136 74 20174 108
rect 20208 74 20246 108
rect 20280 74 20318 108
rect 20352 74 20390 108
rect 20424 74 20462 108
rect 20496 74 20534 108
rect 20568 74 20606 108
rect 20640 74 20678 108
rect 20712 74 20750 108
rect 20784 74 20822 108
rect 20856 74 20894 108
rect 20928 74 20966 108
rect 21000 74 21038 108
rect 21072 74 21110 108
rect 21144 74 21182 108
rect 21216 74 21254 108
rect 21288 74 21326 108
rect 21360 74 21398 108
rect 21432 74 21470 108
rect 21504 74 21542 108
rect 21576 74 21614 108
rect 21648 74 21686 108
rect 21720 74 21758 108
rect 21792 74 21830 108
rect 21864 74 21902 108
rect 21936 74 21974 108
rect 22008 74 22046 108
rect 22080 74 22118 108
rect 22152 74 22190 108
rect 22224 74 22262 108
rect 22296 74 22334 108
rect 22368 74 22406 108
rect 22440 74 22478 108
rect 22512 74 22550 108
rect 22584 74 22622 108
rect 22656 74 22694 108
rect 22728 74 22766 108
rect 22800 74 22812 108
rect 18680 68 18740 69
rect 18742 68 22812 74
tri 11389 62 11395 68 se
rect 11395 62 11441 68
tri 11441 62 11447 68 nw
tri 11363 36 11389 62 se
rect 11389 36 11415 62
tri 11415 36 11441 62 nw
rect 332 4 11383 36
tri 11383 4 11415 36 nw
<< rmetal1 >>
rect 3806 194 3808 195
rect 3806 150 3807 194
rect 3806 149 3808 150
rect 3868 194 3870 195
rect 3869 150 3870 194
rect 4240 194 4242 195
rect 4302 194 4304 195
rect 3868 149 3870 150
rect 4240 150 4241 194
rect 4303 150 4304 194
rect 8404 194 8406 195
rect 8466 194 8468 195
rect 4240 149 4242 150
rect 4302 149 4304 150
rect 8404 150 8405 194
rect 8467 150 8468 194
rect 11544 194 11546 195
rect 11606 194 11608 195
rect 8404 149 8406 150
rect 8466 149 8468 150
rect 11544 150 11545 194
rect 11607 150 11608 194
rect 14687 194 14689 195
rect 14749 194 14751 195
rect 11544 149 11546 150
rect 11606 149 11608 150
rect 14687 150 14688 194
rect 14750 150 14751 194
rect 18789 194 18791 195
rect 18851 194 18853 195
rect 14687 149 14689 150
rect 14749 149 14751 150
rect 18789 150 18790 194
rect 18852 150 18853 194
rect 22928 194 22930 195
rect 22990 194 22992 195
rect 18789 149 18791 150
rect 18851 149 18853 150
rect 22928 150 22929 194
rect 22991 150 22992 194
rect 22928 149 22930 150
rect 22990 149 22992 150
rect 4000 113 4002 114
rect 4062 113 4064 114
rect 4000 69 4001 113
rect 4063 69 4064 113
rect 8179 113 8181 114
rect 8241 113 8243 114
rect 4000 68 4002 69
rect 4062 68 4064 69
rect 8179 69 8180 113
rect 8242 69 8243 113
rect 14504 113 14506 114
rect 14566 113 14568 114
rect 8179 68 8181 69
rect 8241 68 8243 69
rect 14504 69 14505 113
rect 14567 69 14568 113
rect 18678 113 18680 114
rect 18740 113 18742 114
rect 14504 68 14506 69
rect 14566 68 14568 69
rect 18678 69 18679 113
rect 18741 69 18742 113
rect 18678 68 18680 69
rect 18740 68 18742 69
use sky130_fd_io__tk_em1o_cdns_5595914180840  sky130_fd_io__tk_em1o_cdns_5595914180840_0
timestamp 1666199351
transform 1 0 3754 0 -1 195
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_55959141808161  sky130_fd_io__tk_em1s_cdns_55959141808161_0
timestamp 1666199351
transform 1 0 3948 0 -1 114
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_55959141808161  sky130_fd_io__tk_em1s_cdns_55959141808161_1
timestamp 1666199351
transform 1 0 8127 0 -1 114
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_55959141808161  sky130_fd_io__tk_em1s_cdns_55959141808161_2
timestamp 1666199351
transform 1 0 4188 0 -1 195
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_55959141808161  sky130_fd_io__tk_em1s_cdns_55959141808161_3
timestamp 1666199351
transform 1 0 8352 0 -1 195
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_55959141808161  sky130_fd_io__tk_em1s_cdns_55959141808161_4
timestamp 1666199351
transform 1 0 11492 0 -1 195
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_55959141808161  sky130_fd_io__tk_em1s_cdns_55959141808161_5
timestamp 1666199351
transform 1 0 14635 0 -1 195
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_55959141808161  sky130_fd_io__tk_em1s_cdns_55959141808161_6
timestamp 1666199351
transform 1 0 18737 0 -1 195
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_55959141808161  sky130_fd_io__tk_em1s_cdns_55959141808161_7
timestamp 1666199351
transform 1 0 22876 0 -1 195
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_55959141808161  sky130_fd_io__tk_em1s_cdns_55959141808161_8
timestamp 1666199351
transform -1 0 18794 0 -1 114
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_55959141808161  sky130_fd_io__tk_em1s_cdns_55959141808161_9
timestamp 1666199351
transform -1 0 14620 0 -1 114
box 0 0 1 1
use sky130_fd_pr__pfet_01v8__example_55959141808162  sky130_fd_pr__pfet_01v8__example_55959141808162_0
timestamp 1666199351
transform 0 1 11462 1 0 119
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808162  sky130_fd_pr__pfet_01v8__example_55959141808162_1
timestamp 1666199351
transform 0 -1 11288 1 0 119
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808164  sky130_fd_pr__pfet_01v8__example_55959141808164_0
timestamp 1666199351
transform 0 1 14636 1 0 119
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808164  sky130_fd_pr__pfet_01v8__example_55959141808164_1
timestamp 1666199351
transform 0 1 14636 1 0 119
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808164  sky130_fd_pr__pfet_01v8__example_55959141808164_2
timestamp 1666199351
transform 0 1 18810 1 0 119
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808164  sky130_fd_pr__pfet_01v8__example_55959141808164_3
timestamp 1666199351
transform 0 -1 8114 1 0 119
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808164  sky130_fd_pr__pfet_01v8__example_55959141808164_4
timestamp 1666199351
transform 0 -1 3940 1 0 119
box -1 0 101 1
<< labels >>
flabel comment s 639 21 639 21 0 FreeSans 200 0 0 0 PGHS_H_LATCH
flabel comment s 381 98 381 98 0 FreeSans 200 0 0 0 PGHS_H
<< properties >>
string GDS_END 34172612
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 34164850
<< end >>
