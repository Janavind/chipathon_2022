magic
tech sky130B
magscale 1 2
timestamp 1666199351
<< nwell >>
rect -38 261 1326 582
<< pwell >>
rect 834 157 1287 203
rect 1 21 1287 157
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 351 47 381 131
rect 435 47 465 131
rect 543 47 573 119
rect 629 47 659 119
rect 724 47 754 131
rect 912 47 942 177
rect 996 47 1026 177
rect 1179 47 1209 177
<< scpmoshvt >>
rect 79 363 109 491
rect 163 363 193 491
rect 351 369 381 497
rect 435 369 465 497
rect 531 413 561 497
rect 652 413 682 497
rect 724 413 754 497
rect 912 297 942 497
rect 996 297 1026 497
rect 1179 297 1209 497
<< ndiff >>
rect 27 119 79 131
rect 27 85 35 119
rect 69 85 79 119
rect 27 47 79 85
rect 109 93 163 131
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 119 245 131
rect 193 85 203 119
rect 237 85 245 119
rect 193 47 245 85
rect 299 119 351 131
rect 299 85 307 119
rect 341 85 351 119
rect 299 47 351 85
rect 381 89 435 131
rect 381 55 391 89
rect 425 55 435 89
rect 381 47 435 55
rect 465 119 515 131
rect 860 165 912 177
rect 860 131 868 165
rect 902 131 912 165
rect 674 119 724 131
rect 465 47 543 119
rect 573 107 629 119
rect 573 73 584 107
rect 618 73 629 107
rect 573 47 629 73
rect 659 47 724 119
rect 754 106 806 131
rect 754 72 764 106
rect 798 72 806 106
rect 754 47 806 72
rect 860 97 912 131
rect 860 63 868 97
rect 902 63 912 97
rect 860 47 912 63
rect 942 47 996 177
rect 1026 93 1179 177
rect 1026 59 1053 93
rect 1087 59 1134 93
rect 1168 59 1179 93
rect 1026 47 1179 59
rect 1209 133 1261 177
rect 1209 99 1219 133
rect 1253 99 1261 133
rect 1209 47 1261 99
<< pdiff >>
rect 27 477 79 491
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 363 79 375
rect 109 461 163 491
rect 109 427 119 461
rect 153 427 163 461
rect 109 363 163 427
rect 193 477 245 491
rect 193 443 203 477
rect 237 443 245 477
rect 193 409 245 443
rect 193 375 203 409
rect 237 375 245 409
rect 193 363 245 375
rect 299 483 351 497
rect 299 449 307 483
rect 341 449 351 483
rect 299 415 351 449
rect 299 381 307 415
rect 341 381 351 415
rect 299 369 351 381
rect 381 485 435 497
rect 381 451 391 485
rect 425 451 435 485
rect 381 417 435 451
rect 381 383 391 417
rect 425 383 435 417
rect 381 369 435 383
rect 465 413 531 497
rect 561 485 652 497
rect 561 451 596 485
rect 630 451 652 485
rect 561 413 652 451
rect 682 413 724 497
rect 754 477 806 497
rect 754 443 764 477
rect 798 443 806 477
rect 754 413 806 443
rect 860 485 912 497
rect 860 451 868 485
rect 902 451 912 485
rect 465 369 515 413
rect 860 297 912 451
rect 942 471 996 497
rect 942 437 952 471
rect 986 437 996 471
rect 942 368 996 437
rect 942 334 952 368
rect 986 334 996 368
rect 942 297 996 334
rect 1026 485 1179 497
rect 1026 451 1053 485
rect 1087 451 1135 485
rect 1169 451 1179 485
rect 1026 297 1179 451
rect 1209 475 1261 497
rect 1209 441 1219 475
rect 1253 441 1261 475
rect 1209 384 1261 441
rect 1209 350 1219 384
rect 1253 350 1261 384
rect 1209 297 1261 350
<< ndiffc >>
rect 35 85 69 119
rect 119 59 153 93
rect 203 85 237 119
rect 307 85 341 119
rect 391 55 425 89
rect 868 131 902 165
rect 584 73 618 107
rect 764 72 798 106
rect 868 63 902 97
rect 1053 59 1087 93
rect 1134 59 1168 93
rect 1219 99 1253 133
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 119 427 153 461
rect 203 443 237 477
rect 203 375 237 409
rect 307 449 341 483
rect 307 381 341 415
rect 391 451 425 485
rect 391 383 425 417
rect 596 451 630 485
rect 764 443 798 477
rect 868 451 902 485
rect 952 437 986 471
rect 952 334 986 368
rect 1053 451 1087 485
rect 1135 451 1169 485
rect 1219 441 1253 475
rect 1219 350 1253 384
<< poly >>
rect 79 491 109 517
rect 163 491 193 517
rect 351 497 381 523
rect 435 497 465 523
rect 531 497 561 523
rect 652 497 682 523
rect 724 497 754 523
rect 912 497 942 523
rect 996 497 1026 523
rect 1179 497 1209 523
rect 79 348 109 363
rect 46 318 109 348
rect 46 280 76 318
rect 21 264 76 280
rect 163 274 193 363
rect 21 230 32 264
rect 66 230 76 264
rect 21 214 76 230
rect 118 264 193 274
rect 118 230 134 264
rect 168 230 193 264
rect 351 241 381 369
rect 118 220 193 230
rect 46 176 76 214
rect 46 146 109 176
rect 79 131 109 146
rect 163 131 193 220
rect 298 225 381 241
rect 298 191 308 225
rect 342 191 381 225
rect 435 219 465 369
rect 531 337 561 413
rect 652 375 682 413
rect 507 321 561 337
rect 603 365 682 375
rect 603 331 619 365
rect 653 331 682 365
rect 603 321 682 331
rect 724 373 754 413
rect 724 357 812 373
rect 724 323 768 357
rect 802 323 812 357
rect 507 287 517 321
rect 551 287 561 321
rect 507 279 561 287
rect 724 307 812 323
rect 507 271 659 279
rect 531 249 659 271
rect 298 175 381 191
rect 351 131 381 175
rect 424 203 478 219
rect 424 169 434 203
rect 468 169 478 203
rect 424 153 478 169
rect 533 191 587 207
rect 533 157 543 191
rect 577 157 587 191
rect 435 131 465 153
rect 533 141 587 157
rect 543 119 573 141
rect 629 119 659 249
rect 724 131 754 307
rect 912 259 942 297
rect 996 265 1026 297
rect 1179 265 1209 297
rect 796 249 942 259
rect 796 215 812 249
rect 846 215 942 249
rect 796 205 942 215
rect 912 177 942 205
rect 986 249 1040 265
rect 986 215 996 249
rect 1030 215 1040 249
rect 986 199 1040 215
rect 1141 249 1209 265
rect 1141 215 1151 249
rect 1185 215 1209 249
rect 1141 199 1209 215
rect 996 177 1026 199
rect 1179 177 1209 199
rect 79 21 109 47
rect 163 21 193 47
rect 351 21 381 47
rect 435 21 465 47
rect 543 21 573 47
rect 629 21 659 47
rect 724 21 754 47
rect 912 21 942 47
rect 996 21 1026 47
rect 1179 21 1209 47
<< polycont >>
rect 32 230 66 264
rect 134 230 168 264
rect 308 191 342 225
rect 619 331 653 365
rect 768 323 802 357
rect 517 287 551 321
rect 434 169 468 203
rect 543 157 577 191
rect 812 215 846 249
rect 996 215 1030 249
rect 1151 215 1185 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 35 477 69 493
rect 35 409 69 443
rect 103 461 169 527
rect 103 427 119 461
rect 153 427 169 461
rect 203 477 248 493
rect 391 485 454 527
rect 237 443 248 477
rect 203 409 248 443
rect 69 375 156 393
rect 35 359 156 375
rect 17 264 66 325
rect 17 230 32 264
rect 17 197 66 230
rect 122 323 156 359
rect 122 280 156 289
rect 237 391 248 409
rect 203 357 214 375
rect 203 337 248 357
rect 291 449 307 483
rect 341 449 357 483
rect 291 415 357 449
rect 291 381 307 415
rect 341 381 357 415
rect 122 264 168 280
rect 122 230 134 264
rect 122 214 168 230
rect 122 161 156 214
rect 35 127 156 161
rect 35 119 69 127
rect 203 119 237 337
rect 291 333 357 381
rect 425 451 454 485
rect 580 451 596 485
rect 630 451 730 485
rect 391 417 454 451
rect 425 383 454 417
rect 391 367 454 383
rect 494 391 551 401
rect 528 357 551 391
rect 291 299 428 333
rect 292 225 358 265
rect 292 191 308 225
rect 342 191 358 225
rect 394 219 428 299
rect 494 321 551 357
rect 494 287 517 321
rect 494 271 551 287
rect 585 365 653 399
rect 585 331 619 365
rect 585 323 653 331
rect 585 289 586 323
rect 620 289 653 323
rect 585 283 653 289
rect 394 203 468 219
rect 585 207 619 283
rect 696 265 730 451
rect 764 477 822 527
rect 798 443 822 477
rect 764 427 822 443
rect 860 485 916 527
rect 860 451 868 485
rect 902 451 916 485
rect 860 427 916 451
rect 950 471 988 493
rect 950 437 952 471
rect 986 437 988 471
rect 950 373 988 437
rect 1022 485 1185 527
rect 1022 451 1053 485
rect 1087 451 1135 485
rect 1169 451 1185 485
rect 1022 427 1185 451
rect 1219 475 1271 491
rect 1253 441 1271 475
rect 1219 384 1271 441
rect 764 368 1185 373
rect 764 357 952 368
rect 764 323 768 357
rect 802 334 952 357
rect 986 334 1185 368
rect 802 323 1185 334
rect 764 307 1185 323
rect 696 249 866 265
rect 394 169 434 203
rect 394 157 468 169
rect 35 69 69 85
rect 103 59 119 93
rect 153 59 169 93
rect 203 69 237 85
rect 307 153 468 157
rect 543 191 619 207
rect 577 157 619 191
rect 307 123 428 153
rect 543 141 619 157
rect 666 215 812 249
rect 846 215 866 249
rect 666 205 866 215
rect 900 249 1087 265
rect 900 215 996 249
rect 1030 215 1087 249
rect 307 119 341 123
rect 666 107 700 205
rect 900 199 1087 215
rect 1121 249 1185 307
rect 1121 215 1151 249
rect 1121 165 1185 215
rect 307 69 341 85
rect 103 17 169 59
rect 375 55 391 89
rect 425 55 441 89
rect 568 73 584 107
rect 618 73 700 107
rect 848 131 868 165
rect 902 131 1185 165
rect 1253 350 1271 384
rect 1219 133 1271 350
rect 375 17 441 55
rect 748 72 764 106
rect 798 72 814 106
rect 748 17 814 72
rect 848 97 918 131
rect 1253 99 1271 133
rect 848 63 868 97
rect 902 63 918 97
rect 848 51 918 63
rect 1019 93 1185 97
rect 1019 59 1053 93
rect 1087 59 1134 93
rect 1168 59 1185 93
rect 1219 83 1271 99
rect 1019 17 1185 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 122 289 156 323
rect 214 375 237 391
rect 237 375 248 391
rect 214 357 248 375
rect 494 357 528 391
rect 586 289 620 323
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
<< metal1 >>
rect 0 561 1288 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 0 496 1288 527
rect 202 391 260 397
rect 202 357 214 391
rect 248 388 260 391
rect 482 391 540 397
rect 482 388 494 391
rect 248 360 494 388
rect 248 357 260 360
rect 202 351 260 357
rect 482 357 494 360
rect 528 357 540 391
rect 482 351 540 357
rect 110 323 168 329
rect 110 289 122 323
rect 156 320 168 323
rect 574 323 632 329
rect 574 320 586 323
rect 156 292 586 320
rect 156 289 168 292
rect 110 283 168 289
rect 574 289 586 292
rect 620 289 632 323
rect 574 283 632 289
rect 0 17 1288 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
rect 0 -48 1288 -17
<< labels >>
flabel locali s 958 221 992 255 0 FreeSans 200 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1050 221 1084 255 0 FreeSans 200 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1230 153 1264 187 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 1230 221 1264 255 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 310 221 344 255 0 FreeSans 200 0 0 0 D
port 1 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 GATE_N
port 2 nsew clock input
flabel locali s 1230 357 1264 391 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 30 289 64 323 0 FreeSans 200 0 0 0 GATE_N
port 2 nsew clock input
flabel locali s 1230 425 1264 459 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 1230 85 1264 119 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 1230 289 1264 323 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel metal1 s 46 0 46 0 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel metal1 s 47 544 47 544 0 FreeSans 200 0 0 0 VPWR
port 7 nsew
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel nwell s 47 544 47 544 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel nwell s 47 544 47 544 0 FreeSans 200 0 0 0 VPB
port 6 nsew
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel pwell s 47 0 47 0 0 FreeSans 200 0 0 0 VNB
port 5 nsew
flabel pwell s 47 0 47 0 0 FreeSans 200 0 0 0 VNB
port 5 nsew
rlabel comment s 0 0 0 0 4 dlrtn_1
rlabel metal1 s 0 -48 1288 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1288 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1288 544
string GDS_END 2709276
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2697696
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
