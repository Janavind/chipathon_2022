magic
tech sky130A
magscale 1 2
timestamp 1666464484
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 2 67 631 203
rect 2 21 443 67
rect 30 -17 64 21
<< scnmos >>
rect 83 47 113 177
rect 167 47 197 177
rect 251 47 281 177
rect 335 47 365 177
rect 523 93 553 177
<< scpmoshvt >>
rect 83 297 113 497
rect 167 297 197 497
rect 251 297 281 497
rect 335 297 365 497
rect 523 413 553 497
<< ndiff >>
rect 28 163 83 177
rect 28 129 39 163
rect 73 129 83 163
rect 28 95 83 129
rect 28 61 39 95
rect 73 61 83 95
rect 28 47 83 61
rect 113 163 167 177
rect 113 129 123 163
rect 157 129 167 163
rect 113 95 167 129
rect 113 61 123 95
rect 157 61 167 95
rect 113 47 167 61
rect 197 95 251 177
rect 197 61 207 95
rect 241 61 251 95
rect 197 47 251 61
rect 281 163 335 177
rect 281 129 291 163
rect 325 129 335 163
rect 281 95 335 129
rect 281 61 291 95
rect 325 61 335 95
rect 281 47 335 61
rect 365 163 417 177
rect 365 129 375 163
rect 409 129 417 163
rect 365 95 417 129
rect 365 61 375 95
rect 409 61 417 95
rect 471 153 523 177
rect 471 119 479 153
rect 513 119 523 153
rect 471 93 523 119
rect 553 153 605 177
rect 553 119 563 153
rect 597 119 605 153
rect 553 93 605 119
rect 365 47 417 61
<< pdiff >>
rect 27 477 83 497
rect 27 443 39 477
rect 73 443 83 477
rect 27 409 83 443
rect 27 375 39 409
rect 73 375 83 409
rect 27 341 83 375
rect 27 307 39 341
rect 73 307 83 341
rect 27 297 83 307
rect 113 485 167 497
rect 113 451 123 485
rect 157 451 167 485
rect 113 417 167 451
rect 113 383 123 417
rect 157 383 167 417
rect 113 297 167 383
rect 197 477 251 497
rect 197 443 207 477
rect 241 443 251 477
rect 197 409 251 443
rect 197 375 207 409
rect 241 375 251 409
rect 197 341 251 375
rect 197 307 207 341
rect 241 307 251 341
rect 197 297 251 307
rect 281 409 335 497
rect 281 375 291 409
rect 325 375 335 409
rect 281 341 335 375
rect 281 307 291 341
rect 325 307 335 341
rect 281 297 335 307
rect 365 479 417 497
rect 365 445 375 479
rect 409 445 417 479
rect 365 411 417 445
rect 471 473 523 497
rect 471 439 479 473
rect 513 439 523 473
rect 471 413 523 439
rect 553 479 605 497
rect 553 445 563 479
rect 597 445 605 479
rect 553 413 605 445
rect 365 377 375 411
rect 409 377 417 411
rect 365 343 417 377
rect 365 309 375 343
rect 409 309 417 343
rect 365 297 417 309
<< ndiffc >>
rect 39 129 73 163
rect 39 61 73 95
rect 123 129 157 163
rect 123 61 157 95
rect 207 61 241 95
rect 291 129 325 163
rect 291 61 325 95
rect 375 129 409 163
rect 375 61 409 95
rect 479 119 513 153
rect 563 119 597 153
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 39 307 73 341
rect 123 451 157 485
rect 123 383 157 417
rect 207 443 241 477
rect 207 375 241 409
rect 207 307 241 341
rect 291 375 325 409
rect 291 307 325 341
rect 375 445 409 479
rect 479 439 513 473
rect 563 445 597 479
rect 375 377 409 411
rect 375 309 409 343
<< poly >>
rect 83 497 113 523
rect 167 497 197 523
rect 251 497 281 523
rect 335 497 365 523
rect 523 497 553 523
rect 83 265 113 297
rect 167 265 197 297
rect 83 249 197 265
rect 83 215 112 249
rect 146 215 197 249
rect 83 199 197 215
rect 83 177 113 199
rect 167 177 197 199
rect 251 265 281 297
rect 335 265 365 297
rect 523 265 553 413
rect 251 249 441 265
rect 251 215 391 249
rect 425 215 441 249
rect 251 199 441 215
rect 523 249 580 265
rect 523 215 536 249
rect 570 215 580 249
rect 523 199 580 215
rect 251 177 281 199
rect 335 177 365 199
rect 523 177 553 199
rect 83 21 113 47
rect 167 21 197 47
rect 251 21 281 47
rect 335 21 365 47
rect 523 21 553 93
<< polycont >>
rect 112 215 146 249
rect 391 215 425 249
rect 536 215 570 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 17 477 81 493
rect 17 443 39 477
rect 73 443 81 477
rect 17 409 81 443
rect 17 375 39 409
rect 73 375 81 409
rect 17 341 81 375
rect 115 485 165 527
rect 115 451 123 485
rect 157 451 165 485
rect 115 417 165 451
rect 115 383 123 417
rect 157 383 165 417
rect 115 365 165 383
rect 199 479 425 493
rect 199 477 375 479
rect 199 443 207 477
rect 241 459 375 477
rect 241 443 249 459
rect 199 409 249 443
rect 367 445 375 459
rect 409 445 425 479
rect 199 375 207 409
rect 241 375 249 409
rect 17 307 39 341
rect 73 331 81 341
rect 199 341 249 375
rect 199 331 207 341
rect 73 307 207 331
rect 241 307 249 341
rect 17 289 249 307
rect 283 409 333 425
rect 283 375 291 409
rect 325 375 333 409
rect 283 341 333 375
rect 283 307 291 341
rect 325 307 333 341
rect 96 249 184 255
rect 96 215 112 249
rect 146 215 184 249
rect 96 213 184 215
rect 283 179 333 307
rect 367 411 425 445
rect 367 377 375 411
rect 409 378 425 411
rect 479 473 513 492
rect 409 377 418 378
rect 367 343 418 377
rect 367 309 375 343
rect 409 309 418 343
rect 479 323 513 439
rect 555 479 605 527
rect 555 445 563 479
rect 597 445 605 479
rect 555 429 605 445
rect 367 289 418 309
rect 452 289 513 323
rect 452 249 486 289
rect 582 255 625 393
rect 375 215 391 249
rect 425 215 486 249
rect 443 179 486 215
rect 520 249 625 255
rect 520 215 536 249
rect 570 215 625 249
rect 520 213 625 215
rect 17 163 73 179
rect 17 129 39 163
rect 17 95 73 129
rect 17 61 39 95
rect 17 17 73 61
rect 107 163 341 179
rect 107 129 123 163
rect 157 145 291 163
rect 157 129 173 145
rect 107 95 173 129
rect 275 129 291 145
rect 325 129 341 163
rect 107 61 123 95
rect 157 61 173 95
rect 107 51 173 61
rect 207 95 241 111
rect 207 17 241 61
rect 275 95 341 129
rect 275 61 291 95
rect 325 61 341 95
rect 275 51 341 61
rect 375 163 409 179
rect 443 153 513 179
rect 443 145 479 153
rect 375 95 409 129
rect 479 89 513 119
rect 555 153 606 169
rect 555 119 563 153
rect 597 119 606 153
rect 375 17 409 61
rect 555 17 606 119
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
flabel locali s 582 221 616 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 122 221 156 255 0 FreeSans 200 0 0 0 SLEEP
port 2 nsew signal input
flabel locali s 306 85 340 119 0 FreeSans 400 0 0 0 X
port 7 nsew signal output
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 lpflow_isobufsrc_2
rlabel metal1 s 0 -48 644 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 644 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 644 544
string GDS_END 2363572
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2357630
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 16.100 0.000 
<< end >>
