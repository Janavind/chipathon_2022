magic
tech sky130B
magscale 1 2
timestamp 1666464484
<< nwell >>
rect 0 2152 1591 2424
rect 0 272 272 2152
rect 1319 272 1591 2152
rect 0 0 1591 272
<< pwell >>
rect 332 332 1259 2092
<< locali >>
rect 66 2305 1525 2358
rect 66 2271 307 2305
rect 341 2271 379 2305
rect 413 2271 451 2305
rect 485 2271 523 2305
rect 557 2271 595 2305
rect 629 2271 959 2305
rect 993 2271 1031 2305
rect 1065 2271 1103 2305
rect 1137 2271 1175 2305
rect 1209 2271 1247 2305
rect 1281 2271 1525 2305
rect 66 2218 1525 2271
rect 66 2035 206 2218
rect 66 2001 119 2035
rect 153 2001 206 2035
rect 66 1963 206 2001
rect 66 1929 119 1963
rect 153 1929 206 1963
rect 66 1891 206 1929
rect 66 1857 119 1891
rect 153 1857 206 1891
rect 66 1819 206 1857
rect 66 1785 119 1819
rect 153 1785 206 1819
rect 66 1747 206 1785
rect 66 1713 119 1747
rect 153 1713 206 1747
rect 66 1675 206 1713
rect 66 1641 119 1675
rect 153 1641 206 1675
rect 66 1603 206 1641
rect 66 1569 119 1603
rect 153 1569 206 1603
rect 66 1531 206 1569
rect 66 1497 119 1531
rect 153 1497 206 1531
rect 66 1459 206 1497
rect 66 1425 119 1459
rect 153 1425 206 1459
rect 66 1387 206 1425
rect 66 1353 119 1387
rect 153 1353 206 1387
rect 66 1315 206 1353
rect 66 1281 119 1315
rect 153 1281 206 1315
rect 66 1243 206 1281
rect 66 1209 119 1243
rect 153 1209 206 1243
rect 66 1171 206 1209
rect 66 1137 119 1171
rect 153 1137 206 1171
rect 66 1099 206 1137
rect 66 1065 119 1099
rect 153 1065 206 1099
rect 66 1027 206 1065
rect 66 993 119 1027
rect 153 993 206 1027
rect 66 955 206 993
rect 66 921 119 955
rect 153 921 206 955
rect 66 883 206 921
rect 66 849 119 883
rect 153 849 206 883
rect 66 811 206 849
rect 66 777 119 811
rect 153 777 206 811
rect 66 739 206 777
rect 66 705 119 739
rect 153 705 206 739
rect 66 667 206 705
rect 66 633 119 667
rect 153 633 206 667
rect 66 595 206 633
rect 66 561 119 595
rect 153 561 206 595
rect 66 523 206 561
rect 66 489 119 523
rect 153 489 206 523
rect 66 451 206 489
rect 66 417 119 451
rect 153 417 206 451
rect 66 379 206 417
rect 66 345 119 379
rect 153 345 206 379
rect 358 2003 1233 2066
rect 358 1969 454 2003
rect 488 1969 526 2003
rect 560 1969 598 2003
rect 632 1969 928 2003
rect 962 1969 1000 2003
rect 1034 1969 1072 2003
rect 1106 1969 1233 2003
rect 358 1924 1233 1969
rect 358 1803 498 1924
rect 358 1769 395 1803
rect 429 1769 498 1803
rect 662 1847 927 1867
rect 662 1813 725 1847
rect 759 1813 797 1847
rect 831 1813 927 1847
rect 662 1785 927 1813
rect 1093 1803 1233 1924
rect 358 1731 498 1769
rect 1093 1769 1146 1803
rect 1180 1769 1233 1803
rect 358 1697 395 1731
rect 429 1697 498 1731
rect 358 1659 498 1697
rect 358 1625 395 1659
rect 429 1625 498 1659
rect 358 1587 498 1625
rect 358 1553 395 1587
rect 429 1553 498 1587
rect 358 1515 498 1553
rect 358 1481 395 1515
rect 429 1481 498 1515
rect 358 1443 498 1481
rect 358 1409 395 1443
rect 429 1409 498 1443
rect 358 1371 498 1409
rect 358 1337 395 1371
rect 429 1337 498 1371
rect 358 1299 498 1337
rect 358 1265 395 1299
rect 429 1265 498 1299
rect 358 1227 498 1265
rect 358 1193 395 1227
rect 429 1193 498 1227
rect 358 1155 498 1193
rect 358 1121 395 1155
rect 429 1121 498 1155
rect 358 1083 498 1121
rect 358 1049 395 1083
rect 429 1049 498 1083
rect 358 1011 498 1049
rect 358 977 395 1011
rect 429 977 498 1011
rect 358 939 498 977
rect 358 905 395 939
rect 429 905 498 939
rect 358 867 498 905
rect 358 833 395 867
rect 429 833 498 867
rect 358 795 498 833
rect 358 761 395 795
rect 429 761 498 795
rect 358 723 498 761
rect 358 689 395 723
rect 429 689 498 723
rect 358 651 498 689
rect 593 1583 701 1751
rect 593 1549 621 1583
rect 655 1549 701 1583
rect 593 1511 701 1549
rect 593 1477 621 1511
rect 655 1477 701 1511
rect 593 1439 701 1477
rect 593 1405 621 1439
rect 655 1405 701 1439
rect 593 1367 701 1405
rect 593 1333 621 1367
rect 655 1333 701 1367
rect 593 1295 701 1333
rect 593 1261 621 1295
rect 655 1261 701 1295
rect 593 1223 701 1261
rect 593 1189 621 1223
rect 655 1189 701 1223
rect 593 1151 701 1189
rect 593 1117 621 1151
rect 655 1117 701 1151
rect 593 1079 701 1117
rect 593 1045 621 1079
rect 655 1045 701 1079
rect 593 1007 701 1045
rect 593 973 621 1007
rect 655 973 701 1007
rect 593 935 701 973
rect 593 901 621 935
rect 655 901 701 935
rect 593 863 701 901
rect 593 829 621 863
rect 655 829 701 863
rect 593 791 701 829
rect 593 757 621 791
rect 655 757 701 791
rect 593 672 701 757
rect 888 1583 996 1751
rect 888 1549 915 1583
rect 949 1549 996 1583
rect 888 1511 996 1549
rect 888 1477 915 1511
rect 949 1477 996 1511
rect 888 1439 996 1477
rect 888 1405 915 1439
rect 949 1405 996 1439
rect 888 1367 996 1405
rect 888 1333 915 1367
rect 949 1333 996 1367
rect 888 1295 996 1333
rect 888 1261 915 1295
rect 949 1261 996 1295
rect 888 1223 996 1261
rect 888 1189 915 1223
rect 949 1189 996 1223
rect 888 1151 996 1189
rect 888 1117 915 1151
rect 949 1117 996 1151
rect 888 1079 996 1117
rect 888 1045 915 1079
rect 949 1045 996 1079
rect 888 1007 996 1045
rect 888 973 915 1007
rect 949 973 996 1007
rect 888 935 996 973
rect 888 901 915 935
rect 949 901 996 935
rect 888 863 996 901
rect 888 829 915 863
rect 949 829 996 863
rect 888 791 996 829
rect 888 757 915 791
rect 949 757 996 791
rect 888 672 996 757
rect 1093 1731 1233 1769
rect 1093 1697 1146 1731
rect 1180 1697 1233 1731
rect 1093 1659 1233 1697
rect 1093 1625 1146 1659
rect 1180 1625 1233 1659
rect 1093 1587 1233 1625
rect 1093 1553 1146 1587
rect 1180 1553 1233 1587
rect 1093 1515 1233 1553
rect 1093 1481 1146 1515
rect 1180 1481 1233 1515
rect 1093 1443 1233 1481
rect 1093 1409 1146 1443
rect 1180 1409 1233 1443
rect 1093 1371 1233 1409
rect 1093 1337 1146 1371
rect 1180 1337 1233 1371
rect 1093 1299 1233 1337
rect 1093 1265 1146 1299
rect 1180 1265 1233 1299
rect 1093 1227 1233 1265
rect 1093 1193 1146 1227
rect 1180 1193 1233 1227
rect 1093 1155 1233 1193
rect 1093 1121 1146 1155
rect 1180 1121 1233 1155
rect 1093 1083 1233 1121
rect 1093 1049 1146 1083
rect 1180 1049 1233 1083
rect 1093 1011 1233 1049
rect 1093 977 1146 1011
rect 1180 977 1233 1011
rect 1093 939 1233 977
rect 1093 905 1146 939
rect 1180 905 1233 939
rect 1093 867 1233 905
rect 1093 833 1146 867
rect 1180 833 1233 867
rect 1093 795 1233 833
rect 1093 761 1146 795
rect 1180 761 1233 795
rect 1093 723 1233 761
rect 1093 689 1146 723
rect 1180 689 1233 723
rect 358 617 395 651
rect 429 617 498 651
rect 358 579 498 617
rect 358 545 395 579
rect 429 545 498 579
rect 358 507 498 545
rect 358 473 395 507
rect 429 498 498 507
rect 1093 651 1233 689
rect 1093 617 1146 651
rect 1180 617 1233 651
rect 1093 579 1233 617
rect 1093 545 1146 579
rect 1180 545 1233 579
rect 1093 507 1233 545
rect 1093 498 1146 507
rect 429 473 1146 498
rect 1180 473 1233 507
rect 358 435 1233 473
rect 358 401 395 435
rect 429 401 1146 435
rect 1180 401 1233 435
rect 358 358 1233 401
rect 1385 2035 1525 2218
rect 1385 2001 1438 2035
rect 1472 2001 1525 2035
rect 1385 1963 1525 2001
rect 1385 1929 1438 1963
rect 1472 1929 1525 1963
rect 1385 1891 1525 1929
rect 1385 1857 1438 1891
rect 1472 1857 1525 1891
rect 1385 1819 1525 1857
rect 1385 1785 1438 1819
rect 1472 1785 1525 1819
rect 1385 1747 1525 1785
rect 1385 1713 1438 1747
rect 1472 1713 1525 1747
rect 1385 1675 1525 1713
rect 1385 1641 1438 1675
rect 1472 1641 1525 1675
rect 1385 1603 1525 1641
rect 1385 1569 1438 1603
rect 1472 1569 1525 1603
rect 1385 1531 1525 1569
rect 1385 1497 1438 1531
rect 1472 1497 1525 1531
rect 1385 1459 1525 1497
rect 1385 1425 1438 1459
rect 1472 1425 1525 1459
rect 1385 1387 1525 1425
rect 1385 1353 1438 1387
rect 1472 1353 1525 1387
rect 1385 1315 1525 1353
rect 1385 1281 1438 1315
rect 1472 1281 1525 1315
rect 1385 1243 1525 1281
rect 1385 1209 1438 1243
rect 1472 1209 1525 1243
rect 1385 1171 1525 1209
rect 1385 1137 1438 1171
rect 1472 1137 1525 1171
rect 1385 1099 1525 1137
rect 1385 1065 1438 1099
rect 1472 1065 1525 1099
rect 1385 1027 1525 1065
rect 1385 993 1438 1027
rect 1472 993 1525 1027
rect 1385 955 1525 993
rect 1385 921 1438 955
rect 1472 921 1525 955
rect 1385 883 1525 921
rect 1385 849 1438 883
rect 1472 849 1525 883
rect 1385 811 1525 849
rect 1385 777 1438 811
rect 1472 777 1525 811
rect 1385 739 1525 777
rect 1385 705 1438 739
rect 1472 705 1525 739
rect 1385 667 1525 705
rect 1385 633 1438 667
rect 1472 633 1525 667
rect 1385 595 1525 633
rect 1385 561 1438 595
rect 1472 561 1525 595
rect 1385 523 1525 561
rect 1385 489 1438 523
rect 1472 489 1525 523
rect 1385 451 1525 489
rect 1385 417 1438 451
rect 1472 417 1525 451
rect 1385 379 1525 417
rect 66 307 206 345
rect 66 273 119 307
rect 153 273 206 307
rect 66 206 206 273
rect 1385 345 1438 379
rect 1472 345 1525 379
rect 1385 307 1525 345
rect 1385 273 1438 307
rect 1472 273 1525 307
rect 1385 206 1525 273
rect 66 142 1525 206
rect 66 108 1118 142
rect 1152 108 1190 142
rect 1224 108 1262 142
rect 1296 108 1525 142
rect 66 66 1525 108
<< viali >>
rect 307 2271 341 2305
rect 379 2271 413 2305
rect 451 2271 485 2305
rect 523 2271 557 2305
rect 595 2271 629 2305
rect 959 2271 993 2305
rect 1031 2271 1065 2305
rect 1103 2271 1137 2305
rect 1175 2271 1209 2305
rect 1247 2271 1281 2305
rect 119 2001 153 2035
rect 119 1929 153 1963
rect 119 1857 153 1891
rect 119 1785 153 1819
rect 119 1713 153 1747
rect 119 1641 153 1675
rect 119 1569 153 1603
rect 119 1497 153 1531
rect 119 1425 153 1459
rect 119 1353 153 1387
rect 119 1281 153 1315
rect 119 1209 153 1243
rect 119 1137 153 1171
rect 119 1065 153 1099
rect 119 993 153 1027
rect 119 921 153 955
rect 119 849 153 883
rect 119 777 153 811
rect 119 705 153 739
rect 119 633 153 667
rect 119 561 153 595
rect 119 489 153 523
rect 119 417 153 451
rect 119 345 153 379
rect 454 1969 488 2003
rect 526 1969 560 2003
rect 598 1969 632 2003
rect 928 1969 962 2003
rect 1000 1969 1034 2003
rect 1072 1969 1106 2003
rect 395 1769 429 1803
rect 725 1813 759 1847
rect 797 1813 831 1847
rect 1146 1769 1180 1803
rect 395 1697 429 1731
rect 395 1625 429 1659
rect 395 1553 429 1587
rect 395 1481 429 1515
rect 395 1409 429 1443
rect 395 1337 429 1371
rect 395 1265 429 1299
rect 395 1193 429 1227
rect 395 1121 429 1155
rect 395 1049 429 1083
rect 395 977 429 1011
rect 395 905 429 939
rect 395 833 429 867
rect 395 761 429 795
rect 395 689 429 723
rect 621 1549 655 1583
rect 621 1477 655 1511
rect 621 1405 655 1439
rect 621 1333 655 1367
rect 621 1261 655 1295
rect 621 1189 655 1223
rect 621 1117 655 1151
rect 621 1045 655 1079
rect 621 973 655 1007
rect 621 901 655 935
rect 621 829 655 863
rect 621 757 655 791
rect 915 1549 949 1583
rect 915 1477 949 1511
rect 915 1405 949 1439
rect 915 1333 949 1367
rect 915 1261 949 1295
rect 915 1189 949 1223
rect 915 1117 949 1151
rect 915 1045 949 1079
rect 915 973 949 1007
rect 915 901 949 935
rect 915 829 949 863
rect 915 757 949 791
rect 1146 1697 1180 1731
rect 1146 1625 1180 1659
rect 1146 1553 1180 1587
rect 1146 1481 1180 1515
rect 1146 1409 1180 1443
rect 1146 1337 1180 1371
rect 1146 1265 1180 1299
rect 1146 1193 1180 1227
rect 1146 1121 1180 1155
rect 1146 1049 1180 1083
rect 1146 977 1180 1011
rect 1146 905 1180 939
rect 1146 833 1180 867
rect 1146 761 1180 795
rect 1146 689 1180 723
rect 395 617 429 651
rect 395 545 429 579
rect 395 473 429 507
rect 1146 617 1180 651
rect 1146 545 1180 579
rect 1146 473 1180 507
rect 395 401 429 435
rect 1146 401 1180 435
rect 1438 2001 1472 2035
rect 1438 1929 1472 1963
rect 1438 1857 1472 1891
rect 1438 1785 1472 1819
rect 1438 1713 1472 1747
rect 1438 1641 1472 1675
rect 1438 1569 1472 1603
rect 1438 1497 1472 1531
rect 1438 1425 1472 1459
rect 1438 1353 1472 1387
rect 1438 1281 1472 1315
rect 1438 1209 1472 1243
rect 1438 1137 1472 1171
rect 1438 1065 1472 1099
rect 1438 993 1472 1027
rect 1438 921 1472 955
rect 1438 849 1472 883
rect 1438 777 1472 811
rect 1438 705 1472 739
rect 1438 633 1472 667
rect 1438 561 1472 595
rect 1438 489 1472 523
rect 1438 417 1472 451
rect 119 273 153 307
rect 1438 345 1472 379
rect 1438 273 1472 307
rect 1118 108 1152 142
rect 1190 108 1224 142
rect 1262 108 1296 142
<< metal1 >>
tri 66 2216 208 2358 se
rect 208 2305 669 2358
rect 208 2271 307 2305
rect 341 2271 379 2305
rect 413 2271 451 2305
rect 485 2271 523 2305
rect 557 2271 595 2305
rect 629 2271 669 2305
rect 208 2218 669 2271
rect 208 2216 286 2218
tri 286 2216 288 2218 nw
rect 66 2035 206 2216
tri 206 2136 286 2216 nw
rect 66 2001 119 2035
rect 153 2001 206 2035
rect 66 1963 206 2001
rect 66 1929 119 1963
rect 153 1929 206 1963
rect 66 1891 206 1929
rect 66 1857 119 1891
rect 153 1857 206 1891
rect 66 1819 206 1857
rect 66 1785 119 1819
rect 153 1785 206 1819
rect 66 1747 206 1785
rect 66 1713 119 1747
rect 153 1713 206 1747
rect 66 1675 206 1713
rect 66 1641 119 1675
rect 153 1641 206 1675
rect 66 1603 206 1641
rect 66 1569 119 1603
rect 153 1569 206 1603
rect 66 1531 206 1569
rect 66 1497 119 1531
rect 153 1497 206 1531
rect 66 1459 206 1497
rect 66 1425 119 1459
rect 153 1425 206 1459
rect 66 1387 206 1425
rect 66 1353 119 1387
rect 153 1353 206 1387
rect 66 1315 206 1353
rect 66 1281 119 1315
rect 153 1281 206 1315
rect 66 1243 206 1281
rect 66 1209 119 1243
rect 153 1209 206 1243
rect 66 1171 206 1209
rect 66 1137 119 1171
rect 153 1137 206 1171
rect 66 1099 206 1137
rect 66 1065 119 1099
rect 153 1065 206 1099
rect 66 1027 206 1065
rect 66 993 119 1027
rect 153 993 206 1027
rect 66 955 206 993
rect 66 921 119 955
rect 153 921 206 955
rect 66 883 206 921
rect 66 849 119 883
rect 153 849 206 883
rect 66 811 206 849
rect 66 777 119 811
rect 153 777 206 811
rect 66 739 206 777
rect 66 705 119 739
rect 153 705 206 739
rect 66 667 206 705
rect 66 633 119 667
rect 153 633 206 667
rect 66 595 206 633
rect 66 561 119 595
rect 153 561 206 595
rect 66 523 206 561
rect 66 489 119 523
rect 153 489 206 523
rect 66 451 206 489
rect 66 417 119 451
rect 153 417 206 451
rect 66 379 206 417
rect 66 345 119 379
rect 153 345 206 379
rect 66 307 206 345
rect 66 273 119 307
rect 153 273 206 307
rect 66 69 206 273
rect 66 66 203 69
tri 358 2000 424 2066 se
rect 424 2003 669 2066
rect 424 2000 454 2003
rect 358 1969 454 2000
rect 488 1969 526 2003
rect 560 1969 598 2003
rect 632 1969 669 2003
rect 358 1901 669 1969
rect 358 1803 536 1901
tri 536 1826 611 1901 nw
rect 703 1847 852 2359
rect 886 2305 1383 2358
rect 886 2271 959 2305
rect 993 2271 1031 2305
rect 1065 2271 1103 2305
rect 1137 2271 1175 2305
rect 1209 2271 1247 2305
rect 1281 2271 1383 2305
rect 886 2218 1383 2271
tri 1289 2216 1291 2218 ne
rect 1291 2216 1383 2218
tri 1383 2216 1525 2358 sw
tri 1291 2136 1371 2216 ne
rect 1371 2136 1525 2216
tri 1371 2124 1383 2136 ne
rect 1383 2124 1525 2136
tri 1383 2122 1385 2124 ne
rect 886 2003 1167 2066
rect 886 1969 928 2003
rect 962 1969 1000 2003
rect 1034 1969 1072 2003
rect 1106 2000 1167 2003
tri 1167 2000 1233 2066 sw
rect 1106 1969 1233 2000
rect 886 1901 1233 1969
rect 358 1769 395 1803
rect 429 1769 536 1803
rect 703 1813 725 1847
rect 759 1813 797 1847
rect 831 1813 852 1847
tri 1012 1826 1087 1901 ne
rect 1087 1826 1233 1901
tri 1087 1820 1093 1826 ne
rect 703 1791 852 1813
rect 1093 1803 1233 1826
rect 358 1731 536 1769
rect 1093 1769 1146 1803
rect 1180 1769 1233 1803
rect 358 1697 395 1731
rect 429 1697 536 1731
rect 358 1659 536 1697
rect 358 1625 395 1659
rect 429 1625 536 1659
rect 358 1587 536 1625
rect 358 1553 395 1587
rect 429 1553 536 1587
rect 358 1515 536 1553
rect 358 1481 395 1515
rect 429 1481 536 1515
rect 358 1443 536 1481
rect 358 1409 395 1443
rect 429 1409 536 1443
rect 358 1371 536 1409
rect 358 1337 395 1371
rect 429 1337 536 1371
rect 358 1299 536 1337
rect 358 1265 395 1299
rect 429 1265 536 1299
rect 358 1227 536 1265
rect 358 1193 395 1227
rect 429 1193 536 1227
rect 358 1155 536 1193
rect 358 1121 395 1155
rect 429 1121 536 1155
rect 358 1083 536 1121
rect 358 1049 395 1083
rect 429 1049 536 1083
rect 358 1011 536 1049
rect 358 977 395 1011
rect 429 977 536 1011
rect 358 939 536 977
rect 358 905 395 939
rect 429 905 536 939
rect 358 867 536 905
rect 358 833 395 867
rect 429 833 536 867
rect 358 795 536 833
rect 358 761 395 795
rect 429 761 536 795
rect 358 723 536 761
rect 358 689 395 723
rect 429 689 536 723
rect 358 651 536 689
rect 358 617 395 651
rect 429 617 536 651
rect 358 579 536 617
rect 358 545 395 579
rect 429 545 536 579
rect 358 507 536 545
rect 358 473 395 507
rect 429 473 536 507
rect 358 435 536 473
rect 358 401 395 435
rect 429 401 536 435
rect 358 69 536 401
rect 358 66 533 69
rect 572 1583 772 1709
rect 572 1549 621 1583
rect 655 1549 772 1583
rect 572 1511 772 1549
rect 572 1477 621 1511
rect 655 1477 772 1511
rect 572 1439 772 1477
rect 572 1405 621 1439
rect 655 1405 772 1439
rect 572 1367 772 1405
rect 572 1333 621 1367
rect 655 1333 772 1367
rect 572 1295 772 1333
rect 572 1261 621 1295
rect 655 1261 772 1295
rect 572 1223 772 1261
rect 572 1189 621 1223
rect 655 1189 772 1223
rect 572 1151 772 1189
rect 572 1117 621 1151
rect 655 1117 772 1151
rect 572 1079 772 1117
rect 572 1045 621 1079
rect 655 1045 772 1079
rect 572 1007 772 1045
rect 572 973 621 1007
rect 655 973 772 1007
rect 572 935 772 973
rect 572 901 621 935
rect 655 901 772 935
rect 572 863 772 901
rect 572 829 621 863
rect 655 829 772 863
rect 572 791 772 829
rect 572 757 621 791
rect 655 757 772 791
rect 572 66 772 757
rect 831 1583 1031 1752
rect 831 1549 915 1583
rect 949 1549 1031 1583
rect 831 1511 1031 1549
rect 831 1477 915 1511
rect 949 1477 1031 1511
rect 831 1439 1031 1477
rect 831 1405 915 1439
rect 949 1405 1031 1439
rect 831 1367 1031 1405
rect 831 1333 915 1367
rect 949 1333 1031 1367
rect 831 1295 1031 1333
rect 831 1261 915 1295
rect 949 1261 1031 1295
rect 831 1223 1031 1261
rect 831 1189 915 1223
rect 949 1189 1031 1223
rect 831 1151 1031 1189
rect 831 1117 915 1151
rect 949 1117 1031 1151
rect 831 1079 1031 1117
rect 831 1045 915 1079
rect 949 1045 1031 1079
rect 831 1007 1031 1045
rect 831 973 915 1007
rect 949 973 1031 1007
rect 831 935 1031 973
rect 831 901 915 935
rect 949 901 1031 935
rect 831 863 1031 901
rect 831 829 915 863
rect 949 829 1031 863
rect 831 791 1031 829
rect 831 757 915 791
rect 949 757 1031 791
rect 831 66 1031 757
rect 1093 1731 1233 1769
rect 1093 1697 1146 1731
rect 1180 1697 1233 1731
rect 1093 1659 1233 1697
rect 1093 1625 1146 1659
rect 1180 1625 1233 1659
rect 1093 1587 1233 1625
rect 1093 1553 1146 1587
rect 1180 1553 1233 1587
rect 1093 1515 1233 1553
rect 1093 1481 1146 1515
rect 1180 1481 1233 1515
rect 1093 1443 1233 1481
rect 1093 1409 1146 1443
rect 1180 1409 1233 1443
rect 1093 1371 1233 1409
rect 1093 1337 1146 1371
rect 1180 1337 1233 1371
rect 1093 1299 1233 1337
rect 1093 1265 1146 1299
rect 1180 1265 1233 1299
rect 1093 1227 1233 1265
rect 1093 1193 1146 1227
rect 1180 1193 1233 1227
rect 1093 1155 1233 1193
rect 1093 1121 1146 1155
rect 1180 1121 1233 1155
rect 1093 1083 1233 1121
rect 1093 1049 1146 1083
rect 1180 1049 1233 1083
rect 1093 1011 1233 1049
rect 1093 977 1146 1011
rect 1180 977 1233 1011
rect 1093 939 1233 977
rect 1093 905 1146 939
rect 1180 905 1233 939
rect 1093 867 1233 905
rect 1093 833 1146 867
rect 1180 833 1233 867
rect 1093 795 1233 833
rect 1093 761 1146 795
rect 1180 761 1233 795
rect 1093 723 1233 761
rect 1093 689 1146 723
rect 1180 689 1233 723
rect 1093 651 1233 689
rect 1093 617 1146 651
rect 1180 617 1233 651
rect 1093 579 1233 617
rect 1093 545 1146 579
rect 1180 545 1233 579
rect 1093 507 1233 545
rect 1093 473 1146 507
rect 1180 473 1233 507
rect 1093 435 1233 473
rect 1093 401 1146 435
rect 1180 401 1233 435
rect 1093 358 1233 401
rect 1385 2035 1525 2124
rect 1385 2001 1438 2035
rect 1472 2001 1525 2035
rect 1385 1963 1525 2001
rect 1385 1929 1438 1963
rect 1472 1929 1525 1963
rect 1385 1891 1525 1929
rect 1385 1857 1438 1891
rect 1472 1857 1525 1891
rect 1385 1819 1525 1857
rect 1385 1785 1438 1819
rect 1472 1785 1525 1819
rect 1385 1747 1525 1785
rect 1385 1713 1438 1747
rect 1472 1713 1525 1747
rect 1385 1675 1525 1713
rect 1385 1641 1438 1675
rect 1472 1641 1525 1675
rect 1385 1603 1525 1641
rect 1385 1569 1438 1603
rect 1472 1569 1525 1603
rect 1385 1531 1525 1569
rect 1385 1497 1438 1531
rect 1472 1497 1525 1531
rect 1385 1459 1525 1497
rect 1385 1425 1438 1459
rect 1472 1425 1525 1459
rect 1385 1387 1525 1425
rect 1385 1353 1438 1387
rect 1472 1353 1525 1387
rect 1385 1315 1525 1353
rect 1385 1281 1438 1315
rect 1472 1281 1525 1315
rect 1385 1243 1525 1281
rect 1385 1209 1438 1243
rect 1472 1209 1525 1243
rect 1385 1171 1525 1209
rect 1385 1137 1438 1171
rect 1472 1137 1525 1171
rect 1385 1099 1525 1137
rect 1385 1065 1438 1099
rect 1472 1065 1525 1099
rect 1385 1027 1525 1065
rect 1385 993 1438 1027
rect 1472 993 1525 1027
rect 1385 955 1525 993
rect 1385 921 1438 955
rect 1472 921 1525 955
rect 1385 883 1525 921
rect 1385 849 1438 883
rect 1472 849 1525 883
rect 1385 811 1525 849
rect 1385 777 1438 811
rect 1472 777 1525 811
rect 1385 739 1525 777
rect 1385 705 1438 739
rect 1472 705 1525 739
rect 1385 667 1525 705
rect 1385 633 1438 667
rect 1472 633 1525 667
rect 1385 595 1525 633
rect 1385 561 1438 595
rect 1472 561 1525 595
rect 1385 523 1525 561
rect 1385 489 1438 523
rect 1472 489 1525 523
rect 1385 451 1525 489
rect 1385 417 1438 451
rect 1472 417 1525 451
rect 1385 379 1525 417
rect 1385 345 1438 379
rect 1472 345 1525 379
rect 1385 307 1525 345
tri 1289 206 1385 302 se
rect 1385 273 1438 307
rect 1472 273 1525 307
rect 1385 208 1525 273
rect 1385 206 1386 208
rect 1070 142 1386 206
rect 1070 108 1118 142
rect 1152 108 1190 142
rect 1224 108 1262 142
rect 1296 108 1386 142
rect 1070 69 1386 108
tri 1386 69 1525 208 nw
rect 1070 66 1383 69
tri 1383 66 1386 69 nw
<< obsm1 >>
rect 203 66 206 69
rect 533 66 536 69
<< labels >>
rlabel metal1 s 703 1791 852 2359 6 GATE
port 1 nsew
rlabel viali s 797 1813 831 1847 6 GATE
port 1 nsew
rlabel viali s 725 1813 759 1847 6 GATE
port 1 nsew
rlabel locali s 662 1785 927 1867 6 GATE
port 1 nsew
rlabel metal1 s 1070 66 1383 69 6 NWELLRING
port 2 nsew
rlabel metal1 s 66 66 203 69 6 NWELLRING
port 2 nsew
rlabel metal1 s 1070 69 1386 206 6 NWELLRING
port 2 nsew
rlabel metal1 s 1385 206 1386 208 6 NWELLRING
port 2 nsew
rlabel metal1 s 1385 208 1525 2124 6 NWELLRING
port 2 nsew
rlabel metal1 s 1383 2124 1525 2136 6 NWELLRING
port 2 nsew
rlabel metal1 s 1371 2136 1525 2216 6 NWELLRING
port 2 nsew
rlabel metal1 s 66 69 206 2216 6 NWELLRING
port 2 nsew
rlabel metal1 s 1291 2216 1383 2218 6 NWELLRING
port 2 nsew
rlabel metal1 s 208 2216 286 2218 6 NWELLRING
port 2 nsew
rlabel metal1 s 886 2218 1383 2358 6 NWELLRING
port 2 nsew
rlabel metal1 s 208 2218 669 2358 6 NWELLRING
port 2 nsew
rlabel viali s 1262 108 1296 142 6 NWELLRING
port 2 nsew
rlabel viali s 1190 108 1224 142 6 NWELLRING
port 2 nsew
rlabel viali s 1118 108 1152 142 6 NWELLRING
port 2 nsew
rlabel viali s 1438 273 1472 307 6 NWELLRING
port 2 nsew
rlabel viali s 1438 345 1472 379 6 NWELLRING
port 2 nsew
rlabel viali s 1438 417 1472 451 6 NWELLRING
port 2 nsew
rlabel viali s 1438 489 1472 523 6 NWELLRING
port 2 nsew
rlabel viali s 1438 561 1472 595 6 NWELLRING
port 2 nsew
rlabel viali s 1438 633 1472 667 6 NWELLRING
port 2 nsew
rlabel viali s 1438 705 1472 739 6 NWELLRING
port 2 nsew
rlabel viali s 1438 777 1472 811 6 NWELLRING
port 2 nsew
rlabel viali s 1438 849 1472 883 6 NWELLRING
port 2 nsew
rlabel viali s 1438 921 1472 955 6 NWELLRING
port 2 nsew
rlabel viali s 1438 993 1472 1027 6 NWELLRING
port 2 nsew
rlabel viali s 1438 1065 1472 1099 6 NWELLRING
port 2 nsew
rlabel viali s 1438 1137 1472 1171 6 NWELLRING
port 2 nsew
rlabel viali s 1438 1209 1472 1243 6 NWELLRING
port 2 nsew
rlabel viali s 1438 1281 1472 1315 6 NWELLRING
port 2 nsew
rlabel viali s 1438 1353 1472 1387 6 NWELLRING
port 2 nsew
rlabel viali s 1438 1425 1472 1459 6 NWELLRING
port 2 nsew
rlabel viali s 1438 1497 1472 1531 6 NWELLRING
port 2 nsew
rlabel viali s 1438 1569 1472 1603 6 NWELLRING
port 2 nsew
rlabel viali s 1438 1641 1472 1675 6 NWELLRING
port 2 nsew
rlabel viali s 1438 1713 1472 1747 6 NWELLRING
port 2 nsew
rlabel viali s 1438 1785 1472 1819 6 NWELLRING
port 2 nsew
rlabel viali s 1438 1857 1472 1891 6 NWELLRING
port 2 nsew
rlabel viali s 1438 1929 1472 1963 6 NWELLRING
port 2 nsew
rlabel viali s 1438 2001 1472 2035 6 NWELLRING
port 2 nsew
rlabel viali s 119 273 153 307 6 NWELLRING
port 2 nsew
rlabel viali s 119 345 153 379 6 NWELLRING
port 2 nsew
rlabel viali s 119 417 153 451 6 NWELLRING
port 2 nsew
rlabel viali s 119 489 153 523 6 NWELLRING
port 2 nsew
rlabel viali s 119 561 153 595 6 NWELLRING
port 2 nsew
rlabel viali s 119 633 153 667 6 NWELLRING
port 2 nsew
rlabel viali s 119 705 153 739 6 NWELLRING
port 2 nsew
rlabel viali s 119 777 153 811 6 NWELLRING
port 2 nsew
rlabel viali s 119 849 153 883 6 NWELLRING
port 2 nsew
rlabel viali s 119 921 153 955 6 NWELLRING
port 2 nsew
rlabel viali s 119 993 153 1027 6 NWELLRING
port 2 nsew
rlabel viali s 119 1065 153 1099 6 NWELLRING
port 2 nsew
rlabel viali s 119 1137 153 1171 6 NWELLRING
port 2 nsew
rlabel viali s 119 1209 153 1243 6 NWELLRING
port 2 nsew
rlabel viali s 119 1281 153 1315 6 NWELLRING
port 2 nsew
rlabel viali s 119 1353 153 1387 6 NWELLRING
port 2 nsew
rlabel viali s 119 1425 153 1459 6 NWELLRING
port 2 nsew
rlabel viali s 119 1497 153 1531 6 NWELLRING
port 2 nsew
rlabel viali s 119 1569 153 1603 6 NWELLRING
port 2 nsew
rlabel viali s 119 1641 153 1675 6 NWELLRING
port 2 nsew
rlabel viali s 119 1713 153 1747 6 NWELLRING
port 2 nsew
rlabel viali s 119 1785 153 1819 6 NWELLRING
port 2 nsew
rlabel viali s 119 1857 153 1891 6 NWELLRING
port 2 nsew
rlabel viali s 119 1929 153 1963 6 NWELLRING
port 2 nsew
rlabel viali s 119 2001 153 2035 6 NWELLRING
port 2 nsew
rlabel viali s 1247 2271 1281 2305 6 NWELLRING
port 2 nsew
rlabel viali s 1175 2271 1209 2305 6 NWELLRING
port 2 nsew
rlabel viali s 1103 2271 1137 2305 6 NWELLRING
port 2 nsew
rlabel viali s 1031 2271 1065 2305 6 NWELLRING
port 2 nsew
rlabel viali s 959 2271 993 2305 6 NWELLRING
port 2 nsew
rlabel viali s 595 2271 629 2305 6 NWELLRING
port 2 nsew
rlabel viali s 523 2271 557 2305 6 NWELLRING
port 2 nsew
rlabel viali s 451 2271 485 2305 6 NWELLRING
port 2 nsew
rlabel viali s 379 2271 413 2305 6 NWELLRING
port 2 nsew
rlabel viali s 307 2271 341 2305 6 NWELLRING
port 2 nsew
rlabel locali s 66 66 1525 206 6 NWELLRING
port 2 nsew
rlabel locali s 1385 206 1525 2218 6 NWELLRING
port 2 nsew
rlabel locali s 66 206 206 2218 6 NWELLRING
port 2 nsew
rlabel locali s 66 2218 1525 2358 6 NWELLRING
port 2 nsew
rlabel nwell s 0 0 1591 272 6 NWELLRING
port 2 nsew
rlabel nwell s 1319 272 1591 2152 6 NWELLRING
port 2 nsew
rlabel nwell s 0 272 272 2152 6 NWELLRING
port 2 nsew
rlabel nwell s 0 2152 1591 2424 6 NWELLRING
port 2 nsew
rlabel metal1 s 572 66 772 1709 6 VGND
port 3 nsew ground default
rlabel viali s 621 757 655 791 6 VGND
port 3 nsew ground default
rlabel viali s 621 829 655 863 6 VGND
port 3 nsew ground default
rlabel viali s 621 901 655 935 6 VGND
port 3 nsew ground default
rlabel viali s 621 973 655 1007 6 VGND
port 3 nsew ground default
rlabel viali s 621 1045 655 1079 6 VGND
port 3 nsew ground default
rlabel viali s 621 1117 655 1151 6 VGND
port 3 nsew ground default
rlabel viali s 621 1189 655 1223 6 VGND
port 3 nsew ground default
rlabel viali s 621 1261 655 1295 6 VGND
port 3 nsew ground default
rlabel viali s 621 1333 655 1367 6 VGND
port 3 nsew ground default
rlabel viali s 621 1405 655 1439 6 VGND
port 3 nsew ground default
rlabel viali s 621 1477 655 1511 6 VGND
port 3 nsew ground default
rlabel viali s 621 1549 655 1583 6 VGND
port 3 nsew ground default
rlabel locali s 593 672 701 1751 6 VGND
port 3 nsew ground default
rlabel metal1 s 358 66 533 69 6 NBODY
port 4 nsew
rlabel metal1 s 1093 358 1233 1826 6 NBODY
port 4 nsew
rlabel metal1 s 1087 1826 1233 1901 6 NBODY
port 4 nsew
rlabel metal1 s 358 69 536 1901 6 NBODY
port 4 nsew
rlabel metal1 s 886 1901 1233 2000 6 NBODY
port 4 nsew
rlabel metal1 s 886 2000 1167 2066 6 NBODY
port 4 nsew
rlabel metal1 s 358 1901 669 2000 6 NBODY
port 4 nsew
rlabel metal1 s 424 2000 669 2066 6 NBODY
port 4 nsew
rlabel viali s 1146 401 1180 435 6 NBODY
port 4 nsew
rlabel viali s 395 401 429 435 6 NBODY
port 4 nsew
rlabel viali s 1146 473 1180 507 6 NBODY
port 4 nsew
rlabel viali s 1146 545 1180 579 6 NBODY
port 4 nsew
rlabel viali s 1146 617 1180 651 6 NBODY
port 4 nsew
rlabel viali s 1146 689 1180 723 6 NBODY
port 4 nsew
rlabel viali s 1146 761 1180 795 6 NBODY
port 4 nsew
rlabel viali s 1146 833 1180 867 6 NBODY
port 4 nsew
rlabel viali s 1146 905 1180 939 6 NBODY
port 4 nsew
rlabel viali s 1146 977 1180 1011 6 NBODY
port 4 nsew
rlabel viali s 1146 1049 1180 1083 6 NBODY
port 4 nsew
rlabel viali s 1146 1121 1180 1155 6 NBODY
port 4 nsew
rlabel viali s 1146 1193 1180 1227 6 NBODY
port 4 nsew
rlabel viali s 1146 1265 1180 1299 6 NBODY
port 4 nsew
rlabel viali s 1146 1337 1180 1371 6 NBODY
port 4 nsew
rlabel viali s 1146 1409 1180 1443 6 NBODY
port 4 nsew
rlabel viali s 1146 1481 1180 1515 6 NBODY
port 4 nsew
rlabel viali s 1146 1553 1180 1587 6 NBODY
port 4 nsew
rlabel viali s 1146 1625 1180 1659 6 NBODY
port 4 nsew
rlabel viali s 1146 1697 1180 1731 6 NBODY
port 4 nsew
rlabel viali s 1146 1769 1180 1803 6 NBODY
port 4 nsew
rlabel viali s 395 473 429 507 6 NBODY
port 4 nsew
rlabel viali s 395 545 429 579 6 NBODY
port 4 nsew
rlabel viali s 395 617 429 651 6 NBODY
port 4 nsew
rlabel viali s 395 689 429 723 6 NBODY
port 4 nsew
rlabel viali s 395 761 429 795 6 NBODY
port 4 nsew
rlabel viali s 395 833 429 867 6 NBODY
port 4 nsew
rlabel viali s 395 905 429 939 6 NBODY
port 4 nsew
rlabel viali s 395 977 429 1011 6 NBODY
port 4 nsew
rlabel viali s 395 1049 429 1083 6 NBODY
port 4 nsew
rlabel viali s 395 1121 429 1155 6 NBODY
port 4 nsew
rlabel viali s 395 1193 429 1227 6 NBODY
port 4 nsew
rlabel viali s 395 1265 429 1299 6 NBODY
port 4 nsew
rlabel viali s 395 1337 429 1371 6 NBODY
port 4 nsew
rlabel viali s 395 1409 429 1443 6 NBODY
port 4 nsew
rlabel viali s 395 1481 429 1515 6 NBODY
port 4 nsew
rlabel viali s 395 1553 429 1587 6 NBODY
port 4 nsew
rlabel viali s 395 1625 429 1659 6 NBODY
port 4 nsew
rlabel viali s 395 1697 429 1731 6 NBODY
port 4 nsew
rlabel viali s 395 1769 429 1803 6 NBODY
port 4 nsew
rlabel viali s 1072 1969 1106 2003 6 NBODY
port 4 nsew
rlabel viali s 1000 1969 1034 2003 6 NBODY
port 4 nsew
rlabel viali s 928 1969 962 2003 6 NBODY
port 4 nsew
rlabel viali s 598 1969 632 2003 6 NBODY
port 4 nsew
rlabel viali s 526 1969 560 2003 6 NBODY
port 4 nsew
rlabel viali s 454 1969 488 2003 6 NBODY
port 4 nsew
rlabel locali s 358 358 1233 498 6 NBODY
port 4 nsew
rlabel locali s 1093 498 1233 1924 6 NBODY
port 4 nsew
rlabel locali s 358 498 498 1924 6 NBODY
port 4 nsew
rlabel locali s 358 1924 1233 2066 6 NBODY
port 4 nsew
rlabel pwell s 332 332 1259 2092 6 NBODY
port 4 nsew
rlabel metal1 s 831 66 1031 1752 6 IN
port 5 nsew
rlabel viali s 915 757 949 791 6 IN
port 5 nsew
rlabel viali s 915 829 949 863 6 IN
port 5 nsew
rlabel viali s 915 901 949 935 6 IN
port 5 nsew
rlabel viali s 915 973 949 1007 6 IN
port 5 nsew
rlabel viali s 915 1045 949 1079 6 IN
port 5 nsew
rlabel viali s 915 1117 949 1151 6 IN
port 5 nsew
rlabel viali s 915 1189 949 1223 6 IN
port 5 nsew
rlabel viali s 915 1261 949 1295 6 IN
port 5 nsew
rlabel viali s 915 1333 949 1367 6 IN
port 5 nsew
rlabel viali s 915 1405 949 1439 6 IN
port 5 nsew
rlabel viali s 915 1477 949 1511 6 IN
port 5 nsew
rlabel viali s 915 1549 949 1583 6 IN
port 5 nsew
rlabel locali s 888 672 996 1751 6 IN
port 5 nsew
<< properties >>
string FIXED_BBOX 0 0 1591 2424
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 3868322
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 3863558
<< end >>
