magic
tech sky130A
magscale 1 2
timestamp 1666199351
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_0
timestamp 1666199351
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_1
timestamp 1666199351
transform 1 0 36 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_2
timestamp 1666199351
transform 1 0 128 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_3
timestamp 1666199351
transform 1 0 220 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_4
timestamp 1666199351
transform 1 0 312 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_5
timestamp 1666199351
transform 1 0 404 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_6
timestamp 1666199351
transform 1 0 496 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_7
timestamp 1666199351
transform 1 0 588 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_8
timestamp 1666199351
transform 1 0 680 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_9
timestamp 1666199351
transform 1 0 772 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_10
timestamp 1666199351
transform 1 0 864 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 8190306
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 8184736
<< end >>
