magic
tech sky130A
magscale 1 2
timestamp 1666199351
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 1 21 640 203
rect 29 -17 63 21
<< locali >>
rect 388 333 454 493
rect 328 299 454 333
rect 17 197 87 257
rect 121 199 200 265
rect 121 56 165 199
rect 328 158 362 299
rect 489 265 523 485
rect 406 215 523 265
rect 557 215 627 257
rect 312 86 362 158
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 30 291 80 527
rect 114 333 164 493
rect 198 367 354 527
rect 114 299 268 333
rect 234 265 268 299
rect 234 199 294 265
rect 18 17 85 163
rect 234 165 268 199
rect 200 56 268 165
rect 564 291 614 527
rect 396 145 622 181
rect 396 85 454 145
rect 488 17 522 111
rect 556 55 622 145
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel locali s 17 197 87 257 6 A1_N
port 1 nsew signal input
rlabel locali s 121 56 165 199 6 A2_N
port 2 nsew signal input
rlabel locali s 121 199 200 265 6 A2_N
port 2 nsew signal input
rlabel locali s 557 215 627 257 6 B1
port 3 nsew signal input
rlabel locali s 406 215 523 265 6 B2
port 4 nsew signal input
rlabel locali s 489 265 523 485 6 B2
port 4 nsew signal input
rlabel metal1 s 0 -48 644 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 21 640 203 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 682 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 644 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 312 86 362 158 6 Y
port 9 nsew signal output
rlabel locali s 328 158 362 299 6 Y
port 9 nsew signal output
rlabel locali s 328 299 454 333 6 Y
port 9 nsew signal output
rlabel locali s 388 333 454 493 6 Y
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 644 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1241466
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1235296
<< end >>
