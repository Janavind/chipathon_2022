magic
tech sky130B
magscale 1 2
timestamp 1666464484
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 1 21 558 203
rect 31 -17 65 21
<< scnmos >>
rect 79 47 109 177
rect 164 47 194 177
rect 250 47 280 177
rect 351 47 381 177
rect 450 47 480 177
<< scpmoshvt >>
rect 79 297 109 497
rect 164 297 194 497
rect 250 297 280 497
rect 346 297 376 497
rect 445 297 475 497
<< ndiff >>
rect 27 161 79 177
rect 27 127 35 161
rect 69 127 79 161
rect 27 93 79 127
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 47 164 177
rect 194 47 250 177
rect 280 101 351 177
rect 280 67 307 101
rect 341 67 351 101
rect 280 47 351 67
rect 381 97 450 177
rect 381 63 397 97
rect 431 63 450 97
rect 381 47 450 63
rect 480 129 532 177
rect 480 95 490 129
rect 524 95 532 129
rect 480 47 532 95
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 349 79 383
rect 27 315 35 349
rect 69 315 79 349
rect 27 297 79 315
rect 109 445 164 497
rect 109 411 120 445
rect 154 411 164 445
rect 109 377 164 411
rect 109 343 120 377
rect 154 343 164 377
rect 109 297 164 343
rect 194 433 250 497
rect 194 399 204 433
rect 238 399 250 433
rect 194 297 250 399
rect 280 469 346 497
rect 280 435 290 469
rect 324 435 346 469
rect 280 297 346 435
rect 376 297 445 497
rect 475 433 527 497
rect 475 399 485 433
rect 519 399 527 433
rect 475 365 527 399
rect 475 331 485 365
rect 519 331 527 365
rect 475 297 527 331
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 307 67 341 101
rect 397 63 431 97
rect 490 95 524 129
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 120 411 154 445
rect 120 343 154 377
rect 204 399 238 433
rect 290 435 324 469
rect 485 399 519 433
rect 485 331 519 365
<< poly >>
rect 79 497 109 523
rect 164 497 194 523
rect 250 497 280 523
rect 346 497 376 523
rect 445 497 475 523
rect 79 282 109 297
rect 21 249 109 282
rect 164 265 194 297
rect 250 265 280 297
rect 346 265 376 297
rect 445 265 475 297
rect 21 215 31 249
rect 65 215 109 249
rect 21 199 109 215
rect 151 249 205 265
rect 151 215 161 249
rect 195 215 205 249
rect 151 199 205 215
rect 247 249 301 265
rect 247 215 257 249
rect 291 215 301 249
rect 247 199 301 215
rect 343 249 397 265
rect 343 215 353 249
rect 387 215 397 249
rect 343 199 397 215
rect 445 249 533 265
rect 445 215 489 249
rect 523 215 533 249
rect 445 199 533 215
rect 79 177 109 199
rect 164 177 194 199
rect 250 177 280 199
rect 351 177 381 199
rect 450 177 480 199
rect 79 21 109 47
rect 164 21 194 47
rect 250 21 280 47
rect 351 21 381 47
rect 450 21 480 47
<< polycont >>
rect 31 215 65 249
rect 161 215 195 249
rect 257 215 291 249
rect 353 215 387 249
rect 489 215 523 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 19 485 85 527
rect 19 451 35 485
rect 69 451 85 485
rect 19 417 85 451
rect 19 383 35 417
rect 69 383 85 417
rect 19 349 85 383
rect 19 315 35 349
rect 69 315 85 349
rect 120 445 154 461
rect 120 377 154 411
rect 188 433 240 527
rect 188 399 204 433
rect 238 399 240 433
rect 188 383 240 399
rect 274 435 290 469
rect 324 435 340 469
rect 274 349 308 435
rect 390 401 446 471
rect 154 343 308 349
rect 120 315 308 343
rect 342 367 446 401
rect 482 433 530 467
rect 482 399 485 433
rect 519 399 530 433
rect 19 299 85 315
rect 18 249 84 265
rect 18 215 31 249
rect 65 215 84 249
rect 18 195 84 215
rect 120 249 205 265
rect 120 215 161 249
rect 195 215 205 249
rect 120 199 205 215
rect 239 249 291 265
rect 239 215 257 249
rect 239 199 291 215
rect 342 249 387 367
rect 482 365 530 399
rect 482 333 485 365
rect 342 215 353 249
rect 342 199 387 215
rect 421 331 485 333
rect 519 331 530 365
rect 421 299 530 331
rect 19 127 35 161
rect 69 127 85 161
rect 19 93 85 127
rect 19 59 35 93
rect 69 59 85 93
rect 19 17 85 59
rect 120 53 159 199
rect 239 132 273 199
rect 421 165 455 299
rect 489 249 537 265
rect 523 215 537 249
rect 489 199 537 215
rect 193 53 273 132
rect 307 131 530 165
rect 307 101 341 131
rect 481 129 530 131
rect 307 51 341 67
rect 381 63 397 97
rect 431 63 447 97
rect 381 17 447 63
rect 481 95 490 129
rect 524 95 530 129
rect 481 59 530 95
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
flabel locali s 29 221 63 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 493 85 527 119 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 491 221 525 255 0 FreeSans 200 0 0 0 C1
port 5 nsew signal input
flabel locali s 493 425 527 459 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 401 425 435 459 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 123 153 157 187 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 217 85 251 119 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 123 85 157 119 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 121 221 155 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 493 357 527 391 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel nwell s 31 527 65 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel pwell s 31 -17 65 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel metal1 s 31 527 65 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
flabel metal1 s 31 -17 65 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
rlabel comment s 0 0 0 0 4 a311oi_1
rlabel metal1 s 0 -48 644 48 1 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 644 592 1 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 644 544
string GDS_END 3726804
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3720650
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 16.100 0.000 
<< end >>
