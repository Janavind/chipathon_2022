magic
tech sky130B
magscale 1 2
timestamp 1666199351
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 54 21 641 203
rect 54 17 63 21
rect 29 -17 63 17
<< locali >>
rect 158 405 205 493
rect 350 405 419 493
rect 17 357 419 405
rect 17 177 63 357
rect 454 323 523 474
rect 97 215 163 323
rect 17 51 138 177
rect 205 51 271 323
rect 305 199 363 323
rect 397 199 523 323
rect 557 201 623 323
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 58 439 124 527
rect 242 451 308 527
rect 557 359 623 527
rect 350 125 623 165
rect 350 51 419 125
rect 457 17 523 91
rect 557 51 623 125
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel locali s 557 201 623 323 6 A1
port 1 nsew signal input
rlabel locali s 397 199 523 323 6 A2
port 2 nsew signal input
rlabel locali s 454 323 523 474 6 A2
port 2 nsew signal input
rlabel locali s 305 199 363 323 6 B1
port 3 nsew signal input
rlabel locali s 205 51 271 323 6 C1
port 4 nsew signal input
rlabel locali s 97 215 163 323 6 D1
port 5 nsew signal input
rlabel metal1 s 0 -48 644 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 17 8 VNB
port 7 nsew ground bidirectional
rlabel pwell s 54 17 63 21 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 54 21 641 203 6 VNB
port 7 nsew ground bidirectional
rlabel nwell s -38 261 682 582 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 496 644 592 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 17 51 138 177 6 Y
port 10 nsew signal output
rlabel locali s 17 177 63 357 6 Y
port 10 nsew signal output
rlabel locali s 17 357 419 405 6 Y
port 10 nsew signal output
rlabel locali s 350 405 419 493 6 Y
port 10 nsew signal output
rlabel locali s 158 405 205 493 6 Y
port 10 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 644 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 951098
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 945062
<< end >>
