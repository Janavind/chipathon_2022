magic
tech sky130A
timestamp 1666464484
<< properties >>
string GDS_END 35994136
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 35993364
<< end >>
