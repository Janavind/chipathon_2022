magic
tech sky130B
magscale 1 2
timestamp 1666464484
<< pwell >>
rect -13 -26 73 2246
rect 256 567 277 616
rect 467 -26 553 2246
<< locali >>
rect 13 0 47 2220
rect 493 0 527 2220
<< metal1 >>
rect 14 2213 526 2220
rect 14 2161 44 2213
rect 96 2161 284 2213
rect 336 2161 364 2213
rect 416 2161 444 2213
rect 496 2161 526 2213
rect 14 2154 526 2161
rect 14 126 46 2154
rect 74 66 106 2094
rect 134 126 166 2154
rect 194 66 226 2094
rect 254 126 286 2154
rect 314 66 346 2094
rect 374 126 406 2154
rect 434 66 466 2094
rect 494 126 526 2154
rect 60 59 480 66
rect 60 7 84 59
rect 136 7 164 59
rect 216 7 244 59
rect 296 7 324 59
rect 376 7 404 59
rect 456 7 480 59
rect 60 0 480 7
<< via1 >>
rect 44 2161 96 2213
rect 284 2161 336 2213
rect 364 2161 416 2213
rect 444 2161 496 2213
rect 84 7 136 59
rect 164 7 216 59
rect 244 7 296 59
rect 324 7 376 59
rect 404 7 456 59
<< metal2 >>
rect 14 2215 166 2220
rect 14 2159 42 2215
rect 98 2159 166 2215
rect 14 2154 166 2159
rect 14 126 46 2154
rect 74 66 106 2094
rect 134 126 166 2154
rect 194 66 226 2220
rect 254 2215 526 2220
rect 254 2159 282 2215
rect 338 2159 362 2215
rect 418 2159 442 2215
rect 498 2159 526 2215
rect 254 2154 526 2159
rect 254 126 286 2154
rect 314 66 346 2094
rect 374 126 406 2154
rect 434 66 466 2094
rect 494 126 526 2154
rect 60 61 480 66
rect 60 5 82 61
rect 138 5 162 61
rect 218 5 242 61
rect 298 5 322 61
rect 378 5 402 61
rect 458 5 480 61
rect 60 0 480 5
<< via2 >>
rect 42 2213 98 2215
rect 42 2161 44 2213
rect 44 2161 96 2213
rect 96 2161 98 2213
rect 42 2159 98 2161
rect 282 2213 338 2215
rect 282 2161 284 2213
rect 284 2161 336 2213
rect 336 2161 338 2213
rect 282 2159 338 2161
rect 362 2213 418 2215
rect 362 2161 364 2213
rect 364 2161 416 2213
rect 416 2161 418 2213
rect 362 2159 418 2161
rect 442 2213 498 2215
rect 442 2161 444 2213
rect 444 2161 496 2213
rect 496 2161 498 2213
rect 442 2159 498 2161
rect 82 59 138 61
rect 82 7 84 59
rect 84 7 136 59
rect 136 7 138 59
rect 82 5 138 7
rect 162 59 218 61
rect 162 7 164 59
rect 164 7 216 59
rect 216 7 218 59
rect 162 5 218 7
rect 242 59 298 61
rect 242 7 244 59
rect 244 7 296 59
rect 296 7 298 59
rect 242 5 298 7
rect 322 59 378 61
rect 322 7 324 59
rect 324 7 376 59
rect 376 7 378 59
rect 322 5 378 7
rect 402 59 458 61
rect 402 7 404 59
rect 404 7 456 59
rect 456 7 458 59
rect 402 5 458 7
<< metal3 >>
rect 0 2219 540 2220
rect 0 2155 38 2219
rect 102 2155 118 2219
rect 182 2155 198 2219
rect 262 2155 278 2219
rect 342 2155 358 2219
rect 422 2155 438 2219
rect 502 2155 540 2219
rect 0 2154 540 2155
rect 0 126 60 2154
rect 120 66 180 2094
rect 240 126 300 2154
rect 360 66 420 2094
rect 480 126 540 2154
rect 60 65 480 66
rect 60 1 78 65
rect 142 1 158 65
rect 222 1 238 65
rect 302 1 318 65
rect 382 1 398 65
rect 462 1 480 65
rect 60 0 480 1
<< via3 >>
rect 38 2215 102 2219
rect 38 2159 42 2215
rect 42 2159 98 2215
rect 98 2159 102 2215
rect 38 2155 102 2159
rect 118 2155 182 2219
rect 198 2155 262 2219
rect 278 2215 342 2219
rect 278 2159 282 2215
rect 282 2159 338 2215
rect 338 2159 342 2215
rect 278 2155 342 2159
rect 358 2215 422 2219
rect 358 2159 362 2215
rect 362 2159 418 2215
rect 418 2159 422 2215
rect 358 2155 422 2159
rect 438 2215 502 2219
rect 438 2159 442 2215
rect 442 2159 498 2215
rect 498 2159 502 2215
rect 438 2155 502 2159
rect 78 61 142 65
rect 78 5 82 61
rect 82 5 138 61
rect 138 5 142 61
rect 78 1 142 5
rect 158 61 222 65
rect 158 5 162 61
rect 162 5 218 61
rect 218 5 222 61
rect 158 1 222 5
rect 238 61 302 65
rect 238 5 242 61
rect 242 5 298 61
rect 298 5 302 61
rect 238 1 302 5
rect 318 61 382 65
rect 318 5 322 61
rect 322 5 378 61
rect 378 5 382 61
rect 318 1 382 5
rect 398 61 462 65
rect 398 5 402 61
rect 402 5 458 61
rect 458 5 462 61
rect 398 1 462 5
<< metal4 >>
rect 0 2219 540 2220
rect 0 2155 38 2219
rect 102 2155 118 2219
rect 182 2155 198 2219
rect 262 2155 278 2219
rect 342 2155 358 2219
rect 422 2155 438 2219
rect 502 2155 540 2219
rect 0 2154 540 2155
rect 0 126 60 2154
rect 120 66 180 2094
rect 240 126 300 2154
rect 360 66 420 2094
rect 480 126 540 2154
rect 60 65 480 66
rect 60 1 78 65
rect 142 1 158 65
rect 222 1 238 65
rect 302 1 318 65
rect 382 1 398 65
rect 462 1 480 65
rect 60 0 480 1
<< labels >>
flabel metal2 s 139 265 158 285 0 FreeSans 200 0 0 0 C0
port 1 nsew
flabel metal2 s 286 16 322 52 0 FreeSans 200 0 0 0 C1
port 2 nsew
flabel pwell s 256 567 277 616 0 FreeSans 400 0 0 0 SUB
port 3 nsew
<< properties >>
string GDS_END 18284
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 10556
string path 6.750 53.850 6.750 3.150 
string device primitive
<< end >>
