magic
tech sky130B
magscale 1 2
timestamp 1666464484
use sky130_fd_pr__hvdfl1sd2__example_55959141808140  sky130_fd_pr__hvdfl1sd2__example_55959141808140_0
timestamp 1666464484
transform 1 0 120 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808100  sky130_fd_pr__hvdfl1sd__example_55959141808100_0
timestamp 1666464484
transform -1 0 0 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 31674132
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 31673204
<< end >>
