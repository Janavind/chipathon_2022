magic
tech sky130B
magscale 1 2
timestamp 1666199351
<< nwell >>
rect -38 261 1142 582
<< pwell >>
rect 1 21 1060 203
rect 30 -17 64 21
<< scnmos >>
rect 83 47 113 177
rect 167 47 197 177
rect 251 47 281 177
rect 335 47 365 177
rect 525 47 555 177
rect 609 47 639 177
rect 700 47 730 177
rect 784 47 814 177
rect 868 47 898 177
rect 952 47 982 177
<< scpmoshvt >>
rect 83 297 113 497
rect 167 297 197 497
rect 251 297 281 497
rect 335 297 365 497
rect 525 297 555 497
rect 609 297 639 497
rect 700 297 730 497
rect 784 297 814 497
rect 868 297 898 497
rect 952 297 982 497
<< ndiff >>
rect 27 163 83 177
rect 27 129 39 163
rect 73 129 83 163
rect 27 95 83 129
rect 27 61 39 95
rect 73 61 83 95
rect 27 47 83 61
rect 113 163 167 177
rect 113 129 123 163
rect 157 129 167 163
rect 113 95 167 129
rect 113 61 123 95
rect 157 61 167 95
rect 113 47 167 61
rect 197 163 251 177
rect 197 129 207 163
rect 241 129 251 163
rect 197 47 251 129
rect 281 95 335 177
rect 281 61 291 95
rect 325 61 335 95
rect 281 47 335 61
rect 365 95 417 177
rect 365 61 375 95
rect 409 61 417 95
rect 365 47 417 61
rect 471 95 525 177
rect 471 61 481 95
rect 515 61 525 95
rect 471 47 525 61
rect 555 163 609 177
rect 555 129 565 163
rect 599 129 609 163
rect 555 47 609 129
rect 639 163 700 177
rect 639 129 649 163
rect 683 129 700 163
rect 639 95 700 129
rect 639 61 649 95
rect 683 61 700 95
rect 639 47 700 61
rect 730 95 784 177
rect 730 61 740 95
rect 774 61 784 95
rect 730 47 784 61
rect 814 163 868 177
rect 814 129 824 163
rect 858 129 868 163
rect 814 95 868 129
rect 814 61 824 95
rect 858 61 868 95
rect 814 47 868 61
rect 898 95 952 177
rect 898 61 908 95
rect 942 61 952 95
rect 898 47 952 61
rect 982 163 1034 177
rect 982 129 992 163
rect 1026 129 1034 163
rect 982 95 1034 129
rect 982 61 992 95
rect 1026 61 1034 95
rect 982 47 1034 61
<< pdiff >>
rect 27 477 83 497
rect 27 443 39 477
rect 73 443 83 477
rect 27 409 83 443
rect 27 375 39 409
rect 73 375 83 409
rect 27 297 83 375
rect 113 477 167 497
rect 113 443 123 477
rect 157 443 167 477
rect 113 409 167 443
rect 113 375 123 409
rect 157 375 167 409
rect 113 297 167 375
rect 197 477 251 497
rect 197 443 207 477
rect 241 443 251 477
rect 197 297 251 443
rect 281 409 335 497
rect 281 375 291 409
rect 325 375 335 409
rect 281 297 335 375
rect 365 477 525 497
rect 365 443 375 477
rect 409 443 481 477
rect 515 443 525 477
rect 365 297 525 443
rect 555 477 609 497
rect 555 443 565 477
rect 599 443 609 477
rect 555 409 609 443
rect 555 375 565 409
rect 599 375 609 409
rect 555 341 609 375
rect 555 307 565 341
rect 599 307 609 341
rect 555 297 609 307
rect 639 477 700 497
rect 639 443 649 477
rect 683 443 700 477
rect 639 297 700 443
rect 730 477 784 497
rect 730 443 740 477
rect 774 443 784 477
rect 730 297 784 443
rect 814 409 868 497
rect 814 375 824 409
rect 858 375 868 409
rect 814 297 868 375
rect 898 477 952 497
rect 898 443 908 477
rect 942 443 952 477
rect 898 409 952 443
rect 898 375 908 409
rect 942 375 952 409
rect 898 297 952 375
rect 982 477 1039 497
rect 982 443 993 477
rect 1027 443 1039 477
rect 982 409 1039 443
rect 982 375 993 409
rect 1027 375 1039 409
rect 982 297 1039 375
<< ndiffc >>
rect 39 129 73 163
rect 39 61 73 95
rect 123 129 157 163
rect 123 61 157 95
rect 207 129 241 163
rect 291 61 325 95
rect 375 61 409 95
rect 481 61 515 95
rect 565 129 599 163
rect 649 129 683 163
rect 649 61 683 95
rect 740 61 774 95
rect 824 129 858 163
rect 824 61 858 95
rect 908 61 942 95
rect 992 129 1026 163
rect 992 61 1026 95
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 123 443 157 477
rect 123 375 157 409
rect 207 443 241 477
rect 291 375 325 409
rect 375 443 409 477
rect 481 443 515 477
rect 565 443 599 477
rect 565 375 599 409
rect 565 307 599 341
rect 649 443 683 477
rect 740 443 774 477
rect 824 375 858 409
rect 908 443 942 477
rect 908 375 942 409
rect 993 443 1027 477
rect 993 375 1027 409
<< poly >>
rect 83 497 113 523
rect 167 497 197 523
rect 251 497 281 523
rect 335 497 365 523
rect 525 497 555 523
rect 609 497 639 523
rect 700 497 730 523
rect 784 497 814 523
rect 868 497 898 523
rect 952 497 982 523
rect 83 265 113 297
rect 167 265 197 297
rect 251 265 281 297
rect 335 265 365 297
rect 525 265 555 297
rect 609 265 639 297
rect 700 265 730 297
rect 784 265 814 297
rect 868 265 898 297
rect 59 249 125 265
rect 59 215 75 249
rect 109 215 125 249
rect 59 199 125 215
rect 167 249 281 265
rect 167 215 206 249
rect 240 215 281 249
rect 167 199 281 215
rect 323 249 389 265
rect 323 215 339 249
rect 373 215 389 249
rect 323 199 389 215
rect 465 249 639 265
rect 465 215 481 249
rect 515 215 639 249
rect 465 199 639 215
rect 688 249 742 265
rect 688 215 698 249
rect 732 215 742 249
rect 688 199 742 215
rect 784 249 898 265
rect 784 215 824 249
rect 858 215 898 249
rect 784 199 898 215
rect 83 177 113 199
rect 167 177 197 199
rect 251 177 281 199
rect 335 177 365 199
rect 525 177 555 199
rect 609 177 639 199
rect 700 177 730 199
rect 784 177 814 199
rect 868 177 898 199
rect 952 265 982 297
rect 952 249 1006 265
rect 952 215 962 249
rect 996 215 1006 249
rect 952 199 1006 215
rect 952 177 982 199
rect 83 21 113 47
rect 167 21 197 47
rect 251 21 281 47
rect 335 21 365 47
rect 525 21 555 47
rect 609 21 639 47
rect 700 21 730 47
rect 784 21 814 47
rect 868 21 898 47
rect 952 21 982 47
<< polycont >>
rect 75 215 109 249
rect 206 215 240 249
rect 339 215 373 249
rect 481 215 515 249
rect 698 215 732 249
rect 824 215 858 249
rect 962 215 996 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 30 477 80 527
rect 30 443 39 477
rect 73 443 80 477
rect 30 409 80 443
rect 30 375 39 409
rect 73 375 80 409
rect 30 359 80 375
rect 115 477 165 493
rect 115 443 123 477
rect 157 443 165 477
rect 115 409 165 443
rect 199 477 249 527
rect 199 443 207 477
rect 241 443 249 477
rect 199 427 249 443
rect 367 477 515 527
rect 367 443 375 477
rect 409 443 481 477
rect 367 427 515 443
rect 549 477 607 493
rect 549 443 565 477
rect 599 443 607 477
rect 115 375 123 409
rect 157 393 165 409
rect 283 409 333 425
rect 283 393 291 409
rect 157 375 291 393
rect 325 393 333 409
rect 549 409 607 443
rect 641 477 698 527
rect 641 443 649 477
rect 683 443 698 477
rect 641 425 698 443
rect 732 477 950 493
rect 732 443 740 477
rect 774 459 908 477
rect 774 443 782 459
rect 732 425 782 443
rect 900 443 908 459
rect 942 443 950 477
rect 325 375 457 393
rect 115 357 457 375
rect 18 289 389 323
rect 18 249 125 289
rect 18 215 75 249
rect 109 215 125 249
rect 159 249 280 255
rect 159 215 206 249
rect 240 215 280 249
rect 323 249 389 289
rect 323 215 339 249
rect 373 215 389 249
rect 423 265 457 357
rect 549 375 565 409
rect 599 391 607 409
rect 816 409 866 425
rect 816 391 824 409
rect 599 375 824 391
rect 858 375 866 409
rect 549 357 866 375
rect 900 409 950 443
rect 900 375 908 409
rect 942 375 950 409
rect 900 357 950 375
rect 993 477 1034 527
rect 1027 443 1034 477
rect 993 409 1034 443
rect 1027 375 1034 409
rect 993 359 1034 375
rect 549 341 643 357
rect 549 307 565 341
rect 599 307 643 341
rect 423 249 515 265
rect 423 215 481 249
rect 423 199 515 215
rect 549 215 643 307
rect 682 289 1087 323
rect 682 249 748 289
rect 682 215 698 249
rect 732 215 748 249
rect 792 249 900 255
rect 792 215 824 249
rect 858 215 900 249
rect 946 249 1087 289
rect 946 215 962 249
rect 996 215 1087 249
rect 423 181 457 199
rect 39 163 73 179
rect 39 95 73 129
rect 107 163 157 179
rect 107 129 123 163
rect 191 163 457 181
rect 191 129 207 163
rect 241 145 457 163
rect 549 163 615 215
rect 241 129 257 145
rect 549 129 565 163
rect 599 129 615 163
rect 649 163 1042 181
rect 683 147 824 163
rect 683 129 706 147
rect 107 95 157 129
rect 375 95 409 111
rect 107 61 123 95
rect 157 61 291 95
rect 325 61 341 95
rect 39 17 73 61
rect 375 17 409 61
rect 465 95 515 111
rect 649 95 706 129
rect 808 129 824 147
rect 858 145 992 163
rect 858 129 874 145
rect 465 61 481 95
rect 515 61 649 95
rect 683 61 706 95
rect 465 51 706 61
rect 740 95 774 111
rect 740 17 774 61
rect 808 95 874 129
rect 976 129 992 145
rect 1026 129 1042 163
rect 808 61 824 95
rect 858 61 874 95
rect 808 51 874 61
rect 908 95 942 111
rect 908 17 942 61
rect 976 95 1042 129
rect 976 61 992 95
rect 1026 61 1042 95
rect 976 51 1042 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
<< metal1 >>
rect 0 561 1104 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 0 496 1104 527
rect 0 17 1104 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
rect 0 -48 1104 -17
<< labels >>
flabel locali s 862 221 896 255 0 FreeSans 400 180 0 0 B2
port 4 nsew signal input
flabel locali s 586 289 620 323 0 FreeSans 400 0 0 0 Y
port 9 nsew signal output
flabel locali s 30 221 64 255 0 FreeSans 400 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 214 221 248 255 0 FreeSans 400 0 0 0 A2_N
port 2 nsew signal input
flabel locali s 1041 221 1075 255 0 FreeSans 400 180 0 0 B1
port 3 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 o2bb2ai_2
rlabel metal1 s 0 -48 1104 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1104 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1104 544
string GDS_END 1250022
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1241524
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 5.520 0.000 
<< end >>
