magic
tech sky130A
magscale 1 2
timestamp 1666199351
use sky130_fd_pr__hvdftpm1s2__example_55959141808659  sky130_fd_pr__hvdftpm1s2__example_55959141808659_0
timestamp 1666199351
transform 1 0 641 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpm1s2__example_55959141808659  sky130_fd_pr__hvdftpm1s2__example_55959141808659_1
timestamp 1666199351
transform 1 0 1633 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpm1s2__example_55959141808659  sky130_fd_pr__hvdftpm1s2__example_55959141808659_2
timestamp 1666199351
transform 1 0 2625 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpm1s2__example_55959141808659  sky130_fd_pr__hvdftpm1s2__example_55959141808659_3
timestamp 1666199351
transform 1 0 3617 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpm1s2__example_55959141808659  sky130_fd_pr__hvdftpm1s2__example_55959141808659_4
timestamp 1666199351
transform 1 0 4609 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpm1s2__example_55959141808659  sky130_fd_pr__hvdftpm1s2__example_55959141808659_5
timestamp 1666199351
transform 1 0 5601 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpm1s2__example_55959141808659  sky130_fd_pr__hvdftpm1s2__example_55959141808659_6
timestamp 1666199351
transform 1 0 6593 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpm1s2__example_55959141808659  sky130_fd_pr__hvdftpm1s2__example_55959141808659_7
timestamp 1666199351
transform 1 0 7585 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpm1s2__example_55959141808659  sky130_fd_pr__hvdftpm1s2__example_55959141808659_8
timestamp 1666199351
transform 1 0 8577 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpm1s2__example_55959141808659  sky130_fd_pr__hvdftpm1s2__example_55959141808659_9
timestamp 1666199351
transform 1 0 9569 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpm1s2__example_55959141808659  sky130_fd_pr__hvdftpm1s2__example_55959141808659_10
timestamp 1666199351
transform 1 0 10561 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpm1s2__example_55959141808659  sky130_fd_pr__hvdftpm1s2__example_55959141808659_11
timestamp 1666199351
transform 1 0 11553 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpm1s2__example_55959141808659  sky130_fd_pr__hvdftpm1s2__example_55959141808659_12
timestamp 1666199351
transform 1 0 12545 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 2366972
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 2352840
<< end >>
