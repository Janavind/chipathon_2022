magic
tech sky130B
magscale 1 2
timestamp 1666464484
<< nwell >>
rect -66 377 738 897
<< pwell >>
rect 4 43 586 283
rect -26 -43 698 43
<< mvnmos >>
rect 87 107 187 257
rect 247 107 347 257
rect 403 107 503 257
<< mvpmos >>
rect 105 443 205 743
rect 247 443 347 743
rect 403 443 503 743
<< mvndiff >>
rect 30 249 87 257
rect 30 215 42 249
rect 76 215 87 249
rect 30 149 87 215
rect 30 115 42 149
rect 76 115 87 149
rect 30 107 87 115
rect 187 167 247 257
rect 187 133 198 167
rect 232 133 247 167
rect 187 107 247 133
rect 347 249 403 257
rect 347 215 358 249
rect 392 215 403 249
rect 347 149 403 215
rect 347 115 358 149
rect 392 115 403 149
rect 347 107 403 115
rect 503 249 560 257
rect 503 215 514 249
rect 548 215 560 249
rect 503 149 560 215
rect 503 115 514 149
rect 548 115 560 149
rect 503 107 560 115
<< mvpdiff >>
rect 48 735 105 743
rect 48 701 60 735
rect 94 701 105 735
rect 48 652 105 701
rect 48 618 60 652
rect 94 618 105 652
rect 48 568 105 618
rect 48 534 60 568
rect 94 534 105 568
rect 48 485 105 534
rect 48 451 60 485
rect 94 451 105 485
rect 48 443 105 451
rect 205 443 247 743
rect 347 735 403 743
rect 347 701 358 735
rect 392 701 403 735
rect 347 652 403 701
rect 347 618 358 652
rect 392 618 403 652
rect 347 568 403 618
rect 347 534 358 568
rect 392 534 403 568
rect 347 485 403 534
rect 347 451 358 485
rect 392 451 403 485
rect 347 443 403 451
rect 503 735 560 743
rect 503 701 514 735
rect 548 701 560 735
rect 503 655 560 701
rect 503 621 514 655
rect 548 621 560 655
rect 503 574 560 621
rect 503 540 514 574
rect 548 540 560 574
rect 503 494 560 540
rect 503 460 514 494
rect 548 460 560 494
rect 503 443 560 460
<< mvndiffc >>
rect 42 215 76 249
rect 42 115 76 149
rect 198 133 232 167
rect 358 215 392 249
rect 358 115 392 149
rect 514 215 548 249
rect 514 115 548 149
<< mvpdiffc >>
rect 60 701 94 735
rect 60 618 94 652
rect 60 534 94 568
rect 60 451 94 485
rect 358 701 392 735
rect 358 618 392 652
rect 358 534 392 568
rect 358 451 392 485
rect 514 701 548 735
rect 514 621 548 655
rect 514 540 548 574
rect 514 460 548 494
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 672 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
<< poly >>
rect 105 743 205 769
rect 247 743 347 769
rect 403 743 503 769
rect 105 417 205 443
rect 87 383 205 417
rect 21 351 205 383
rect 21 317 41 351
rect 75 317 121 351
rect 155 317 205 351
rect 21 283 205 317
rect 247 343 347 443
rect 247 309 267 343
rect 301 309 347 343
rect 87 257 187 283
rect 247 257 347 309
rect 403 417 503 443
rect 403 395 535 417
rect 403 361 481 395
rect 515 361 535 395
rect 403 283 535 361
rect 403 257 503 283
rect 87 81 187 107
rect 247 81 347 107
rect 403 81 503 107
<< polycont >>
rect 41 317 75 351
rect 121 317 155 351
rect 267 309 301 343
rect 481 361 515 395
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 672 831
rect 18 735 208 751
rect 18 701 24 735
rect 58 701 60 735
rect 94 701 96 735
rect 130 701 168 735
rect 202 701 208 735
rect 18 652 208 701
rect 18 618 60 652
rect 94 618 208 652
rect 18 568 208 618
rect 18 534 60 568
rect 94 534 208 568
rect 18 485 208 534
rect 18 451 60 485
rect 94 451 208 485
rect 18 435 208 451
rect 313 735 408 751
rect 313 701 358 735
rect 392 701 408 735
rect 313 652 408 701
rect 313 618 358 652
rect 392 618 408 652
rect 313 568 408 618
rect 313 534 358 568
rect 392 534 408 568
rect 313 485 408 534
rect 313 451 358 485
rect 392 451 408 485
rect 444 735 634 751
rect 444 701 450 735
rect 484 701 514 735
rect 556 701 594 735
rect 628 701 634 735
rect 444 655 634 701
rect 444 621 514 655
rect 548 621 634 655
rect 444 574 634 621
rect 444 540 514 574
rect 548 540 634 574
rect 444 494 634 540
rect 444 460 514 494
rect 548 460 634 494
rect 313 422 408 451
rect 313 388 429 422
rect 25 351 171 367
rect 25 317 41 351
rect 75 317 121 351
rect 155 317 171 351
rect 25 301 171 317
rect 213 343 359 352
rect 213 309 267 343
rect 301 309 359 343
rect 213 301 359 309
rect 395 325 429 388
rect 465 395 647 424
rect 465 361 481 395
rect 515 361 647 395
rect 395 291 564 325
rect 26 255 92 265
rect 26 249 408 255
rect 26 215 42 249
rect 76 221 358 249
rect 76 215 92 221
rect 26 149 92 215
rect 342 215 358 221
rect 392 215 408 249
rect 26 115 42 149
rect 76 115 92 149
rect 26 99 92 115
rect 128 167 306 185
rect 128 133 198 167
rect 232 133 306 167
rect 128 113 306 133
rect 162 79 200 113
rect 234 79 272 113
rect 342 149 408 215
rect 342 115 358 149
rect 392 115 408 149
rect 342 99 408 115
rect 498 249 564 291
rect 498 215 514 249
rect 548 215 564 249
rect 498 149 564 215
rect 498 115 514 149
rect 548 115 564 149
rect 498 99 564 115
rect 128 73 306 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 24 701 58 735
rect 96 701 130 735
rect 168 701 202 735
rect 450 701 484 735
rect 522 701 548 735
rect 548 701 556 735
rect 594 701 628 735
rect 128 79 162 113
rect 200 79 234 113
rect 272 79 306 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 831 672 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 672 831
rect 0 791 672 797
rect 0 735 672 763
rect 0 701 24 735
rect 58 701 96 735
rect 130 701 168 735
rect 202 701 450 735
rect 484 701 522 735
rect 556 701 594 735
rect 628 701 672 735
rect 0 689 672 701
rect 0 113 672 125
rect 0 79 128 113
rect 162 79 200 113
rect 234 79 272 113
rect 306 79 672 113
rect 0 51 672 79
rect 0 17 672 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -23 672 -17
<< labels >>
rlabel comment s 0 0 0 0 4 o21ai_1
flabel metal1 s 0 51 672 125 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 0 0 672 23 0 FreeSans 340 0 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 0 689 672 763 0 FreeSans 340 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 791 672 814 0 FreeSans 340 0 0 0 VPB
port 6 nsew power bidirectional
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 319 464 353 498 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 319 538 353 572 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
flabel locali s 319 612 353 646 0 FreeSans 340 0 0 0 Y
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 672 814
string GDS_END 407940
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 398986
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
<< end >>
