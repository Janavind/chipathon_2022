magic
tech sky130B
magscale 1 2
timestamp 1666464484
<< dnwell >>
rect 16073 -8402 21019 -6652
rect 16073 -11421 20759 -8402
<< nwell >>
rect 15993 -6858 21099 -6572
rect 15993 -10351 16279 -6858
rect 18191 -8459 18262 -8079
rect 20813 -8196 21099 -6858
rect 20553 -8482 21099 -8196
rect 20553 -9772 20839 -8482
rect 15993 -10783 16404 -10351
rect 17657 -10665 18843 -9868
rect 20104 -10204 20176 -9872
rect 20514 -10204 20839 -9772
rect 15993 -11215 16279 -10783
rect 20553 -11215 20839 -10204
rect 22343 -10544 23737 -10378
rect 15993 -11501 20839 -11215
rect 22486 -12089 24604 -11923
<< pwell >>
rect 18322 -9193 19422 -9107
rect 18735 -9535 19149 -9193
rect 20148 -9283 20492 -8079
rect 19441 -9377 20492 -9283
rect 19441 -9535 20122 -9377
rect 17166 -10320 17518 -10127
rect 16959 -10522 17518 -10320
rect 17166 -10541 17518 -10522
rect 22409 -11492 26270 -11406
<< mvnmos >>
rect 18814 -9509 18914 -9309
rect 18970 -9509 19070 -9309
rect 19520 -9509 19620 -9309
rect 19676 -9509 19776 -9309
rect 19943 -9509 20043 -9309
rect 17192 -10306 17492 -10206
rect 17192 -10462 17492 -10362
<< mvpmos >>
rect 17857 -10530 18257 -10380
rect 18313 -10530 18713 -10380
<< mvndiff >>
rect 18761 -9321 18814 -9309
rect 18761 -9355 18769 -9321
rect 18803 -9355 18814 -9321
rect 18761 -9389 18814 -9355
rect 18761 -9423 18769 -9389
rect 18803 -9423 18814 -9389
rect 18761 -9457 18814 -9423
rect 18761 -9491 18769 -9457
rect 18803 -9491 18814 -9457
rect 18761 -9509 18814 -9491
rect 18914 -9321 18970 -9309
rect 18914 -9355 18925 -9321
rect 18959 -9355 18970 -9321
rect 18914 -9389 18970 -9355
rect 18914 -9423 18925 -9389
rect 18959 -9423 18970 -9389
rect 18914 -9457 18970 -9423
rect 18914 -9491 18925 -9457
rect 18959 -9491 18970 -9457
rect 18914 -9509 18970 -9491
rect 19070 -9321 19123 -9309
rect 19070 -9355 19081 -9321
rect 19115 -9355 19123 -9321
rect 19070 -9389 19123 -9355
rect 19070 -9423 19081 -9389
rect 19115 -9423 19123 -9389
rect 19070 -9457 19123 -9423
rect 19070 -9491 19081 -9457
rect 19115 -9491 19123 -9457
rect 19070 -9509 19123 -9491
rect 19467 -9327 19520 -9309
rect 19467 -9361 19475 -9327
rect 19509 -9361 19520 -9327
rect 19467 -9395 19520 -9361
rect 19467 -9429 19475 -9395
rect 19509 -9429 19520 -9395
rect 19467 -9463 19520 -9429
rect 19467 -9497 19475 -9463
rect 19509 -9497 19520 -9463
rect 19467 -9509 19520 -9497
rect 19620 -9327 19676 -9309
rect 19620 -9361 19631 -9327
rect 19665 -9361 19676 -9327
rect 19620 -9395 19676 -9361
rect 19620 -9429 19631 -9395
rect 19665 -9429 19676 -9395
rect 19620 -9463 19676 -9429
rect 19620 -9497 19631 -9463
rect 19665 -9497 19676 -9463
rect 19620 -9509 19676 -9497
rect 19776 -9327 19829 -9309
rect 19776 -9361 19787 -9327
rect 19821 -9361 19829 -9327
rect 19776 -9395 19829 -9361
rect 19776 -9429 19787 -9395
rect 19821 -9429 19829 -9395
rect 19776 -9463 19829 -9429
rect 19776 -9497 19787 -9463
rect 19821 -9497 19829 -9463
rect 19776 -9509 19829 -9497
rect 19890 -9327 19943 -9309
rect 19890 -9361 19898 -9327
rect 19932 -9361 19943 -9327
rect 19890 -9395 19943 -9361
rect 19890 -9429 19898 -9395
rect 19932 -9429 19943 -9395
rect 19890 -9463 19943 -9429
rect 19890 -9497 19898 -9463
rect 19932 -9497 19943 -9463
rect 19890 -9509 19943 -9497
rect 20043 -9327 20096 -9309
rect 20043 -9361 20054 -9327
rect 20088 -9361 20096 -9327
rect 20043 -9395 20096 -9361
rect 20043 -9429 20054 -9395
rect 20088 -9429 20096 -9395
rect 20043 -9463 20096 -9429
rect 20043 -9497 20054 -9463
rect 20088 -9497 20096 -9463
rect 20043 -9509 20096 -9497
rect 17192 -10161 17492 -10153
rect 17192 -10195 17242 -10161
rect 17276 -10195 17310 -10161
rect 17344 -10195 17378 -10161
rect 17412 -10195 17446 -10161
rect 17480 -10195 17492 -10161
rect 17192 -10206 17492 -10195
rect 17192 -10317 17492 -10306
rect 17192 -10351 17242 -10317
rect 17276 -10351 17310 -10317
rect 17344 -10351 17378 -10317
rect 17412 -10351 17446 -10317
rect 17480 -10351 17492 -10317
rect 17192 -10362 17492 -10351
rect 17192 -10473 17492 -10462
rect 17192 -10507 17242 -10473
rect 17276 -10507 17310 -10473
rect 17344 -10507 17378 -10473
rect 17412 -10507 17446 -10473
rect 17480 -10507 17492 -10473
rect 17192 -10515 17492 -10507
<< mvpdiff >>
rect 17804 -10416 17857 -10380
rect 17804 -10450 17812 -10416
rect 17846 -10450 17857 -10416
rect 17804 -10484 17857 -10450
rect 17804 -10518 17812 -10484
rect 17846 -10518 17857 -10484
rect 17804 -10530 17857 -10518
rect 18257 -10416 18313 -10380
rect 18257 -10450 18268 -10416
rect 18302 -10450 18313 -10416
rect 18257 -10484 18313 -10450
rect 18257 -10518 18268 -10484
rect 18302 -10518 18313 -10484
rect 18257 -10530 18313 -10518
rect 18713 -10416 18766 -10380
rect 18713 -10450 18724 -10416
rect 18758 -10450 18766 -10416
rect 18713 -10484 18766 -10450
rect 18713 -10518 18724 -10484
rect 18758 -10518 18766 -10484
rect 18713 -10530 18766 -10518
<< mvndiffc >>
rect 18769 -9355 18803 -9321
rect 18769 -9423 18803 -9389
rect 18769 -9491 18803 -9457
rect 18925 -9355 18959 -9321
rect 18925 -9423 18959 -9389
rect 18925 -9491 18959 -9457
rect 19081 -9355 19115 -9321
rect 19081 -9423 19115 -9389
rect 19081 -9491 19115 -9457
rect 19475 -9361 19509 -9327
rect 19475 -9429 19509 -9395
rect 19475 -9497 19509 -9463
rect 19631 -9361 19665 -9327
rect 19631 -9429 19665 -9395
rect 19631 -9497 19665 -9463
rect 19787 -9361 19821 -9327
rect 19787 -9429 19821 -9395
rect 19787 -9497 19821 -9463
rect 19898 -9361 19932 -9327
rect 19898 -9429 19932 -9395
rect 19898 -9497 19932 -9463
rect 20054 -9361 20088 -9327
rect 20054 -9429 20088 -9395
rect 20054 -9497 20088 -9463
rect 17242 -10195 17276 -10161
rect 17310 -10195 17344 -10161
rect 17378 -10195 17412 -10161
rect 17446 -10195 17480 -10161
rect 17242 -10351 17276 -10317
rect 17310 -10351 17344 -10317
rect 17378 -10351 17412 -10317
rect 17446 -10351 17480 -10317
rect 17242 -10507 17276 -10473
rect 17310 -10507 17344 -10473
rect 17378 -10507 17412 -10473
rect 17446 -10507 17480 -10473
<< mvpdiffc >>
rect 17812 -10450 17846 -10416
rect 17812 -10518 17846 -10484
rect 18268 -10450 18302 -10416
rect 18268 -10518 18302 -10484
rect 18724 -10450 18758 -10416
rect 18724 -10518 18758 -10484
<< psubdiff >>
rect 23669 -11466 23702 -11432
rect 23736 -11466 23771 -11432
rect 23805 -11466 23840 -11432
rect 23874 -11466 23909 -11432
rect 23943 -11466 23978 -11432
rect 24012 -11466 24047 -11432
rect 24081 -11466 24116 -11432
rect 24150 -11466 24185 -11432
rect 24219 -11466 24254 -11432
rect 24288 -11466 24323 -11432
rect 24357 -11466 24392 -11432
rect 24426 -11466 24461 -11432
rect 24495 -11466 24530 -11432
rect 24564 -11466 24599 -11432
rect 24633 -11466 24668 -11432
rect 24702 -11466 24737 -11432
rect 24771 -11466 24806 -11432
rect 24840 -11466 24875 -11432
rect 24909 -11466 24944 -11432
rect 24978 -11466 25013 -11432
rect 25047 -11466 25082 -11432
rect 25116 -11466 25151 -11432
rect 25185 -11466 25220 -11432
rect 25254 -11466 25289 -11432
rect 25323 -11466 25358 -11432
rect 25392 -11466 25427 -11432
rect 25461 -11466 25496 -11432
rect 25530 -11466 25565 -11432
rect 25599 -11466 25634 -11432
rect 25668 -11466 25703 -11432
rect 25737 -11466 25772 -11432
rect 25806 -11466 25841 -11432
rect 25875 -11466 25910 -11432
rect 25944 -11466 25979 -11432
rect 26013 -11466 26048 -11432
rect 26082 -11466 26117 -11432
rect 26151 -11466 26186 -11432
rect 26220 -11466 26244 -11432
<< mvpsubdiff >>
rect 20174 -8139 20466 -8105
rect 20208 -8173 20260 -8139
rect 20294 -8173 20346 -8139
rect 20380 -8173 20432 -8139
rect 20174 -8210 20466 -8173
rect 20208 -8244 20260 -8210
rect 20294 -8244 20346 -8210
rect 20380 -8244 20432 -8210
rect 20174 -8281 20466 -8244
rect 20208 -8315 20260 -8281
rect 20294 -8315 20346 -8281
rect 20380 -8315 20432 -8281
rect 20174 -8352 20466 -8315
rect 20208 -8386 20260 -8352
rect 20294 -8386 20346 -8352
rect 20380 -8386 20432 -8352
rect 20174 -8423 20466 -8386
rect 20208 -8457 20260 -8423
rect 20294 -8457 20346 -8423
rect 20380 -8457 20432 -8423
rect 20174 -8494 20466 -8457
rect 20208 -8528 20260 -8494
rect 20294 -8528 20346 -8494
rect 20380 -8528 20432 -8494
rect 20174 -8565 20466 -8528
rect 20208 -8599 20260 -8565
rect 20294 -8599 20346 -8565
rect 20380 -8599 20432 -8565
rect 20174 -8636 20466 -8599
rect 20208 -8670 20260 -8636
rect 20294 -8670 20346 -8636
rect 20380 -8670 20432 -8636
rect 20174 -8707 20466 -8670
rect 20208 -8741 20260 -8707
rect 20294 -8741 20346 -8707
rect 20380 -8741 20432 -8707
rect 20174 -8779 20466 -8741
rect 20208 -8813 20260 -8779
rect 20294 -8813 20346 -8779
rect 20380 -8813 20432 -8779
rect 20174 -8851 20466 -8813
rect 20208 -8885 20260 -8851
rect 20294 -8885 20346 -8851
rect 20380 -8885 20432 -8851
rect 20174 -8923 20466 -8885
rect 20208 -8957 20260 -8923
rect 20294 -8957 20346 -8923
rect 20380 -8957 20432 -8923
rect 20174 -8995 20466 -8957
rect 20208 -9029 20260 -8995
rect 20294 -9029 20346 -8995
rect 20380 -9029 20432 -8995
rect 20174 -9067 20466 -9029
rect 20208 -9101 20260 -9067
rect 20294 -9101 20346 -9067
rect 20380 -9101 20432 -9067
rect 18348 -9167 18372 -9133
rect 18406 -9167 18441 -9133
rect 18475 -9167 18510 -9133
rect 18544 -9167 18579 -9133
rect 18613 -9167 18648 -9133
rect 18682 -9167 18717 -9133
rect 18751 -9167 18786 -9133
rect 18820 -9167 18855 -9133
rect 18889 -9167 18924 -9133
rect 18958 -9167 18993 -9133
rect 19027 -9167 19062 -9133
rect 19096 -9167 19131 -9133
rect 19165 -9167 19200 -9133
rect 19234 -9167 19269 -9133
rect 19303 -9167 19338 -9133
rect 19372 -9167 19396 -9133
rect 20174 -9139 20466 -9101
rect 20208 -9173 20260 -9139
rect 20294 -9173 20346 -9139
rect 20380 -9173 20432 -9139
rect 20174 -9211 20466 -9173
rect 20208 -9245 20260 -9211
rect 20294 -9245 20346 -9211
rect 20380 -9245 20432 -9211
rect 20174 -9283 20466 -9245
rect 20208 -9317 20260 -9283
rect 20294 -9317 20346 -9283
rect 20380 -9317 20432 -9283
rect 20174 -9351 20466 -9317
rect 16985 -10370 17101 -10346
rect 17019 -10404 17067 -10370
rect 16985 -10438 17101 -10404
rect 17019 -10472 17067 -10438
rect 16985 -10496 17101 -10472
rect 22435 -11466 22459 -11432
rect 22493 -11466 22529 -11432
rect 22563 -11466 22598 -11432
rect 22632 -11466 22667 -11432
rect 22701 -11466 22736 -11432
rect 22770 -11466 22805 -11432
rect 22839 -11466 22874 -11432
rect 22908 -11466 22943 -11432
rect 22977 -11466 23012 -11432
rect 23046 -11466 23081 -11432
rect 23115 -11466 23150 -11432
rect 23184 -11466 23219 -11432
rect 23253 -11466 23288 -11432
rect 23322 -11466 23357 -11432
rect 23391 -11466 23426 -11432
rect 23460 -11466 23495 -11432
rect 23529 -11466 23564 -11432
rect 23598 -11466 23633 -11432
rect 23667 -11466 23669 -11432
<< mvnsubdiff >>
rect 16119 -6732 16247 -6698
rect 16281 -6732 16315 -6698
rect 16349 -6732 16383 -6698
rect 16417 -6732 16451 -6698
rect 16485 -6732 16519 -6698
rect 16553 -6732 16587 -6698
rect 16621 -6732 16655 -6698
rect 16689 -6732 16723 -6698
rect 16757 -6732 16791 -6698
rect 16825 -6732 16859 -6698
rect 16893 -6732 16927 -6698
rect 16961 -6732 16995 -6698
rect 17029 -6732 17063 -6698
rect 17097 -6732 17131 -6698
rect 17165 -6732 17199 -6698
rect 17233 -6732 17267 -6698
rect 17301 -6732 17335 -6698
rect 17369 -6732 17403 -6698
rect 17437 -6732 17471 -6698
rect 17505 -6732 17539 -6698
rect 17573 -6732 17607 -6698
rect 17641 -6732 17675 -6698
rect 17709 -6732 17743 -6698
rect 17777 -6732 17811 -6698
rect 17845 -6732 17879 -6698
rect 17913 -6732 17947 -6698
rect 17981 -6732 18015 -6698
rect 18049 -6732 18083 -6698
rect 18117 -6732 18151 -6698
rect 18185 -6732 18219 -6698
rect 18253 -6732 18287 -6698
rect 18321 -6732 18355 -6698
rect 18389 -6732 18423 -6698
rect 18457 -6732 18491 -6698
rect 18525 -6732 18559 -6698
rect 18593 -6732 18627 -6698
rect 18661 -6732 18695 -6698
rect 18729 -6732 18763 -6698
rect 18797 -6732 18831 -6698
rect 18865 -6732 18899 -6698
rect 18933 -6732 18967 -6698
rect 19001 -6732 19035 -6698
rect 19069 -6732 19103 -6698
rect 19137 -6732 19171 -6698
rect 19205 -6732 19239 -6698
rect 19273 -6732 19307 -6698
rect 19341 -6732 19375 -6698
rect 19409 -6732 19443 -6698
rect 19477 -6732 19511 -6698
rect 19545 -6732 19579 -6698
rect 19613 -6732 19647 -6698
rect 19681 -6732 19715 -6698
rect 19749 -6732 19783 -6698
rect 19817 -6732 19851 -6698
rect 19885 -6732 19919 -6698
rect 19953 -6732 19987 -6698
rect 20021 -6732 20055 -6698
rect 20089 -6732 20123 -6698
rect 20157 -6732 20191 -6698
rect 20225 -6732 20259 -6698
rect 20293 -6732 20327 -6698
rect 20361 -6732 20395 -6698
rect 20429 -6732 20463 -6698
rect 20497 -6732 20531 -6698
rect 20565 -6732 20599 -6698
rect 20633 -6732 20667 -6698
rect 20701 -6732 20735 -6698
rect 20769 -6732 20803 -6698
rect 20837 -6732 20871 -6698
rect 20905 -6732 20973 -6698
rect 16119 -6766 16153 -6732
rect 16119 -6834 16153 -6800
rect 16119 -6902 16153 -6868
rect 16119 -6970 16153 -6936
rect 16119 -7038 16153 -7004
rect 16119 -7106 16153 -7072
rect 16119 -7174 16153 -7140
rect 16119 -7242 16153 -7208
rect 16119 -7310 16153 -7276
rect 16119 -7378 16153 -7344
rect 16119 -7446 16153 -7412
rect 16119 -7514 16153 -7480
rect 16119 -7582 16153 -7548
rect 16119 -7650 16153 -7616
rect 16119 -7718 16153 -7684
rect 16119 -7786 16153 -7752
rect 16119 -7854 16153 -7820
rect 16119 -7922 16153 -7888
rect 16119 -7990 16153 -7956
rect 16119 -8058 16153 -8024
rect 16119 -8126 16153 -8092
rect 20939 -6826 20973 -6732
rect 20939 -6894 20973 -6860
rect 20939 -6962 20973 -6928
rect 20939 -7030 20973 -6996
rect 20939 -7098 20973 -7064
rect 20939 -7166 20973 -7132
rect 20939 -7234 20973 -7200
rect 20939 -7302 20973 -7268
rect 20939 -7370 20973 -7336
rect 20939 -7438 20973 -7404
rect 20939 -7506 20973 -7472
rect 20939 -7574 20973 -7540
rect 20939 -7642 20973 -7608
rect 20939 -7710 20973 -7676
rect 20939 -7778 20973 -7744
rect 20939 -7846 20973 -7812
rect 20939 -7914 20973 -7880
rect 20939 -7982 20973 -7948
rect 20939 -8050 20973 -8016
rect 16119 -8194 16153 -8160
rect 16119 -8262 16153 -8228
rect 16119 -8330 16153 -8296
rect 16119 -8398 16153 -8364
rect 16119 -8466 16153 -8432
rect 16119 -8534 16153 -8500
rect 16119 -8602 16153 -8568
rect 16119 -8670 16153 -8636
rect 16119 -8738 16153 -8704
rect 16119 -8806 16153 -8772
rect 16119 -8874 16153 -8840
rect 16119 -8942 16153 -8908
rect 16119 -9010 16153 -8976
rect 16119 -9078 16153 -9044
rect 16119 -9146 16153 -9112
rect 20939 -8118 20973 -8084
rect 20939 -8186 20973 -8152
rect 20939 -8254 20973 -8220
rect 20939 -8322 20973 -8288
rect 16119 -9214 16153 -9180
rect 16119 -9282 16153 -9248
rect 16119 -9350 16153 -9316
rect 16119 -9418 16153 -9384
rect 16119 -9486 16153 -9452
rect 20679 -8356 20747 -8322
rect 20781 -8356 20815 -8322
rect 20849 -8356 20973 -8322
rect 20679 -8417 20713 -8356
rect 20679 -8485 20713 -8451
rect 20679 -8553 20713 -8519
rect 20679 -8621 20713 -8587
rect 20679 -8689 20713 -8655
rect 20679 -8757 20713 -8723
rect 20679 -8825 20713 -8791
rect 20679 -8893 20713 -8859
rect 20679 -8961 20713 -8927
rect 20679 -9029 20713 -8995
rect 20679 -9097 20713 -9063
rect 20679 -9165 20713 -9131
rect 20679 -9233 20713 -9199
rect 20679 -9301 20713 -9267
rect 20679 -9369 20713 -9335
rect 20679 -9437 20713 -9403
rect 20679 -9505 20713 -9471
rect 16119 -9554 16153 -9520
rect 16119 -9622 16153 -9588
rect 16119 -9690 16153 -9656
rect 16119 -9758 16153 -9724
rect 16119 -9902 16153 -9792
rect 16119 -9970 16153 -9936
rect 20679 -9573 20713 -9539
rect 20679 -9641 20713 -9607
rect 20679 -9709 20713 -9675
rect 20679 -9777 20713 -9743
rect 20679 -9845 20713 -9811
rect 20679 -9913 20713 -9879
rect 16119 -10038 16153 -10004
rect 16119 -10106 16153 -10072
rect 16119 -10174 16153 -10140
rect 18349 -9962 18383 -9938
rect 18349 -10097 18383 -9996
rect 18349 -10155 18383 -10131
rect 20679 -9981 20713 -9947
rect 20679 -10049 20713 -10015
rect 20679 -10117 20713 -10083
rect 20679 -10185 20713 -10151
rect 16119 -10242 16153 -10208
rect 16119 -10310 16153 -10276
rect 20679 -10253 20713 -10219
rect 16119 -10378 16153 -10344
rect 16119 -10446 16153 -10412
rect 16119 -10514 16153 -10480
rect 20679 -10321 20713 -10287
rect 20679 -10389 20713 -10355
rect 20679 -10457 20713 -10423
rect 22409 -10478 22443 -10444
rect 22477 -10478 22588 -10444
rect 22622 -10478 22733 -10444
rect 22767 -10478 22878 -10444
rect 22912 -10478 23023 -10444
rect 23057 -10478 23168 -10444
rect 23202 -10478 23313 -10444
rect 23347 -10478 23458 -10444
rect 23492 -10478 23603 -10444
rect 23637 -10478 23671 -10444
rect 20679 -10525 20713 -10491
rect 16119 -10582 16153 -10548
rect 16119 -10650 16153 -10616
rect 20679 -10593 20713 -10559
rect 16119 -10718 16153 -10684
rect 16119 -10786 16153 -10752
rect 16119 -10854 16153 -10820
rect 16119 -10922 16153 -10888
rect 16119 -10990 16153 -10956
rect 16119 -11058 16153 -11024
rect 16119 -11126 16153 -11092
rect 16119 -11194 16153 -11160
rect 16119 -11262 16153 -11228
rect 16119 -11341 16153 -11296
rect 20679 -10661 20713 -10627
rect 20679 -10729 20713 -10695
rect 20679 -10797 20713 -10763
rect 20679 -10865 20713 -10831
rect 20679 -10933 20713 -10899
rect 20679 -11001 20713 -10967
rect 20679 -11069 20713 -11035
rect 20679 -11137 20713 -11103
rect 20679 -11205 20713 -11171
rect 20679 -11273 20713 -11239
rect 20679 -11341 20713 -11307
rect 16119 -11375 16187 -11341
rect 16221 -11375 16255 -11341
rect 16289 -11375 16323 -11341
rect 16357 -11375 16391 -11341
rect 16425 -11375 16459 -11341
rect 16493 -11375 16527 -11341
rect 16561 -11375 16595 -11341
rect 16629 -11375 16663 -11341
rect 16697 -11375 16731 -11341
rect 16765 -11375 16799 -11341
rect 16833 -11375 16867 -11341
rect 16901 -11375 16935 -11341
rect 16969 -11375 17003 -11341
rect 17037 -11375 17071 -11341
rect 17105 -11375 17139 -11341
rect 17173 -11375 17207 -11341
rect 17241 -11375 17275 -11341
rect 17309 -11375 17343 -11341
rect 17377 -11375 17411 -11341
rect 17445 -11375 17479 -11341
rect 17513 -11375 17547 -11341
rect 17581 -11375 17615 -11341
rect 17649 -11375 17683 -11341
rect 17717 -11375 17751 -11341
rect 17785 -11375 17819 -11341
rect 17853 -11375 17887 -11341
rect 17921 -11375 17955 -11341
rect 17989 -11375 18023 -11341
rect 18057 -11375 18091 -11341
rect 18125 -11375 18159 -11341
rect 18193 -11375 18227 -11341
rect 18261 -11375 18295 -11341
rect 18329 -11375 18363 -11341
rect 18397 -11375 18431 -11341
rect 18465 -11375 18499 -11341
rect 18533 -11375 18567 -11341
rect 18601 -11375 18635 -11341
rect 18669 -11375 18703 -11341
rect 18737 -11375 18771 -11341
rect 18805 -11375 18839 -11341
rect 18873 -11375 18907 -11341
rect 18941 -11375 18975 -11341
rect 19009 -11375 19043 -11341
rect 19077 -11375 19111 -11341
rect 19145 -11375 19179 -11341
rect 19213 -11375 19247 -11341
rect 19281 -11375 19315 -11341
rect 19349 -11375 19383 -11341
rect 19417 -11375 19451 -11341
rect 19485 -11375 19519 -11341
rect 19553 -11375 19587 -11341
rect 19621 -11375 19655 -11341
rect 19689 -11375 19723 -11341
rect 19757 -11375 19791 -11341
rect 19825 -11375 19859 -11341
rect 19893 -11375 19927 -11341
rect 19961 -11375 19995 -11341
rect 20029 -11375 20063 -11341
rect 20097 -11375 20131 -11341
rect 20165 -11375 20199 -11341
rect 20233 -11375 20267 -11341
rect 20301 -11375 20335 -11341
rect 20369 -11375 20403 -11341
rect 20437 -11375 20471 -11341
rect 20505 -11375 20539 -11341
rect 20573 -11375 20607 -11341
rect 20641 -11375 20713 -11341
rect 22552 -12023 22576 -11989
rect 22610 -12023 22644 -11989
rect 22678 -12023 22712 -11989
rect 22746 -12023 22780 -11989
rect 22814 -12023 22848 -11989
rect 22882 -12023 22916 -11989
rect 22950 -12023 22984 -11989
rect 23018 -12023 23052 -11989
rect 23086 -12023 23120 -11989
rect 23154 -12023 23188 -11989
rect 23222 -12023 23256 -11989
rect 23290 -12023 23324 -11989
rect 23358 -12023 23392 -11989
rect 23426 -12023 23460 -11989
rect 23494 -12023 23528 -11989
rect 23562 -12023 23596 -11989
rect 23630 -12023 23664 -11989
rect 23698 -12023 23732 -11989
rect 23766 -12023 23800 -11989
rect 23834 -12023 23868 -11989
rect 23902 -12023 23936 -11989
rect 23970 -12023 24004 -11989
rect 24038 -12023 24072 -11989
rect 24106 -12023 24140 -11989
rect 24174 -12023 24208 -11989
rect 24242 -12023 24276 -11989
rect 24310 -12023 24344 -11989
rect 24378 -12023 24412 -11989
rect 24446 -12023 24480 -11989
rect 24514 -12023 24538 -11989
<< psubdiffcont >>
rect 23702 -11466 23736 -11432
rect 23771 -11466 23805 -11432
rect 23840 -11466 23874 -11432
rect 23909 -11466 23943 -11432
rect 23978 -11466 24012 -11432
rect 24047 -11466 24081 -11432
rect 24116 -11466 24150 -11432
rect 24185 -11466 24219 -11432
rect 24254 -11466 24288 -11432
rect 24323 -11466 24357 -11432
rect 24392 -11466 24426 -11432
rect 24461 -11466 24495 -11432
rect 24530 -11466 24564 -11432
rect 24599 -11466 24633 -11432
rect 24668 -11466 24702 -11432
rect 24737 -11466 24771 -11432
rect 24806 -11466 24840 -11432
rect 24875 -11466 24909 -11432
rect 24944 -11466 24978 -11432
rect 25013 -11466 25047 -11432
rect 25082 -11466 25116 -11432
rect 25151 -11466 25185 -11432
rect 25220 -11466 25254 -11432
rect 25289 -11466 25323 -11432
rect 25358 -11466 25392 -11432
rect 25427 -11466 25461 -11432
rect 25496 -11466 25530 -11432
rect 25565 -11466 25599 -11432
rect 25634 -11466 25668 -11432
rect 25703 -11466 25737 -11432
rect 25772 -11466 25806 -11432
rect 25841 -11466 25875 -11432
rect 25910 -11466 25944 -11432
rect 25979 -11466 26013 -11432
rect 26048 -11466 26082 -11432
rect 26117 -11466 26151 -11432
rect 26186 -11466 26220 -11432
<< mvpsubdiffcont >>
rect 20174 -8173 20208 -8139
rect 20260 -8173 20294 -8139
rect 20346 -8173 20380 -8139
rect 20432 -8173 20466 -8139
rect 20174 -8244 20208 -8210
rect 20260 -8244 20294 -8210
rect 20346 -8244 20380 -8210
rect 20432 -8244 20466 -8210
rect 20174 -8315 20208 -8281
rect 20260 -8315 20294 -8281
rect 20346 -8315 20380 -8281
rect 20432 -8315 20466 -8281
rect 20174 -8386 20208 -8352
rect 20260 -8386 20294 -8352
rect 20346 -8386 20380 -8352
rect 20432 -8386 20466 -8352
rect 20174 -8457 20208 -8423
rect 20260 -8457 20294 -8423
rect 20346 -8457 20380 -8423
rect 20432 -8457 20466 -8423
rect 20174 -8528 20208 -8494
rect 20260 -8528 20294 -8494
rect 20346 -8528 20380 -8494
rect 20432 -8528 20466 -8494
rect 20174 -8599 20208 -8565
rect 20260 -8599 20294 -8565
rect 20346 -8599 20380 -8565
rect 20432 -8599 20466 -8565
rect 20174 -8670 20208 -8636
rect 20260 -8670 20294 -8636
rect 20346 -8670 20380 -8636
rect 20432 -8670 20466 -8636
rect 20174 -8741 20208 -8707
rect 20260 -8741 20294 -8707
rect 20346 -8741 20380 -8707
rect 20432 -8741 20466 -8707
rect 20174 -8813 20208 -8779
rect 20260 -8813 20294 -8779
rect 20346 -8813 20380 -8779
rect 20432 -8813 20466 -8779
rect 20174 -8885 20208 -8851
rect 20260 -8885 20294 -8851
rect 20346 -8885 20380 -8851
rect 20432 -8885 20466 -8851
rect 20174 -8957 20208 -8923
rect 20260 -8957 20294 -8923
rect 20346 -8957 20380 -8923
rect 20432 -8957 20466 -8923
rect 20174 -9029 20208 -8995
rect 20260 -9029 20294 -8995
rect 20346 -9029 20380 -8995
rect 20432 -9029 20466 -8995
rect 20174 -9101 20208 -9067
rect 20260 -9101 20294 -9067
rect 20346 -9101 20380 -9067
rect 20432 -9101 20466 -9067
rect 18372 -9167 18406 -9133
rect 18441 -9167 18475 -9133
rect 18510 -9167 18544 -9133
rect 18579 -9167 18613 -9133
rect 18648 -9167 18682 -9133
rect 18717 -9167 18751 -9133
rect 18786 -9167 18820 -9133
rect 18855 -9167 18889 -9133
rect 18924 -9167 18958 -9133
rect 18993 -9167 19027 -9133
rect 19062 -9167 19096 -9133
rect 19131 -9167 19165 -9133
rect 19200 -9167 19234 -9133
rect 19269 -9167 19303 -9133
rect 19338 -9167 19372 -9133
rect 20174 -9173 20208 -9139
rect 20260 -9173 20294 -9139
rect 20346 -9173 20380 -9139
rect 20432 -9173 20466 -9139
rect 20174 -9245 20208 -9211
rect 20260 -9245 20294 -9211
rect 20346 -9245 20380 -9211
rect 20432 -9245 20466 -9211
rect 20174 -9317 20208 -9283
rect 20260 -9317 20294 -9283
rect 20346 -9317 20380 -9283
rect 20432 -9317 20466 -9283
rect 16985 -10404 17019 -10370
rect 17067 -10404 17101 -10370
rect 16985 -10472 17019 -10438
rect 17067 -10472 17101 -10438
rect 22459 -11466 22493 -11432
rect 22529 -11466 22563 -11432
rect 22598 -11466 22632 -11432
rect 22667 -11466 22701 -11432
rect 22736 -11466 22770 -11432
rect 22805 -11466 22839 -11432
rect 22874 -11466 22908 -11432
rect 22943 -11466 22977 -11432
rect 23012 -11466 23046 -11432
rect 23081 -11466 23115 -11432
rect 23150 -11466 23184 -11432
rect 23219 -11466 23253 -11432
rect 23288 -11466 23322 -11432
rect 23357 -11466 23391 -11432
rect 23426 -11466 23460 -11432
rect 23495 -11466 23529 -11432
rect 23564 -11466 23598 -11432
rect 23633 -11466 23667 -11432
<< mvnsubdiffcont >>
rect 16247 -6732 16281 -6698
rect 16315 -6732 16349 -6698
rect 16383 -6732 16417 -6698
rect 16451 -6732 16485 -6698
rect 16519 -6732 16553 -6698
rect 16587 -6732 16621 -6698
rect 16655 -6732 16689 -6698
rect 16723 -6732 16757 -6698
rect 16791 -6732 16825 -6698
rect 16859 -6732 16893 -6698
rect 16927 -6732 16961 -6698
rect 16995 -6732 17029 -6698
rect 17063 -6732 17097 -6698
rect 17131 -6732 17165 -6698
rect 17199 -6732 17233 -6698
rect 17267 -6732 17301 -6698
rect 17335 -6732 17369 -6698
rect 17403 -6732 17437 -6698
rect 17471 -6732 17505 -6698
rect 17539 -6732 17573 -6698
rect 17607 -6732 17641 -6698
rect 17675 -6732 17709 -6698
rect 17743 -6732 17777 -6698
rect 17811 -6732 17845 -6698
rect 17879 -6732 17913 -6698
rect 17947 -6732 17981 -6698
rect 18015 -6732 18049 -6698
rect 18083 -6732 18117 -6698
rect 18151 -6732 18185 -6698
rect 18219 -6732 18253 -6698
rect 18287 -6732 18321 -6698
rect 18355 -6732 18389 -6698
rect 18423 -6732 18457 -6698
rect 18491 -6732 18525 -6698
rect 18559 -6732 18593 -6698
rect 18627 -6732 18661 -6698
rect 18695 -6732 18729 -6698
rect 18763 -6732 18797 -6698
rect 18831 -6732 18865 -6698
rect 18899 -6732 18933 -6698
rect 18967 -6732 19001 -6698
rect 19035 -6732 19069 -6698
rect 19103 -6732 19137 -6698
rect 19171 -6732 19205 -6698
rect 19239 -6732 19273 -6698
rect 19307 -6732 19341 -6698
rect 19375 -6732 19409 -6698
rect 19443 -6732 19477 -6698
rect 19511 -6732 19545 -6698
rect 19579 -6732 19613 -6698
rect 19647 -6732 19681 -6698
rect 19715 -6732 19749 -6698
rect 19783 -6732 19817 -6698
rect 19851 -6732 19885 -6698
rect 19919 -6732 19953 -6698
rect 19987 -6732 20021 -6698
rect 20055 -6732 20089 -6698
rect 20123 -6732 20157 -6698
rect 20191 -6732 20225 -6698
rect 20259 -6732 20293 -6698
rect 20327 -6732 20361 -6698
rect 20395 -6732 20429 -6698
rect 20463 -6732 20497 -6698
rect 20531 -6732 20565 -6698
rect 20599 -6732 20633 -6698
rect 20667 -6732 20701 -6698
rect 20735 -6732 20769 -6698
rect 20803 -6732 20837 -6698
rect 20871 -6732 20905 -6698
rect 16119 -6800 16153 -6766
rect 16119 -6868 16153 -6834
rect 16119 -6936 16153 -6902
rect 16119 -7004 16153 -6970
rect 16119 -7072 16153 -7038
rect 16119 -7140 16153 -7106
rect 16119 -7208 16153 -7174
rect 16119 -7276 16153 -7242
rect 16119 -7344 16153 -7310
rect 16119 -7412 16153 -7378
rect 16119 -7480 16153 -7446
rect 16119 -7548 16153 -7514
rect 16119 -7616 16153 -7582
rect 16119 -7684 16153 -7650
rect 16119 -7752 16153 -7718
rect 16119 -7820 16153 -7786
rect 16119 -7888 16153 -7854
rect 16119 -7956 16153 -7922
rect 16119 -8024 16153 -7990
rect 16119 -8092 16153 -8058
rect 20939 -6860 20973 -6826
rect 20939 -6928 20973 -6894
rect 20939 -6996 20973 -6962
rect 20939 -7064 20973 -7030
rect 20939 -7132 20973 -7098
rect 20939 -7200 20973 -7166
rect 20939 -7268 20973 -7234
rect 20939 -7336 20973 -7302
rect 20939 -7404 20973 -7370
rect 20939 -7472 20973 -7438
rect 20939 -7540 20973 -7506
rect 20939 -7608 20973 -7574
rect 20939 -7676 20973 -7642
rect 20939 -7744 20973 -7710
rect 20939 -7812 20973 -7778
rect 20939 -7880 20973 -7846
rect 20939 -7948 20973 -7914
rect 20939 -8016 20973 -7982
rect 20939 -8084 20973 -8050
rect 16119 -8160 16153 -8126
rect 16119 -8228 16153 -8194
rect 16119 -8296 16153 -8262
rect 16119 -8364 16153 -8330
rect 16119 -8432 16153 -8398
rect 16119 -8500 16153 -8466
rect 16119 -8568 16153 -8534
rect 16119 -8636 16153 -8602
rect 16119 -8704 16153 -8670
rect 16119 -8772 16153 -8738
rect 16119 -8840 16153 -8806
rect 16119 -8908 16153 -8874
rect 16119 -8976 16153 -8942
rect 16119 -9044 16153 -9010
rect 16119 -9112 16153 -9078
rect 20939 -8152 20973 -8118
rect 20939 -8220 20973 -8186
rect 20939 -8288 20973 -8254
rect 16119 -9180 16153 -9146
rect 16119 -9248 16153 -9214
rect 16119 -9316 16153 -9282
rect 16119 -9384 16153 -9350
rect 16119 -9452 16153 -9418
rect 16119 -9520 16153 -9486
rect 20747 -8356 20781 -8322
rect 20815 -8356 20849 -8322
rect 20679 -8451 20713 -8417
rect 20679 -8519 20713 -8485
rect 20679 -8587 20713 -8553
rect 20679 -8655 20713 -8621
rect 20679 -8723 20713 -8689
rect 20679 -8791 20713 -8757
rect 20679 -8859 20713 -8825
rect 20679 -8927 20713 -8893
rect 20679 -8995 20713 -8961
rect 20679 -9063 20713 -9029
rect 20679 -9131 20713 -9097
rect 20679 -9199 20713 -9165
rect 20679 -9267 20713 -9233
rect 20679 -9335 20713 -9301
rect 20679 -9403 20713 -9369
rect 20679 -9471 20713 -9437
rect 20679 -9539 20713 -9505
rect 16119 -9588 16153 -9554
rect 16119 -9656 16153 -9622
rect 16119 -9724 16153 -9690
rect 16119 -9792 16153 -9758
rect 16119 -9936 16153 -9902
rect 20679 -9607 20713 -9573
rect 20679 -9675 20713 -9641
rect 20679 -9743 20713 -9709
rect 20679 -9811 20713 -9777
rect 20679 -9879 20713 -9845
rect 16119 -10004 16153 -9970
rect 16119 -10072 16153 -10038
rect 16119 -10140 16153 -10106
rect 18349 -9996 18383 -9962
rect 18349 -10131 18383 -10097
rect 16119 -10208 16153 -10174
rect 20679 -9947 20713 -9913
rect 20679 -10015 20713 -9981
rect 20679 -10083 20713 -10049
rect 20679 -10151 20713 -10117
rect 16119 -10276 16153 -10242
rect 20679 -10219 20713 -10185
rect 20679 -10287 20713 -10253
rect 16119 -10344 16153 -10310
rect 16119 -10412 16153 -10378
rect 16119 -10480 16153 -10446
rect 20679 -10355 20713 -10321
rect 16119 -10548 16153 -10514
rect 20679 -10423 20713 -10389
rect 20679 -10491 20713 -10457
rect 22443 -10478 22477 -10444
rect 22588 -10478 22622 -10444
rect 22733 -10478 22767 -10444
rect 22878 -10478 22912 -10444
rect 23023 -10478 23057 -10444
rect 23168 -10478 23202 -10444
rect 23313 -10478 23347 -10444
rect 23458 -10478 23492 -10444
rect 23603 -10478 23637 -10444
rect 16119 -10616 16153 -10582
rect 20679 -10559 20713 -10525
rect 20679 -10627 20713 -10593
rect 16119 -10684 16153 -10650
rect 16119 -10752 16153 -10718
rect 16119 -10820 16153 -10786
rect 16119 -10888 16153 -10854
rect 16119 -10956 16153 -10922
rect 16119 -11024 16153 -10990
rect 16119 -11092 16153 -11058
rect 16119 -11160 16153 -11126
rect 16119 -11228 16153 -11194
rect 16119 -11296 16153 -11262
rect 20679 -10695 20713 -10661
rect 20679 -10763 20713 -10729
rect 20679 -10831 20713 -10797
rect 20679 -10899 20713 -10865
rect 20679 -10967 20713 -10933
rect 20679 -11035 20713 -11001
rect 20679 -11103 20713 -11069
rect 20679 -11171 20713 -11137
rect 20679 -11239 20713 -11205
rect 20679 -11307 20713 -11273
rect 16187 -11375 16221 -11341
rect 16255 -11375 16289 -11341
rect 16323 -11375 16357 -11341
rect 16391 -11375 16425 -11341
rect 16459 -11375 16493 -11341
rect 16527 -11375 16561 -11341
rect 16595 -11375 16629 -11341
rect 16663 -11375 16697 -11341
rect 16731 -11375 16765 -11341
rect 16799 -11375 16833 -11341
rect 16867 -11375 16901 -11341
rect 16935 -11375 16969 -11341
rect 17003 -11375 17037 -11341
rect 17071 -11375 17105 -11341
rect 17139 -11375 17173 -11341
rect 17207 -11375 17241 -11341
rect 17275 -11375 17309 -11341
rect 17343 -11375 17377 -11341
rect 17411 -11375 17445 -11341
rect 17479 -11375 17513 -11341
rect 17547 -11375 17581 -11341
rect 17615 -11375 17649 -11341
rect 17683 -11375 17717 -11341
rect 17751 -11375 17785 -11341
rect 17819 -11375 17853 -11341
rect 17887 -11375 17921 -11341
rect 17955 -11375 17989 -11341
rect 18023 -11375 18057 -11341
rect 18091 -11375 18125 -11341
rect 18159 -11375 18193 -11341
rect 18227 -11375 18261 -11341
rect 18295 -11375 18329 -11341
rect 18363 -11375 18397 -11341
rect 18431 -11375 18465 -11341
rect 18499 -11375 18533 -11341
rect 18567 -11375 18601 -11341
rect 18635 -11375 18669 -11341
rect 18703 -11375 18737 -11341
rect 18771 -11375 18805 -11341
rect 18839 -11375 18873 -11341
rect 18907 -11375 18941 -11341
rect 18975 -11375 19009 -11341
rect 19043 -11375 19077 -11341
rect 19111 -11375 19145 -11341
rect 19179 -11375 19213 -11341
rect 19247 -11375 19281 -11341
rect 19315 -11375 19349 -11341
rect 19383 -11375 19417 -11341
rect 19451 -11375 19485 -11341
rect 19519 -11375 19553 -11341
rect 19587 -11375 19621 -11341
rect 19655 -11375 19689 -11341
rect 19723 -11375 19757 -11341
rect 19791 -11375 19825 -11341
rect 19859 -11375 19893 -11341
rect 19927 -11375 19961 -11341
rect 19995 -11375 20029 -11341
rect 20063 -11375 20097 -11341
rect 20131 -11375 20165 -11341
rect 20199 -11375 20233 -11341
rect 20267 -11375 20301 -11341
rect 20335 -11375 20369 -11341
rect 20403 -11375 20437 -11341
rect 20471 -11375 20505 -11341
rect 20539 -11375 20573 -11341
rect 20607 -11375 20641 -11341
rect 22576 -12023 22610 -11989
rect 22644 -12023 22678 -11989
rect 22712 -12023 22746 -11989
rect 22780 -12023 22814 -11989
rect 22848 -12023 22882 -11989
rect 22916 -12023 22950 -11989
rect 22984 -12023 23018 -11989
rect 23052 -12023 23086 -11989
rect 23120 -12023 23154 -11989
rect 23188 -12023 23222 -11989
rect 23256 -12023 23290 -11989
rect 23324 -12023 23358 -11989
rect 23392 -12023 23426 -11989
rect 23460 -12023 23494 -11989
rect 23528 -12023 23562 -11989
rect 23596 -12023 23630 -11989
rect 23664 -12023 23698 -11989
rect 23732 -12023 23766 -11989
rect 23800 -12023 23834 -11989
rect 23868 -12023 23902 -11989
rect 23936 -12023 23970 -11989
rect 24004 -12023 24038 -11989
rect 24072 -12023 24106 -11989
rect 24140 -12023 24174 -11989
rect 24208 -12023 24242 -11989
rect 24276 -12023 24310 -11989
rect 24344 -12023 24378 -11989
rect 24412 -12023 24446 -11989
rect 24480 -12023 24514 -11989
<< poly >>
rect 18814 -9227 19070 -9211
rect 18814 -9261 18830 -9227
rect 18864 -9261 18925 -9227
rect 18959 -9261 19020 -9227
rect 19054 -9261 19070 -9227
rect 18814 -9277 19070 -9261
rect 18814 -9309 18914 -9277
rect 18970 -9309 19070 -9277
rect 19520 -9227 20043 -9211
rect 19520 -9261 19536 -9227
rect 19570 -9261 19612 -9227
rect 19646 -9261 19688 -9227
rect 19722 -9261 19764 -9227
rect 19798 -9261 19840 -9227
rect 19874 -9261 19916 -9227
rect 19950 -9261 19993 -9227
rect 20027 -9261 20043 -9227
rect 19520 -9277 20043 -9261
rect 19520 -9309 19620 -9277
rect 19676 -9309 19776 -9277
rect 19943 -9309 20043 -9277
rect 18814 -9541 18914 -9509
rect 18970 -9541 19070 -9509
rect 19520 -9541 19620 -9509
rect 19676 -9541 19776 -9509
rect 19943 -9541 20043 -9509
rect 17015 -10243 17192 -10206
rect 17015 -10277 17031 -10243
rect 17065 -10277 17099 -10243
rect 17133 -10277 17192 -10243
rect 17015 -10306 17192 -10277
rect 17492 -10306 17524 -10206
rect 17160 -10462 17192 -10362
rect 17492 -10378 17590 -10362
rect 17492 -10412 17540 -10378
rect 17574 -10412 17590 -10378
rect 17857 -10380 18257 -10348
rect 18313 -10380 18713 -10348
rect 17492 -10446 17590 -10412
rect 17492 -10462 17540 -10446
rect 17524 -10480 17540 -10462
rect 17574 -10480 17590 -10446
rect 17524 -10496 17590 -10480
rect 17857 -10562 18257 -10530
rect 18313 -10562 18713 -10530
rect 17857 -10578 18713 -10562
rect 17857 -10612 17873 -10578
rect 17907 -10612 17945 -10578
rect 17979 -10612 18017 -10578
rect 18051 -10612 18089 -10578
rect 18123 -10612 18161 -10578
rect 18195 -10612 18233 -10578
rect 18267 -10612 18305 -10578
rect 18339 -10612 18377 -10578
rect 18411 -10612 18449 -10578
rect 18483 -10612 18521 -10578
rect 18555 -10612 18592 -10578
rect 18626 -10612 18663 -10578
rect 18697 -10612 18713 -10578
rect 17857 -10628 18713 -10612
<< polycont >>
rect 18830 -9261 18864 -9227
rect 18925 -9261 18959 -9227
rect 19020 -9261 19054 -9227
rect 19536 -9261 19570 -9227
rect 19612 -9261 19646 -9227
rect 19688 -9261 19722 -9227
rect 19764 -9261 19798 -9227
rect 19840 -9261 19874 -9227
rect 19916 -9261 19950 -9227
rect 19993 -9261 20027 -9227
rect 17031 -10277 17065 -10243
rect 17099 -10277 17133 -10243
rect 17540 -10412 17574 -10378
rect 17540 -10480 17574 -10446
rect 17873 -10612 17907 -10578
rect 17945 -10612 17979 -10578
rect 18017 -10612 18051 -10578
rect 18089 -10612 18123 -10578
rect 18161 -10612 18195 -10578
rect 18233 -10612 18267 -10578
rect 18305 -10612 18339 -10578
rect 18377 -10612 18411 -10578
rect 18449 -10612 18483 -10578
rect 18521 -10612 18555 -10578
rect 18592 -10612 18626 -10578
rect 18663 -10612 18697 -10578
<< locali >>
rect 16119 -6732 16191 -6698
rect 16225 -6732 16247 -6698
rect 16305 -6732 16315 -6698
rect 16349 -6732 16383 -6698
rect 16417 -6732 16451 -6698
rect 16485 -6732 16519 -6698
rect 16553 -6732 16587 -6698
rect 16621 -6732 16655 -6698
rect 16689 -6732 16723 -6698
rect 16757 -6732 16791 -6698
rect 16825 -6732 16859 -6698
rect 16893 -6732 16927 -6698
rect 16961 -6732 16995 -6698
rect 17029 -6732 17063 -6698
rect 17097 -6732 17131 -6698
rect 17165 -6732 17199 -6698
rect 17233 -6732 17267 -6698
rect 17301 -6732 17335 -6698
rect 17369 -6732 17403 -6698
rect 17437 -6732 17471 -6698
rect 17505 -6732 17539 -6698
rect 17573 -6732 17607 -6698
rect 17641 -6732 17675 -6698
rect 17709 -6732 17743 -6698
rect 17777 -6732 17811 -6698
rect 17845 -6732 17879 -6698
rect 17913 -6732 17947 -6698
rect 17981 -6732 18015 -6698
rect 18049 -6732 18083 -6698
rect 18117 -6732 18151 -6698
rect 18185 -6732 18219 -6698
rect 18253 -6732 18287 -6698
rect 18321 -6732 18355 -6698
rect 18389 -6732 18423 -6698
rect 18457 -6732 18491 -6698
rect 18525 -6732 18559 -6698
rect 18593 -6732 18627 -6698
rect 18661 -6732 18695 -6698
rect 18729 -6732 18763 -6698
rect 18797 -6732 18831 -6698
rect 18865 -6732 18899 -6698
rect 18933 -6732 18967 -6698
rect 19001 -6732 19035 -6698
rect 19069 -6732 19103 -6698
rect 19137 -6732 19171 -6698
rect 19205 -6732 19239 -6698
rect 19273 -6732 19307 -6698
rect 19341 -6732 19375 -6698
rect 19409 -6732 19443 -6698
rect 19477 -6732 19511 -6698
rect 19545 -6732 19579 -6698
rect 19613 -6732 19647 -6698
rect 19681 -6732 19715 -6698
rect 19749 -6732 19783 -6698
rect 19817 -6732 19851 -6698
rect 19885 -6732 19919 -6698
rect 19953 -6732 19987 -6698
rect 20021 -6732 20055 -6698
rect 20089 -6732 20123 -6698
rect 20157 -6732 20191 -6698
rect 20225 -6732 20259 -6698
rect 20293 -6732 20327 -6698
rect 20361 -6732 20395 -6698
rect 20429 -6732 20463 -6698
rect 20497 -6732 20531 -6698
rect 20565 -6732 20599 -6698
rect 20633 -6732 20667 -6698
rect 20701 -6732 20735 -6698
rect 20769 -6732 20803 -6698
rect 20837 -6732 20871 -6698
rect 20905 -6732 20973 -6698
rect 16119 -6766 16153 -6732
rect 16119 -6834 16153 -6804
rect 16119 -6902 16153 -6876
rect 16119 -6970 16153 -6948
rect 16119 -7038 16153 -7020
rect 16119 -7106 16153 -7092
rect 16119 -7174 16153 -7164
rect 20939 -6826 20973 -6732
rect 20939 -6894 20973 -6860
rect 20939 -6962 20973 -6928
rect 20939 -7030 20973 -6996
rect 20939 -7098 20973 -7064
rect 20939 -7166 20973 -7132
rect 20939 -7225 20973 -7200
rect 16119 -7242 16153 -7236
rect 16119 -7310 16153 -7308
rect 16119 -7346 16153 -7344
rect 16119 -7418 16153 -7412
rect 16119 -7490 16153 -7480
rect 16119 -7562 16153 -7548
rect 16119 -7634 16153 -7616
rect 16119 -7706 16153 -7684
rect 16119 -7778 16153 -7752
rect 16119 -7850 16153 -7820
rect 16119 -7922 16153 -7888
rect 16119 -7990 16153 -7956
rect 16119 -8058 16153 -8028
rect 16119 -8126 16153 -8100
rect 20954 -7234 20973 -7225
rect 20920 -7268 20939 -7259
rect 20920 -7299 20973 -7268
rect 20954 -7302 20973 -7299
rect 20920 -7336 20939 -7333
rect 20920 -7370 20973 -7336
rect 20920 -7373 20939 -7370
rect 20954 -7407 20973 -7404
rect 20920 -7438 20973 -7407
rect 20920 -7446 20939 -7438
rect 20954 -7480 20973 -7472
rect 20920 -7506 20973 -7480
rect 20920 -7519 20939 -7506
rect 20954 -7553 20973 -7540
rect 20920 -7574 20973 -7553
rect 20920 -7592 20939 -7574
rect 20954 -7626 20973 -7608
rect 20920 -7642 20973 -7626
rect 20920 -7665 20939 -7642
rect 20954 -7699 20973 -7676
rect 20920 -7710 20973 -7699
rect 20920 -7738 20939 -7710
rect 20954 -7772 20973 -7744
rect 20920 -7778 20973 -7772
rect 20920 -7811 20939 -7778
rect 20954 -7845 20973 -7812
rect 20920 -7846 20973 -7845
rect 20920 -7880 20939 -7846
rect 20920 -7884 20973 -7880
rect 20954 -7914 20973 -7884
rect 20920 -7948 20939 -7918
rect 20920 -7957 20973 -7948
rect 20954 -7982 20973 -7957
rect 20920 -8016 20939 -7991
rect 20920 -8030 20973 -8016
rect 20954 -8050 20973 -8030
rect 20920 -8084 20939 -8064
rect 20920 -8103 20973 -8084
rect 16119 -8194 16153 -8172
rect 16119 -8262 16153 -8244
rect 16119 -8330 16153 -8316
rect 16119 -8398 16153 -8388
rect 16119 -8466 16153 -8460
rect 16119 -8534 16153 -8532
rect 16119 -8570 16153 -8568
rect 16119 -8642 16153 -8636
rect 20174 -8139 20466 -8105
rect 20208 -8173 20260 -8139
rect 20294 -8173 20346 -8139
rect 20380 -8173 20432 -8139
rect 20174 -8210 20466 -8173
rect 20208 -8244 20260 -8210
rect 20294 -8244 20346 -8210
rect 20380 -8244 20432 -8210
rect 20174 -8281 20466 -8244
rect 20208 -8315 20260 -8281
rect 20294 -8315 20346 -8281
rect 20380 -8315 20432 -8281
rect 20174 -8352 20466 -8315
rect 20954 -8118 20973 -8103
rect 20920 -8152 20939 -8137
rect 20920 -8176 20973 -8152
rect 20954 -8186 20973 -8176
rect 20920 -8220 20939 -8210
rect 20920 -8249 20973 -8220
rect 20954 -8254 20973 -8249
rect 20920 -8288 20939 -8283
rect 20920 -8322 20973 -8288
rect 20208 -8386 20260 -8352
rect 20294 -8386 20346 -8352
rect 20380 -8386 20432 -8352
rect 20174 -8423 20466 -8386
rect 20208 -8457 20260 -8423
rect 20294 -8457 20346 -8423
rect 20380 -8457 20432 -8423
rect 20174 -8494 20466 -8457
rect 20208 -8528 20260 -8494
rect 20294 -8528 20346 -8494
rect 20380 -8528 20432 -8494
rect 20174 -8565 20466 -8528
rect 20208 -8599 20260 -8565
rect 20294 -8599 20346 -8565
rect 20380 -8599 20432 -8565
rect 20174 -8636 20466 -8599
rect 20208 -8670 20260 -8636
rect 20294 -8670 20346 -8636
rect 20380 -8670 20432 -8636
rect 16119 -8714 16153 -8704
rect 17398 -8680 18957 -8675
rect 17398 -8714 17873 -8680
rect 17907 -8714 17949 -8680
rect 17983 -8714 18025 -8680
rect 18059 -8714 18101 -8680
rect 18135 -8714 18177 -8680
rect 18211 -8714 18254 -8680
rect 18288 -8714 18331 -8680
rect 18365 -8714 18408 -8680
rect 18442 -8714 18485 -8680
rect 18519 -8714 18957 -8680
rect 17398 -8727 18957 -8714
rect 20174 -8707 20466 -8670
rect 16119 -8787 16153 -8772
rect 16119 -8860 16153 -8840
rect 16119 -8933 16153 -8908
rect 16119 -9006 16153 -8976
rect 16119 -9078 16153 -9044
rect 16119 -9146 16153 -9113
rect 20208 -8741 20260 -8707
rect 20294 -8741 20346 -8707
rect 20380 -8741 20432 -8707
rect 20174 -8779 20466 -8741
rect 20208 -8813 20260 -8779
rect 20294 -8813 20346 -8779
rect 20380 -8813 20432 -8779
rect 20174 -8851 20466 -8813
rect 20208 -8885 20260 -8851
rect 20294 -8885 20346 -8851
rect 20380 -8885 20432 -8851
rect 20174 -8923 20466 -8885
rect 20208 -8957 20260 -8923
rect 20294 -8957 20346 -8923
rect 20380 -8957 20432 -8923
rect 20174 -8995 20466 -8957
rect 20208 -9029 20260 -8995
rect 20294 -9029 20346 -8995
rect 20380 -9029 20432 -8995
rect 20174 -9067 20466 -9029
rect 20208 -9101 20260 -9067
rect 20294 -9101 20346 -9067
rect 20380 -9101 20432 -9067
rect 18348 -9167 18372 -9133
rect 18406 -9167 18441 -9133
rect 18475 -9167 18510 -9133
rect 18544 -9167 18579 -9133
rect 18613 -9167 18648 -9133
rect 18682 -9167 18717 -9133
rect 18751 -9167 18786 -9133
rect 18820 -9167 18855 -9133
rect 18889 -9167 18924 -9133
rect 18958 -9167 18993 -9133
rect 19027 -9167 19062 -9133
rect 19096 -9167 19131 -9133
rect 19165 -9167 19200 -9133
rect 19234 -9167 19269 -9133
rect 19303 -9167 19338 -9133
rect 19372 -9167 19396 -9133
rect 20174 -9139 20466 -9101
rect 16119 -9214 16153 -9186
rect 20208 -9173 20260 -9139
rect 20294 -9173 20346 -9139
rect 20380 -9173 20432 -9139
rect 20174 -9211 20466 -9173
rect 18791 -9259 18829 -9225
rect 16119 -9282 16153 -9259
rect 18814 -9261 18830 -9259
rect 18864 -9261 18925 -9227
rect 18959 -9261 19020 -9227
rect 19054 -9261 19070 -9227
rect 19520 -9261 19536 -9227
rect 19570 -9261 19612 -9227
rect 19646 -9261 19688 -9227
rect 19722 -9261 19747 -9227
rect 19798 -9261 19819 -9227
rect 19874 -9261 19916 -9227
rect 19950 -9261 19993 -9227
rect 20027 -9261 20043 -9227
rect 20208 -9245 20260 -9211
rect 20294 -9245 20346 -9211
rect 20380 -9245 20432 -9211
rect 20174 -9283 20466 -9245
rect 16119 -9350 16153 -9332
rect 16119 -9418 16153 -9405
rect 16119 -9486 16153 -9478
rect 16119 -9554 16153 -9551
rect 16119 -9590 16153 -9588
rect 18764 -9305 18808 -9303
rect 18764 -9355 18769 -9305
rect 18803 -9355 18808 -9305
rect 18764 -9377 18808 -9355
rect 18764 -9423 18769 -9377
rect 18803 -9423 18808 -9377
rect 18764 -9449 18808 -9423
rect 18764 -9491 18769 -9449
rect 18803 -9491 18808 -9449
rect 18764 -9620 18808 -9491
rect 18925 -9377 18959 -9355
rect 18925 -9449 18959 -9423
rect 18925 -9507 18959 -9491
rect 19115 -9355 19150 -9310
rect 19081 -9377 19150 -9355
rect 19115 -9423 19150 -9377
rect 19081 -9449 19150 -9423
rect 19115 -9491 19150 -9449
rect 19081 -9507 19150 -9491
rect 19106 -9620 19150 -9507
rect 19458 -9327 19509 -9311
rect 19458 -9369 19475 -9327
rect 19458 -9395 19509 -9369
rect 19458 -9441 19475 -9395
rect 19458 -9463 19509 -9441
rect 19458 -9513 19475 -9463
rect 19631 -9327 19665 -9311
rect 19631 -9395 19665 -9369
rect 19631 -9463 19665 -9441
rect 19787 -9327 19864 -9311
rect 19821 -9369 19864 -9327
rect 19787 -9395 19864 -9369
rect 19821 -9441 19864 -9395
rect 19787 -9463 19864 -9441
rect 19821 -9513 19864 -9463
rect 19898 -9327 19910 -9311
rect 19932 -9361 19944 -9343
rect 19898 -9381 19944 -9361
rect 19898 -9395 19910 -9381
rect 20054 -9324 20088 -9311
rect 20208 -9317 20260 -9283
rect 20294 -9317 20346 -9283
rect 20380 -9317 20432 -9283
rect 20174 -9351 20466 -9317
rect 20679 -8356 20747 -8322
rect 20797 -8356 20815 -8322
rect 20882 -8356 20973 -8322
rect 20679 -8394 20713 -8356
rect 20679 -8468 20713 -8451
rect 20679 -8542 20713 -8519
rect 20679 -8616 20713 -8587
rect 20679 -8689 20713 -8655
rect 20679 -8757 20713 -8724
rect 20679 -8825 20713 -8798
rect 20679 -8893 20713 -8872
rect 20679 -8961 20713 -8946
rect 20679 -9029 20713 -9020
rect 20679 -9097 20713 -9094
rect 20679 -9134 20713 -9131
rect 20679 -9208 20713 -9199
rect 20679 -9282 20713 -9267
rect 20054 -9395 20088 -9361
rect 19898 -9463 19932 -9429
rect 19898 -9513 19932 -9497
rect 20054 -9463 20088 -9430
rect 20054 -9513 20088 -9497
rect 20679 -9356 20713 -9335
rect 20679 -9430 20713 -9403
rect 20679 -9504 20713 -9471
rect 19458 -9620 19502 -9513
rect 16119 -9663 16153 -9656
rect 16119 -9736 16153 -9724
rect 16119 -9809 16153 -9792
rect 16119 -9882 16153 -9843
rect 16119 -9955 16153 -9936
rect 16119 -10028 16153 -10004
rect 16119 -10101 16153 -10072
rect 16119 -10174 16153 -10140
rect 18349 -9962 18383 -9938
rect 18349 -10040 18383 -9996
rect 18349 -10097 18383 -10074
rect 18349 -10155 18383 -10146
rect 17226 -10195 17242 -10161
rect 17276 -10195 17310 -10161
rect 17344 -10195 17378 -10161
rect 17412 -10195 17446 -10161
rect 17480 -10195 17496 -10161
rect 19805 -10163 19864 -9513
rect 20250 -9622 20284 -9584
rect 20679 -9573 20713 -9539
rect 20412 -9665 20446 -9627
rect 20679 -9641 20713 -9612
rect 20330 -9749 20364 -9711
rect 20679 -9709 20713 -9686
rect 20679 -9777 20713 -9760
rect 20679 -9845 20713 -9834
rect 20679 -9913 20713 -9908
rect 20679 -9948 20713 -9947
rect 20679 -10022 20713 -10015
rect 20250 -10112 20284 -10074
rect 20679 -10096 20713 -10083
rect 16119 -10242 16153 -10208
rect 17256 -10229 17294 -10195
rect 17328 -10229 17496 -10195
rect 16634 -10271 16668 -10233
rect 17226 -10235 17496 -10229
rect 20679 -10170 20713 -10151
rect 16119 -10310 16153 -10281
rect 16119 -10378 16153 -10354
rect 17065 -10277 17071 -10243
rect 17133 -10277 17149 -10243
rect 20679 -10244 20713 -10219
rect 16553 -10351 16587 -10313
rect 16715 -10351 16749 -10313
rect 17274 -10317 17327 -10315
rect 17361 -10317 17414 -10315
rect 16985 -10370 17101 -10346
rect 17226 -10349 17240 -10317
rect 17226 -10351 17242 -10349
rect 17276 -10351 17310 -10317
rect 17361 -10349 17378 -10317
rect 17344 -10351 17378 -10349
rect 17412 -10349 17414 -10317
rect 17412 -10351 17446 -10349
rect 17480 -10351 17496 -10317
rect 18280 -10349 18318 -10315
rect 20679 -10318 20713 -10287
rect 17019 -10371 17067 -10370
rect 16119 -10446 16153 -10427
rect 17019 -10404 17063 -10371
rect 17013 -10405 17063 -10404
rect 17097 -10405 17101 -10404
rect 16979 -10438 17101 -10405
rect 16979 -10443 16985 -10438
rect 17019 -10443 17067 -10438
rect 16119 -10514 16153 -10500
rect 17019 -10472 17063 -10443
rect 17540 -10378 17574 -10362
rect 17540 -10429 17541 -10412
rect 17540 -10446 17575 -10429
rect 17574 -10467 17575 -10446
rect 17013 -10477 17063 -10472
rect 17097 -10477 17101 -10472
rect 16478 -10521 16512 -10483
rect 16985 -10496 17101 -10477
rect 17256 -10473 17294 -10468
rect 17276 -10502 17294 -10473
rect 17226 -10507 17242 -10502
rect 17276 -10507 17310 -10502
rect 17344 -10507 17378 -10473
rect 17412 -10507 17446 -10473
rect 17480 -10507 17496 -10473
rect 17540 -10496 17541 -10480
rect 17812 -10416 17846 -10400
rect 17812 -10484 17846 -10458
rect 17812 -10534 17846 -10530
rect 18268 -10416 18302 -10349
rect 20679 -10389 20713 -10355
rect 18268 -10484 18302 -10450
rect 18268 -10534 18302 -10518
rect 18724 -10416 18758 -10400
rect 18724 -10458 18736 -10450
rect 18724 -10484 18770 -10458
rect 18758 -10496 18770 -10484
rect 18724 -10530 18736 -10518
rect 20679 -10457 20713 -10426
rect 22409 -10478 22415 -10444
rect 22477 -10478 22492 -10444
rect 22526 -10478 22569 -10444
rect 22622 -10478 22646 -10444
rect 22680 -10478 22723 -10444
rect 22767 -10478 22800 -10444
rect 22834 -10478 22877 -10444
rect 22912 -10478 22954 -10444
rect 22988 -10478 23023 -10444
rect 23065 -10478 23108 -10444
rect 23142 -10478 23168 -10444
rect 23219 -10478 23261 -10444
rect 23295 -10478 23313 -10444
rect 23371 -10478 23413 -10444
rect 23447 -10478 23458 -10444
rect 23523 -10478 23565 -10444
rect 23599 -10478 23603 -10444
rect 23637 -10478 23671 -10444
rect 20679 -10525 20713 -10499
rect 18724 -10534 18758 -10530
rect 16119 -10582 16153 -10573
rect 16119 -10650 16153 -10646
rect 16635 -10647 16669 -10609
rect 17857 -10612 17873 -10578
rect 17907 -10612 17919 -10578
rect 17979 -10612 17998 -10578
rect 18051 -10612 18077 -10578
rect 18123 -10612 18156 -10578
rect 18195 -10612 18233 -10578
rect 18269 -10612 18305 -10578
rect 18348 -10612 18377 -10578
rect 18427 -10612 18449 -10578
rect 18505 -10612 18521 -10578
rect 18583 -10612 18592 -10578
rect 18626 -10612 18627 -10578
rect 18661 -10612 18663 -10578
rect 18697 -10612 18705 -10578
rect 20679 -10593 20713 -10572
rect 20679 -10661 20713 -10645
rect 16119 -10685 16153 -10684
rect 16119 -10758 16153 -10752
rect 16800 -10747 16834 -10709
rect 20679 -10729 20713 -10718
rect 16119 -10831 16153 -10820
rect 16119 -10904 16153 -10888
rect 16119 -10977 16153 -10956
rect 16119 -11050 16153 -11024
rect 16119 -11123 16153 -11092
rect 16119 -11194 16153 -11160
rect 16119 -11262 16153 -11230
rect 16119 -11341 16153 -11303
rect 20679 -10797 20713 -10791
rect 20679 -10865 20713 -10864
rect 22724 -10845 22758 -10807
rect 22905 -10845 22939 -10807
rect 23054 -10864 23072 -10830
rect 23106 -10864 23119 -10830
rect 20679 -10903 20713 -10899
rect 20679 -10976 20713 -10967
rect 20679 -11049 20713 -11035
rect 23054 -10902 23119 -10864
rect 23054 -10936 23072 -10902
rect 23106 -10936 23119 -10902
rect 23208 -10922 23246 -10888
rect 20679 -11122 20713 -11103
rect 20679 -11195 20713 -11171
rect 22458 -11141 22492 -11103
rect 22548 -11141 22582 -11103
rect 22810 -11141 22844 -11103
rect 23054 -11064 23119 -10936
rect 23054 -11068 23069 -11064
rect 22904 -11134 22938 -11096
rect 23103 -11068 23119 -11064
rect 23069 -11136 23103 -11098
rect 23254 -11136 23288 -11098
rect 23426 -11141 23460 -11103
rect 23514 -11141 23548 -11103
rect 20679 -11268 20713 -11239
rect 20679 -11341 20713 -11307
rect 16119 -11375 16187 -11341
rect 16225 -11375 16255 -11341
rect 16297 -11375 16323 -11341
rect 16369 -11375 16391 -11341
rect 16441 -11375 16459 -11341
rect 16513 -11375 16527 -11341
rect 16585 -11375 16595 -11341
rect 16657 -11375 16663 -11341
rect 16729 -11375 16731 -11341
rect 16765 -11375 16767 -11341
rect 16833 -11375 16839 -11341
rect 16901 -11375 16911 -11341
rect 16969 -11375 16983 -11341
rect 17037 -11375 17055 -11341
rect 17105 -11375 17127 -11341
rect 17173 -11375 17199 -11341
rect 17241 -11375 17271 -11341
rect 17309 -11375 17343 -11341
rect 17377 -11375 17411 -11341
rect 17449 -11375 17479 -11341
rect 17521 -11375 17547 -11341
rect 17593 -11375 17615 -11341
rect 17665 -11375 17683 -11341
rect 17737 -11375 17751 -11341
rect 17809 -11375 17819 -11341
rect 17881 -11375 17887 -11341
rect 17953 -11375 17955 -11341
rect 17989 -11375 17991 -11341
rect 18057 -11375 18063 -11341
rect 18125 -11375 18135 -11341
rect 18193 -11375 18207 -11341
rect 18261 -11375 18279 -11341
rect 18329 -11375 18351 -11341
rect 18397 -11375 18423 -11341
rect 18465 -11375 18495 -11341
rect 18533 -11375 18567 -11341
rect 18601 -11375 18635 -11341
rect 18673 -11375 18703 -11341
rect 18745 -11375 18771 -11341
rect 18817 -11375 18839 -11341
rect 18889 -11375 18907 -11341
rect 18962 -11375 18975 -11341
rect 19035 -11375 19043 -11341
rect 19108 -11375 19111 -11341
rect 19145 -11375 19147 -11341
rect 19213 -11375 19220 -11341
rect 19281 -11375 19293 -11341
rect 19349 -11375 19366 -11341
rect 19417 -11375 19439 -11341
rect 19485 -11375 19512 -11341
rect 19553 -11375 19585 -11341
rect 19621 -11375 19655 -11341
rect 19692 -11375 19723 -11341
rect 19765 -11375 19791 -11341
rect 19838 -11375 19859 -11341
rect 19911 -11375 19927 -11341
rect 19984 -11375 19995 -11341
rect 20057 -11375 20063 -11341
rect 20130 -11375 20131 -11341
rect 20165 -11375 20169 -11341
rect 20233 -11375 20242 -11341
rect 20301 -11375 20315 -11341
rect 20369 -11375 20388 -11341
rect 20437 -11375 20461 -11341
rect 20505 -11375 20534 -11341
rect 20573 -11375 20607 -11341
rect 20641 -11375 20713 -11341
rect 22435 -11466 22459 -11432
rect 22493 -11466 22494 -11432
rect 22528 -11466 22529 -11432
rect 22563 -11466 22567 -11432
rect 22632 -11466 22640 -11432
rect 22701 -11466 22713 -11432
rect 22770 -11466 22786 -11432
rect 22839 -11466 22859 -11432
rect 22908 -11466 22932 -11432
rect 22977 -11466 23005 -11432
rect 23046 -11466 23078 -11432
rect 23115 -11466 23150 -11432
rect 23185 -11466 23219 -11432
rect 23258 -11466 23288 -11432
rect 23331 -11466 23357 -11432
rect 23403 -11466 23426 -11432
rect 23475 -11466 23495 -11432
rect 23547 -11466 23564 -11432
rect 23619 -11466 23633 -11432
rect 23691 -11466 23702 -11432
rect 23763 -11466 23771 -11432
rect 23835 -11466 23840 -11432
rect 23907 -11466 23909 -11432
rect 23943 -11466 23945 -11432
rect 24012 -11466 24017 -11432
rect 24081 -11466 24089 -11432
rect 24150 -11466 24161 -11432
rect 24219 -11466 24233 -11432
rect 24288 -11466 24305 -11432
rect 24357 -11466 24377 -11432
rect 24426 -11466 24449 -11432
rect 24495 -11466 24521 -11432
rect 24564 -11466 24593 -11432
rect 24633 -11466 24665 -11432
rect 24702 -11466 24737 -11432
rect 24771 -11466 24806 -11432
rect 24843 -11466 24875 -11432
rect 24915 -11466 24944 -11432
rect 24987 -11466 25013 -11432
rect 25059 -11466 25082 -11432
rect 25131 -11466 25151 -11432
rect 25203 -11466 25220 -11432
rect 25275 -11466 25289 -11432
rect 25347 -11466 25358 -11432
rect 25419 -11466 25427 -11432
rect 25491 -11466 25496 -11432
rect 25563 -11466 25565 -11432
rect 25599 -11466 25601 -11432
rect 25668 -11466 25673 -11432
rect 25737 -11466 25745 -11432
rect 25806 -11466 25817 -11432
rect 25875 -11466 25889 -11432
rect 25944 -11466 25961 -11432
rect 26013 -11466 26033 -11432
rect 26082 -11466 26105 -11432
rect 26151 -11466 26177 -11432
rect 26220 -11466 26249 -11432
rect 22552 -12023 22576 -11989
rect 22610 -12023 22644 -11989
rect 22678 -12023 22712 -11989
rect 22746 -12023 22780 -11989
rect 22814 -12023 22848 -11989
rect 22882 -12023 22916 -11989
rect 22950 -12023 22984 -11989
rect 23018 -12023 23052 -11989
rect 23086 -12023 23120 -11989
rect 23154 -12023 23188 -11989
rect 23222 -12023 23256 -11989
rect 23290 -12023 23324 -11989
rect 23358 -12023 23392 -11989
rect 23426 -12023 23460 -11989
rect 23494 -12023 23528 -11989
rect 23562 -12023 23596 -11989
rect 23630 -12023 23664 -11989
rect 23698 -12023 23732 -11989
rect 23766 -12023 23800 -11989
rect 23834 -12023 23868 -11989
rect 23902 -12023 23936 -11989
rect 23970 -12023 24004 -11989
rect 24038 -12023 24072 -11989
rect 24106 -12023 24140 -11989
rect 24174 -12023 24208 -11989
rect 24242 -12023 24276 -11989
rect 24310 -12023 24344 -11989
rect 24378 -12023 24412 -11989
rect 24446 -12023 24480 -11989
rect 24514 -12023 24538 -11989
rect 22560 -12088 22594 -12023
rect 22912 -12088 22946 -12023
rect 23264 -12088 23298 -12023
rect 23616 -12088 23650 -12023
rect 23968 -12088 24002 -12023
rect 24320 -12088 24354 -12023
rect 17860 -13575 18062 -13541
<< viali >>
rect 16191 -6732 16225 -6698
rect 16271 -6732 16281 -6698
rect 16281 -6732 16305 -6698
rect 16119 -6800 16153 -6770
rect 16119 -6804 16153 -6800
rect 16119 -6868 16153 -6842
rect 16119 -6876 16153 -6868
rect 16119 -6936 16153 -6914
rect 16119 -6948 16153 -6936
rect 16119 -7004 16153 -6986
rect 16119 -7020 16153 -7004
rect 16119 -7072 16153 -7058
rect 16119 -7092 16153 -7072
rect 16119 -7140 16153 -7130
rect 16119 -7164 16153 -7140
rect 16119 -7208 16153 -7202
rect 16119 -7236 16153 -7208
rect 16119 -7276 16153 -7274
rect 16119 -7308 16153 -7276
rect 16119 -7378 16153 -7346
rect 16119 -7380 16153 -7378
rect 16119 -7446 16153 -7418
rect 16119 -7452 16153 -7446
rect 16119 -7514 16153 -7490
rect 16119 -7524 16153 -7514
rect 16119 -7582 16153 -7562
rect 16119 -7596 16153 -7582
rect 16119 -7650 16153 -7634
rect 16119 -7668 16153 -7650
rect 16119 -7718 16153 -7706
rect 16119 -7740 16153 -7718
rect 16119 -7786 16153 -7778
rect 16119 -7812 16153 -7786
rect 16119 -7854 16153 -7850
rect 16119 -7884 16153 -7854
rect 16119 -7956 16153 -7922
rect 16119 -8024 16153 -7994
rect 16119 -8028 16153 -8024
rect 16119 -8092 16153 -8066
rect 16119 -8100 16153 -8092
rect 20920 -7234 20954 -7225
rect 20920 -7259 20939 -7234
rect 20939 -7259 20954 -7234
rect 20920 -7302 20954 -7299
rect 20920 -7333 20939 -7302
rect 20939 -7333 20954 -7302
rect 20920 -7404 20939 -7373
rect 20939 -7404 20954 -7373
rect 20920 -7407 20954 -7404
rect 20920 -7472 20939 -7446
rect 20939 -7472 20954 -7446
rect 20920 -7480 20954 -7472
rect 20920 -7540 20939 -7519
rect 20939 -7540 20954 -7519
rect 20920 -7553 20954 -7540
rect 20920 -7608 20939 -7592
rect 20939 -7608 20954 -7592
rect 20920 -7626 20954 -7608
rect 20920 -7676 20939 -7665
rect 20939 -7676 20954 -7665
rect 20920 -7699 20954 -7676
rect 20920 -7744 20939 -7738
rect 20939 -7744 20954 -7738
rect 20920 -7772 20954 -7744
rect 20920 -7812 20939 -7811
rect 20939 -7812 20954 -7811
rect 20920 -7845 20954 -7812
rect 20920 -7914 20954 -7884
rect 20920 -7918 20939 -7914
rect 20939 -7918 20954 -7914
rect 20920 -7982 20954 -7957
rect 20920 -7991 20939 -7982
rect 20939 -7991 20954 -7982
rect 20920 -8050 20954 -8030
rect 20920 -8064 20939 -8050
rect 20939 -8064 20954 -8050
rect 16119 -8160 16153 -8138
rect 16119 -8172 16153 -8160
rect 16119 -8228 16153 -8210
rect 16119 -8244 16153 -8228
rect 16119 -8296 16153 -8282
rect 16119 -8316 16153 -8296
rect 16119 -8364 16153 -8354
rect 16119 -8388 16153 -8364
rect 16119 -8432 16153 -8426
rect 16119 -8460 16153 -8432
rect 16119 -8500 16153 -8498
rect 16119 -8532 16153 -8500
rect 16119 -8602 16153 -8570
rect 16119 -8604 16153 -8602
rect 16119 -8670 16153 -8642
rect 16119 -8676 16153 -8670
rect 20920 -8118 20954 -8103
rect 20920 -8137 20939 -8118
rect 20939 -8137 20954 -8118
rect 20920 -8186 20954 -8176
rect 20920 -8210 20939 -8186
rect 20939 -8210 20954 -8186
rect 20920 -8254 20954 -8249
rect 20920 -8283 20939 -8254
rect 20939 -8283 20954 -8254
rect 16119 -8738 16153 -8714
rect 17873 -8714 17907 -8680
rect 17949 -8714 17983 -8680
rect 18025 -8714 18059 -8680
rect 18101 -8714 18135 -8680
rect 18177 -8714 18211 -8680
rect 18254 -8714 18288 -8680
rect 18331 -8714 18365 -8680
rect 18408 -8714 18442 -8680
rect 18485 -8714 18519 -8680
rect 16119 -8748 16153 -8738
rect 16119 -8806 16153 -8787
rect 16119 -8821 16153 -8806
rect 16119 -8874 16153 -8860
rect 16119 -8894 16153 -8874
rect 16119 -8942 16153 -8933
rect 16119 -8967 16153 -8942
rect 16119 -9010 16153 -9006
rect 16119 -9040 16153 -9010
rect 16119 -9112 16153 -9079
rect 16119 -9113 16153 -9112
rect 16119 -9180 16153 -9152
rect 16119 -9186 16153 -9180
rect 16119 -9248 16153 -9225
rect 16119 -9259 16153 -9248
rect 18757 -9259 18791 -9225
rect 18829 -9227 18863 -9225
rect 18829 -9259 18830 -9227
rect 18830 -9259 18863 -9227
rect 19747 -9261 19764 -9227
rect 19764 -9261 19781 -9227
rect 19819 -9261 19840 -9227
rect 19840 -9261 19853 -9227
rect 16119 -9316 16153 -9298
rect 16119 -9332 16153 -9316
rect 16119 -9384 16153 -9371
rect 16119 -9405 16153 -9384
rect 16119 -9452 16153 -9444
rect 16119 -9478 16153 -9452
rect 16119 -9520 16153 -9517
rect 16119 -9551 16153 -9520
rect 16119 -9622 16153 -9590
rect 18769 -9321 18803 -9305
rect 18769 -9339 18803 -9321
rect 18769 -9389 18803 -9377
rect 18769 -9411 18803 -9389
rect 18769 -9457 18803 -9449
rect 18769 -9483 18803 -9457
rect 18925 -9321 18959 -9305
rect 18925 -9339 18959 -9321
rect 18925 -9389 18959 -9377
rect 18925 -9411 18959 -9389
rect 18925 -9457 18959 -9449
rect 18925 -9483 18959 -9457
rect 19081 -9321 19115 -9305
rect 19081 -9339 19115 -9321
rect 19081 -9389 19115 -9377
rect 19081 -9411 19115 -9389
rect 19081 -9457 19115 -9449
rect 19081 -9483 19115 -9457
rect 19475 -9361 19509 -9335
rect 19475 -9369 19509 -9361
rect 19475 -9429 19509 -9407
rect 19475 -9441 19509 -9429
rect 19475 -9497 19509 -9479
rect 19475 -9513 19509 -9497
rect 19631 -9361 19665 -9335
rect 19631 -9369 19665 -9361
rect 19631 -9429 19665 -9407
rect 19631 -9441 19665 -9429
rect 19631 -9497 19665 -9479
rect 19631 -9513 19665 -9497
rect 19787 -9361 19821 -9335
rect 19787 -9369 19821 -9361
rect 19787 -9429 19821 -9407
rect 19787 -9441 19821 -9429
rect 19787 -9497 19821 -9479
rect 19787 -9513 19821 -9497
rect 19910 -9327 19944 -9309
rect 19910 -9343 19932 -9327
rect 19932 -9343 19944 -9327
rect 19910 -9395 19944 -9381
rect 19910 -9415 19932 -9395
rect 19932 -9415 19944 -9395
rect 20054 -9327 20088 -9324
rect 20054 -9358 20088 -9327
rect 20763 -8356 20781 -8322
rect 20781 -8356 20797 -8322
rect 20848 -8356 20849 -8322
rect 20849 -8356 20882 -8322
rect 20679 -8417 20713 -8394
rect 20679 -8428 20713 -8417
rect 20679 -8485 20713 -8468
rect 20679 -8502 20713 -8485
rect 20679 -8553 20713 -8542
rect 20679 -8576 20713 -8553
rect 20679 -8621 20713 -8616
rect 20679 -8650 20713 -8621
rect 20679 -8723 20713 -8690
rect 20679 -8724 20713 -8723
rect 20679 -8791 20713 -8764
rect 20679 -8798 20713 -8791
rect 20679 -8859 20713 -8838
rect 20679 -8872 20713 -8859
rect 20679 -8927 20713 -8912
rect 20679 -8946 20713 -8927
rect 20679 -8995 20713 -8986
rect 20679 -9020 20713 -8995
rect 20679 -9063 20713 -9060
rect 20679 -9094 20713 -9063
rect 20679 -9165 20713 -9134
rect 20679 -9168 20713 -9165
rect 20679 -9233 20713 -9208
rect 20679 -9242 20713 -9233
rect 20679 -9301 20713 -9282
rect 20679 -9316 20713 -9301
rect 20054 -9429 20088 -9396
rect 20054 -9430 20088 -9429
rect 20679 -9369 20713 -9356
rect 20679 -9390 20713 -9369
rect 20679 -9437 20713 -9430
rect 20679 -9464 20713 -9437
rect 20679 -9505 20713 -9504
rect 16119 -9624 16153 -9622
rect 16119 -9690 16153 -9663
rect 16119 -9697 16153 -9690
rect 16119 -9758 16153 -9736
rect 16119 -9770 16153 -9758
rect 16119 -9843 16153 -9809
rect 16119 -9902 16153 -9882
rect 16119 -9916 16153 -9902
rect 16119 -9970 16153 -9955
rect 16119 -9989 16153 -9970
rect 16119 -10038 16153 -10028
rect 16119 -10062 16153 -10038
rect 16119 -10106 16153 -10101
rect 16119 -10135 16153 -10106
rect 18349 -10074 18383 -10040
rect 18349 -10131 18383 -10112
rect 18349 -10146 18383 -10131
rect 16119 -10208 16153 -10174
rect 20679 -9538 20713 -9505
rect 20250 -9584 20284 -9550
rect 20250 -9656 20284 -9622
rect 20412 -9627 20446 -9593
rect 20330 -9711 20364 -9677
rect 20412 -9699 20446 -9665
rect 20679 -9607 20713 -9578
rect 20679 -9612 20713 -9607
rect 20679 -9675 20713 -9652
rect 20679 -9686 20713 -9675
rect 20330 -9783 20364 -9749
rect 20679 -9743 20713 -9726
rect 20679 -9760 20713 -9743
rect 20679 -9811 20713 -9800
rect 20679 -9834 20713 -9811
rect 20679 -9879 20713 -9874
rect 20679 -9908 20713 -9879
rect 20679 -9981 20713 -9948
rect 20679 -9982 20713 -9981
rect 20250 -10074 20284 -10040
rect 20250 -10146 20284 -10112
rect 20679 -10049 20713 -10022
rect 20679 -10056 20713 -10049
rect 20679 -10117 20713 -10096
rect 20679 -10130 20713 -10117
rect 16119 -10276 16153 -10247
rect 16119 -10281 16153 -10276
rect 16634 -10233 16668 -10199
rect 17222 -10229 17256 -10195
rect 17294 -10229 17328 -10195
rect 20679 -10185 20713 -10170
rect 20679 -10204 20713 -10185
rect 16119 -10344 16153 -10320
rect 16119 -10354 16153 -10344
rect 16553 -10313 16587 -10279
rect 16634 -10305 16668 -10271
rect 16999 -10277 17031 -10243
rect 17031 -10277 17033 -10243
rect 17071 -10277 17099 -10243
rect 17099 -10277 17105 -10243
rect 20679 -10253 20713 -10244
rect 20679 -10278 20713 -10253
rect 16553 -10385 16587 -10351
rect 16715 -10313 16749 -10279
rect 17240 -10317 17274 -10315
rect 17327 -10317 17361 -10315
rect 17414 -10317 17448 -10315
rect 16715 -10385 16749 -10351
rect 17240 -10349 17242 -10317
rect 17242 -10349 17274 -10317
rect 17327 -10349 17344 -10317
rect 17344 -10349 17361 -10317
rect 17414 -10349 17446 -10317
rect 17446 -10349 17448 -10317
rect 18246 -10349 18280 -10315
rect 18318 -10349 18352 -10315
rect 20679 -10321 20713 -10318
rect 16119 -10412 16153 -10393
rect 16119 -10427 16153 -10412
rect 16979 -10404 16985 -10371
rect 16985 -10404 17013 -10371
rect 17063 -10404 17067 -10371
rect 17067 -10404 17097 -10371
rect 16979 -10405 17013 -10404
rect 17063 -10405 17097 -10404
rect 16119 -10480 16153 -10466
rect 16119 -10500 16153 -10480
rect 16119 -10548 16153 -10539
rect 16119 -10573 16153 -10548
rect 16478 -10483 16512 -10449
rect 16979 -10472 16985 -10443
rect 16985 -10472 17013 -10443
rect 17063 -10472 17067 -10443
rect 17067 -10472 17097 -10443
rect 17541 -10412 17574 -10395
rect 17574 -10412 17575 -10395
rect 17541 -10429 17575 -10412
rect 16979 -10477 17013 -10472
rect 17063 -10477 17097 -10472
rect 17222 -10473 17256 -10468
rect 17294 -10473 17328 -10468
rect 17222 -10502 17242 -10473
rect 17242 -10502 17256 -10473
rect 17294 -10502 17310 -10473
rect 17310 -10502 17328 -10473
rect 17541 -10480 17574 -10467
rect 17574 -10480 17575 -10467
rect 17541 -10501 17575 -10480
rect 17812 -10450 17846 -10424
rect 17812 -10458 17846 -10450
rect 16478 -10555 16512 -10521
rect 17812 -10518 17846 -10496
rect 17812 -10530 17846 -10518
rect 20679 -10352 20713 -10321
rect 20679 -10423 20713 -10392
rect 18736 -10450 18758 -10424
rect 18758 -10450 18770 -10424
rect 18736 -10458 18770 -10450
rect 18736 -10518 18758 -10496
rect 18758 -10518 18770 -10496
rect 18736 -10530 18770 -10518
rect 20679 -10426 20713 -10423
rect 20679 -10491 20713 -10465
rect 22415 -10478 22443 -10444
rect 22443 -10478 22449 -10444
rect 22492 -10478 22526 -10444
rect 22569 -10478 22588 -10444
rect 22588 -10478 22603 -10444
rect 22646 -10478 22680 -10444
rect 22723 -10478 22733 -10444
rect 22733 -10478 22757 -10444
rect 22800 -10478 22834 -10444
rect 22877 -10478 22878 -10444
rect 22878 -10478 22911 -10444
rect 22954 -10478 22988 -10444
rect 23031 -10478 23057 -10444
rect 23057 -10478 23065 -10444
rect 23108 -10478 23142 -10444
rect 23185 -10478 23202 -10444
rect 23202 -10478 23219 -10444
rect 23261 -10478 23295 -10444
rect 23337 -10478 23347 -10444
rect 23347 -10478 23371 -10444
rect 23413 -10478 23447 -10444
rect 23489 -10478 23492 -10444
rect 23492 -10478 23523 -10444
rect 23565 -10478 23599 -10444
rect 20679 -10499 20713 -10491
rect 20679 -10559 20713 -10538
rect 20679 -10572 20713 -10559
rect 16119 -10616 16153 -10612
rect 16119 -10646 16153 -10616
rect 16635 -10609 16669 -10575
rect 17919 -10612 17945 -10578
rect 17945 -10612 17953 -10578
rect 17998 -10612 18017 -10578
rect 18017 -10612 18032 -10578
rect 18077 -10612 18089 -10578
rect 18089 -10612 18111 -10578
rect 18156 -10612 18161 -10578
rect 18161 -10612 18190 -10578
rect 18235 -10612 18267 -10578
rect 18267 -10612 18269 -10578
rect 18314 -10612 18339 -10578
rect 18339 -10612 18348 -10578
rect 18393 -10612 18411 -10578
rect 18411 -10612 18427 -10578
rect 18471 -10612 18483 -10578
rect 18483 -10612 18505 -10578
rect 18549 -10612 18555 -10578
rect 18555 -10612 18583 -10578
rect 18627 -10612 18661 -10578
rect 18705 -10612 18739 -10578
rect 16635 -10681 16669 -10647
rect 20679 -10627 20713 -10611
rect 20679 -10645 20713 -10627
rect 16119 -10718 16153 -10685
rect 16119 -10719 16153 -10718
rect 16119 -10786 16153 -10758
rect 16800 -10709 16834 -10675
rect 16800 -10781 16834 -10747
rect 20679 -10695 20713 -10684
rect 20679 -10718 20713 -10695
rect 20679 -10763 20713 -10757
rect 16119 -10792 16153 -10786
rect 16119 -10854 16153 -10831
rect 16119 -10865 16153 -10854
rect 16119 -10922 16153 -10904
rect 16119 -10938 16153 -10922
rect 16119 -10990 16153 -10977
rect 16119 -11011 16153 -10990
rect 16119 -11058 16153 -11050
rect 16119 -11084 16153 -11058
rect 16119 -11126 16153 -11123
rect 16119 -11157 16153 -11126
rect 16119 -11228 16153 -11196
rect 16119 -11230 16153 -11228
rect 16119 -11296 16153 -11269
rect 16119 -11303 16153 -11296
rect 20679 -10791 20713 -10763
rect 20679 -10831 20713 -10830
rect 20679 -10864 20713 -10831
rect 22724 -10807 22758 -10773
rect 22724 -10879 22758 -10845
rect 22905 -10807 22939 -10773
rect 22905 -10879 22939 -10845
rect 23072 -10864 23106 -10830
rect 20679 -10933 20713 -10903
rect 20679 -10937 20713 -10933
rect 20679 -11001 20713 -10976
rect 20679 -11010 20713 -11001
rect 20679 -11069 20713 -11049
rect 23072 -10936 23106 -10902
rect 23174 -10922 23208 -10888
rect 23246 -10922 23280 -10888
rect 20679 -11083 20713 -11069
rect 20679 -11137 20713 -11122
rect 20679 -11156 20713 -11137
rect 22458 -11103 22492 -11069
rect 22458 -11175 22492 -11141
rect 22548 -11103 22582 -11069
rect 22548 -11175 22582 -11141
rect 22810 -11103 22844 -11069
rect 22810 -11175 22844 -11141
rect 22904 -11096 22938 -11062
rect 22904 -11168 22938 -11134
rect 23069 -11098 23103 -11064
rect 23069 -11170 23103 -11136
rect 23254 -11098 23288 -11064
rect 23254 -11170 23288 -11136
rect 23426 -11103 23460 -11069
rect 23426 -11175 23460 -11141
rect 23514 -11103 23548 -11069
rect 23514 -11175 23548 -11141
rect 20679 -11205 20713 -11195
rect 20679 -11229 20713 -11205
rect 20679 -11273 20713 -11268
rect 20679 -11302 20713 -11273
rect 16191 -11375 16221 -11341
rect 16221 -11375 16225 -11341
rect 16263 -11375 16289 -11341
rect 16289 -11375 16297 -11341
rect 16335 -11375 16357 -11341
rect 16357 -11375 16369 -11341
rect 16407 -11375 16425 -11341
rect 16425 -11375 16441 -11341
rect 16479 -11375 16493 -11341
rect 16493 -11375 16513 -11341
rect 16551 -11375 16561 -11341
rect 16561 -11375 16585 -11341
rect 16623 -11375 16629 -11341
rect 16629 -11375 16657 -11341
rect 16695 -11375 16697 -11341
rect 16697 -11375 16729 -11341
rect 16767 -11375 16799 -11341
rect 16799 -11375 16801 -11341
rect 16839 -11375 16867 -11341
rect 16867 -11375 16873 -11341
rect 16911 -11375 16935 -11341
rect 16935 -11375 16945 -11341
rect 16983 -11375 17003 -11341
rect 17003 -11375 17017 -11341
rect 17055 -11375 17071 -11341
rect 17071 -11375 17089 -11341
rect 17127 -11375 17139 -11341
rect 17139 -11375 17161 -11341
rect 17199 -11375 17207 -11341
rect 17207 -11375 17233 -11341
rect 17271 -11375 17275 -11341
rect 17275 -11375 17305 -11341
rect 17343 -11375 17377 -11341
rect 17415 -11375 17445 -11341
rect 17445 -11375 17449 -11341
rect 17487 -11375 17513 -11341
rect 17513 -11375 17521 -11341
rect 17559 -11375 17581 -11341
rect 17581 -11375 17593 -11341
rect 17631 -11375 17649 -11341
rect 17649 -11375 17665 -11341
rect 17703 -11375 17717 -11341
rect 17717 -11375 17737 -11341
rect 17775 -11375 17785 -11341
rect 17785 -11375 17809 -11341
rect 17847 -11375 17853 -11341
rect 17853 -11375 17881 -11341
rect 17919 -11375 17921 -11341
rect 17921 -11375 17953 -11341
rect 17991 -11375 18023 -11341
rect 18023 -11375 18025 -11341
rect 18063 -11375 18091 -11341
rect 18091 -11375 18097 -11341
rect 18135 -11375 18159 -11341
rect 18159 -11375 18169 -11341
rect 18207 -11375 18227 -11341
rect 18227 -11375 18241 -11341
rect 18279 -11375 18295 -11341
rect 18295 -11375 18313 -11341
rect 18351 -11375 18363 -11341
rect 18363 -11375 18385 -11341
rect 18423 -11375 18431 -11341
rect 18431 -11375 18457 -11341
rect 18495 -11375 18499 -11341
rect 18499 -11375 18529 -11341
rect 18567 -11375 18601 -11341
rect 18639 -11375 18669 -11341
rect 18669 -11375 18673 -11341
rect 18711 -11375 18737 -11341
rect 18737 -11375 18745 -11341
rect 18783 -11375 18805 -11341
rect 18805 -11375 18817 -11341
rect 18855 -11375 18873 -11341
rect 18873 -11375 18889 -11341
rect 18928 -11375 18941 -11341
rect 18941 -11375 18962 -11341
rect 19001 -11375 19009 -11341
rect 19009 -11375 19035 -11341
rect 19074 -11375 19077 -11341
rect 19077 -11375 19108 -11341
rect 19147 -11375 19179 -11341
rect 19179 -11375 19181 -11341
rect 19220 -11375 19247 -11341
rect 19247 -11375 19254 -11341
rect 19293 -11375 19315 -11341
rect 19315 -11375 19327 -11341
rect 19366 -11375 19383 -11341
rect 19383 -11375 19400 -11341
rect 19439 -11375 19451 -11341
rect 19451 -11375 19473 -11341
rect 19512 -11375 19519 -11341
rect 19519 -11375 19546 -11341
rect 19585 -11375 19587 -11341
rect 19587 -11375 19619 -11341
rect 19658 -11375 19689 -11341
rect 19689 -11375 19692 -11341
rect 19731 -11375 19757 -11341
rect 19757 -11375 19765 -11341
rect 19804 -11375 19825 -11341
rect 19825 -11375 19838 -11341
rect 19877 -11375 19893 -11341
rect 19893 -11375 19911 -11341
rect 19950 -11375 19961 -11341
rect 19961 -11375 19984 -11341
rect 20023 -11375 20029 -11341
rect 20029 -11375 20057 -11341
rect 20096 -11375 20097 -11341
rect 20097 -11375 20130 -11341
rect 20169 -11375 20199 -11341
rect 20199 -11375 20203 -11341
rect 20242 -11375 20267 -11341
rect 20267 -11375 20276 -11341
rect 20315 -11375 20335 -11341
rect 20335 -11375 20349 -11341
rect 20388 -11375 20403 -11341
rect 20403 -11375 20422 -11341
rect 20461 -11375 20471 -11341
rect 20471 -11375 20495 -11341
rect 20534 -11375 20539 -11341
rect 20539 -11375 20568 -11341
rect 20607 -11375 20641 -11341
rect 22494 -11466 22528 -11432
rect 22567 -11466 22598 -11432
rect 22598 -11466 22601 -11432
rect 22640 -11466 22667 -11432
rect 22667 -11466 22674 -11432
rect 22713 -11466 22736 -11432
rect 22736 -11466 22747 -11432
rect 22786 -11466 22805 -11432
rect 22805 -11466 22820 -11432
rect 22859 -11466 22874 -11432
rect 22874 -11466 22893 -11432
rect 22932 -11466 22943 -11432
rect 22943 -11466 22966 -11432
rect 23005 -11466 23012 -11432
rect 23012 -11466 23039 -11432
rect 23078 -11466 23081 -11432
rect 23081 -11466 23112 -11432
rect 23151 -11466 23184 -11432
rect 23184 -11466 23185 -11432
rect 23224 -11466 23253 -11432
rect 23253 -11466 23258 -11432
rect 23297 -11466 23322 -11432
rect 23322 -11466 23331 -11432
rect 23369 -11466 23391 -11432
rect 23391 -11466 23403 -11432
rect 23441 -11466 23460 -11432
rect 23460 -11466 23475 -11432
rect 23513 -11466 23529 -11432
rect 23529 -11466 23547 -11432
rect 23585 -11466 23598 -11432
rect 23598 -11466 23619 -11432
rect 23657 -11466 23667 -11432
rect 23667 -11466 23691 -11432
rect 23729 -11466 23736 -11432
rect 23736 -11466 23763 -11432
rect 23801 -11466 23805 -11432
rect 23805 -11466 23835 -11432
rect 23873 -11466 23874 -11432
rect 23874 -11466 23907 -11432
rect 23945 -11466 23978 -11432
rect 23978 -11466 23979 -11432
rect 24017 -11466 24047 -11432
rect 24047 -11466 24051 -11432
rect 24089 -11466 24116 -11432
rect 24116 -11466 24123 -11432
rect 24161 -11466 24185 -11432
rect 24185 -11466 24195 -11432
rect 24233 -11466 24254 -11432
rect 24254 -11466 24267 -11432
rect 24305 -11466 24323 -11432
rect 24323 -11466 24339 -11432
rect 24377 -11466 24392 -11432
rect 24392 -11466 24411 -11432
rect 24449 -11466 24461 -11432
rect 24461 -11466 24483 -11432
rect 24521 -11466 24530 -11432
rect 24530 -11466 24555 -11432
rect 24593 -11466 24599 -11432
rect 24599 -11466 24627 -11432
rect 24665 -11466 24668 -11432
rect 24668 -11466 24699 -11432
rect 24737 -11466 24771 -11432
rect 24809 -11466 24840 -11432
rect 24840 -11466 24843 -11432
rect 24881 -11466 24909 -11432
rect 24909 -11466 24915 -11432
rect 24953 -11466 24978 -11432
rect 24978 -11466 24987 -11432
rect 25025 -11466 25047 -11432
rect 25047 -11466 25059 -11432
rect 25097 -11466 25116 -11432
rect 25116 -11466 25131 -11432
rect 25169 -11466 25185 -11432
rect 25185 -11466 25203 -11432
rect 25241 -11466 25254 -11432
rect 25254 -11466 25275 -11432
rect 25313 -11466 25323 -11432
rect 25323 -11466 25347 -11432
rect 25385 -11466 25392 -11432
rect 25392 -11466 25419 -11432
rect 25457 -11466 25461 -11432
rect 25461 -11466 25491 -11432
rect 25529 -11466 25530 -11432
rect 25530 -11466 25563 -11432
rect 25601 -11466 25634 -11432
rect 25634 -11466 25635 -11432
rect 25673 -11466 25703 -11432
rect 25703 -11466 25707 -11432
rect 25745 -11466 25772 -11432
rect 25772 -11466 25779 -11432
rect 25817 -11466 25841 -11432
rect 25841 -11466 25851 -11432
rect 25889 -11466 25910 -11432
rect 25910 -11466 25923 -11432
rect 25961 -11466 25979 -11432
rect 25979 -11466 25995 -11432
rect 26033 -11466 26048 -11432
rect 26048 -11466 26067 -11432
rect 26105 -11466 26117 -11432
rect 26117 -11466 26139 -11432
rect 26177 -11466 26186 -11432
rect 26186 -11466 26211 -11432
rect 26249 -11466 26283 -11432
<< metal1 >>
rect 16434 -4653 16462 -4625
rect 17004 -6616 17056 -6610
rect 17004 -6680 17056 -6668
tri 16238 -6692 16244 -6686 se
rect 16244 -6692 16250 -6686
rect 16113 -6698 16250 -6692
rect 16302 -6698 16314 -6686
rect 16113 -6732 16191 -6698
rect 16225 -6732 16250 -6698
rect 16305 -6732 16314 -6698
rect 16113 -6738 16250 -6732
rect 16302 -6738 16314 -6732
rect 16366 -6738 16372 -6686
tri 17056 -6692 17090 -6658 sw
tri 17392 -6692 17426 -6658 se
rect 17472 -6692 17498 -6684
tri 17498 -6692 17506 -6684 nw
tri 17472 -6718 17498 -6692 nw
rect 17004 -6738 17056 -6732
rect 16113 -6770 16159 -6738
rect 16113 -6804 16119 -6770
rect 16153 -6804 16159 -6770
tri 16159 -6772 16193 -6738 nw
rect 16113 -6842 16159 -6804
rect 16113 -6876 16119 -6842
rect 16153 -6876 16159 -6842
rect 16113 -6914 16159 -6876
rect 16113 -6948 16119 -6914
rect 16153 -6948 16159 -6914
rect 16113 -6986 16159 -6948
rect 16113 -7020 16119 -6986
rect 16153 -7020 16159 -6986
rect 16113 -7058 16159 -7020
rect 20221 -6966 20273 -6960
rect 20221 -7030 20273 -7018
rect 16113 -7092 16119 -7058
rect 16153 -7092 16159 -7058
rect 18358 -7089 18386 -7061
rect 18463 -7089 18469 -7037
rect 18521 -7089 18533 -7037
rect 18585 -7089 18591 -7037
rect 20221 -7088 20273 -7082
rect 20388 -7089 20416 -7061
rect 16113 -7130 16159 -7092
rect 16113 -7164 16119 -7130
rect 16153 -7164 16159 -7130
rect 16113 -7202 16159 -7164
rect 16113 -7236 16119 -7202
rect 16153 -7236 16159 -7202
rect 16113 -7274 16159 -7236
rect 18575 -7261 18581 -7209
rect 18633 -7261 18645 -7209
rect 18697 -7261 18703 -7209
rect 20065 -7261 20071 -7209
rect 20123 -7261 20135 -7209
rect 20187 -7261 20193 -7209
rect 20914 -7225 20960 -7213
rect 20914 -7259 20920 -7225
rect 20954 -7259 20960 -7225
rect 16113 -7308 16119 -7274
rect 16153 -7308 16159 -7274
rect 16113 -7346 16159 -7308
rect 16113 -7380 16119 -7346
rect 16153 -7380 16159 -7346
rect 16113 -7418 16159 -7380
rect 18343 -7292 18395 -7286
rect 20914 -7299 20960 -7259
rect 18343 -7356 18395 -7344
rect 18343 -7414 18395 -7408
rect 18543 -7316 18595 -7310
rect 19240 -7356 19499 -7310
rect 18543 -7380 18595 -7368
rect 16113 -7452 16119 -7418
rect 16153 -7452 16159 -7418
rect 20049 -7402 20179 -7354
rect 20404 -7359 20410 -7307
rect 20462 -7359 20474 -7307
rect 20526 -7359 20532 -7307
rect 20914 -7333 20920 -7299
rect 20954 -7333 20960 -7299
rect 20049 -7428 20057 -7402
rect 18543 -7438 18595 -7432
rect 16113 -7490 16159 -7452
rect 20051 -7454 20057 -7428
rect 20109 -7454 20121 -7402
rect 20173 -7454 20179 -7402
rect 20914 -7373 20960 -7333
rect 20914 -7407 20920 -7373
rect 20954 -7407 20960 -7373
rect 21068 -7310 21120 -7304
rect 21068 -7374 21120 -7362
rect 20914 -7446 20960 -7407
rect 16113 -7524 16119 -7490
rect 16153 -7524 16159 -7490
rect 16113 -7562 16159 -7524
rect 16113 -7596 16119 -7562
rect 16153 -7596 16159 -7562
rect 16113 -7634 16159 -7596
rect 16113 -7668 16119 -7634
rect 16153 -7668 16159 -7634
rect 20914 -7480 20920 -7446
rect 20954 -7480 20960 -7446
rect 20914 -7519 20960 -7480
rect 20914 -7553 20920 -7519
rect 20954 -7553 20960 -7519
rect 20988 -7409 21040 -7403
rect 21068 -7432 21120 -7426
rect 20988 -7473 21040 -7461
rect 20988 -7531 21040 -7525
rect 20914 -7592 20960 -7553
rect 20914 -7626 20920 -7592
rect 20954 -7626 20960 -7592
rect 20914 -7665 20960 -7626
rect 16113 -7706 16159 -7668
rect 16113 -7740 16119 -7706
rect 16153 -7740 16159 -7706
rect 17577 -7718 17583 -7666
rect 17635 -7718 17647 -7666
rect 17699 -7718 18909 -7666
rect 18961 -7718 18973 -7666
rect 19025 -7718 19031 -7666
rect 20914 -7699 20920 -7665
rect 20954 -7699 20960 -7665
tri 19549 -7738 19566 -7721 se
rect 19566 -7738 20102 -7721
tri 20102 -7738 20119 -7721 sw
rect 16113 -7778 16159 -7740
tri 19541 -7746 19549 -7738 se
rect 19549 -7746 20119 -7738
tri 20119 -7746 20127 -7738 sw
rect 20587 -7746 20593 -7721
rect 16113 -7812 16119 -7778
rect 16153 -7812 16159 -7778
rect 16113 -7850 16159 -7812
rect 16113 -7884 16119 -7850
rect 16153 -7884 16159 -7850
rect 16113 -7922 16159 -7884
rect 16113 -7956 16119 -7922
rect 16153 -7956 16159 -7922
rect 16678 -7749 20593 -7746
rect 16678 -7772 19596 -7749
tri 19596 -7772 19619 -7749 nw
tri 20049 -7772 20072 -7749 ne
rect 20072 -7772 20593 -7749
rect 16678 -7774 19594 -7772
tri 19594 -7774 19596 -7772 nw
tri 20072 -7774 20074 -7772 ne
rect 20074 -7773 20593 -7772
rect 20645 -7773 20657 -7721
rect 20709 -7773 20715 -7721
rect 20074 -7774 20715 -7773
rect 20914 -7738 20960 -7699
rect 20914 -7772 20920 -7738
rect 20954 -7772 20960 -7738
rect 16678 -7805 16730 -7774
tri 16730 -7808 16764 -7774 nw
tri 19621 -7802 19646 -7777 se
rect 19646 -7802 19993 -7777
tri 19993 -7802 20018 -7777 sw
rect 16778 -7805 20593 -7802
rect 16778 -7808 19696 -7805
tri 19696 -7808 19699 -7805 nw
tri 19940 -7808 19943 -7805 ne
rect 19943 -7808 20593 -7805
rect 16678 -7869 16730 -7857
rect 16678 -7927 16730 -7921
rect 16830 -7811 19693 -7808
tri 19693 -7811 19696 -7808 nw
tri 19943 -7811 19946 -7808 ne
rect 19946 -7811 20593 -7808
rect 16830 -7830 19674 -7811
tri 19674 -7830 19693 -7811 nw
tri 19946 -7830 19965 -7811 ne
rect 19965 -7830 20593 -7811
rect 16830 -7833 16861 -7830
tri 16861 -7833 16864 -7830 nw
rect 16830 -7845 16849 -7833
tri 16849 -7845 16861 -7833 nw
tri 19707 -7845 19719 -7833 se
rect 19719 -7845 19725 -7833
rect 16830 -7858 16836 -7845
tri 16836 -7858 16849 -7845 nw
tri 19694 -7858 19707 -7845 se
rect 19707 -7858 19725 -7845
rect 16778 -7872 16830 -7860
tri 16830 -7864 16836 -7858 nw
tri 16883 -7864 16889 -7858 se
rect 16889 -7864 19725 -7858
tri 16863 -7884 16883 -7864 se
rect 16883 -7884 19725 -7864
tri 16862 -7885 16863 -7884 se
rect 16863 -7885 19725 -7884
rect 19777 -7885 19789 -7833
rect 19841 -7885 19847 -7833
rect 20587 -7854 20593 -7830
rect 20645 -7854 20657 -7802
rect 20709 -7854 20715 -7802
rect 20914 -7811 20960 -7772
rect 20914 -7845 20920 -7811
rect 20954 -7845 20960 -7811
rect 20914 -7884 20960 -7845
rect 16778 -7930 16830 -7924
tri 16858 -7889 16862 -7885 se
rect 16862 -7886 19827 -7885
rect 16862 -7889 16909 -7886
tri 16909 -7889 16912 -7886 nw
rect 16113 -7994 16159 -7956
rect 16113 -8028 16119 -7994
rect 16153 -8028 16159 -7994
rect 16113 -8066 16159 -8028
rect 16113 -8100 16119 -8066
rect 16153 -8100 16159 -8066
rect 16113 -8138 16159 -8100
rect 16453 -7991 16505 -7985
tri 16505 -8030 16534 -8001 sw
tri 16829 -8030 16858 -8001 se
rect 16858 -8030 16886 -7889
tri 16886 -7912 16909 -7889 nw
tri 17104 -7916 17106 -7914 se
rect 17106 -7916 17574 -7914
rect 16505 -8035 16534 -8030
tri 16534 -8035 16539 -8030 sw
tri 16824 -8035 16829 -8030 se
rect 16829 -8035 16886 -8030
rect 16505 -8043 16886 -8035
rect 16453 -8055 16886 -8043
rect 16505 -8063 16886 -8055
rect 16922 -7922 17574 -7916
rect 16974 -7974 17008 -7922
rect 17060 -7974 17574 -7922
rect 16922 -7987 17574 -7974
rect 16974 -8039 17008 -7987
rect 17060 -8039 17574 -7987
rect 16922 -8052 17574 -8039
rect 16505 -8064 16538 -8063
tri 16538 -8064 16539 -8063 nw
rect 16505 -8092 16510 -8064
tri 16510 -8092 16538 -8064 nw
tri 16505 -8097 16510 -8092 nw
rect 16453 -8113 16505 -8107
rect 16974 -8104 17008 -8052
rect 17060 -8104 17574 -8052
rect 16922 -8111 17574 -8104
rect 17868 -7918 18071 -7917
rect 17868 -7970 17874 -7918
rect 17926 -7970 17944 -7918
rect 17996 -7970 18013 -7918
rect 18065 -7970 18071 -7918
rect 17868 -7988 18071 -7970
rect 17868 -8040 17874 -7988
rect 17926 -8040 17944 -7988
rect 17996 -8040 18013 -7988
rect 18065 -8040 18071 -7988
rect 17868 -8058 18071 -8040
rect 17868 -8110 17874 -8058
rect 17926 -8110 17944 -8058
rect 17996 -8110 18013 -8058
rect 18065 -8110 18071 -8058
rect 17868 -8111 18071 -8110
rect 18334 -8111 19106 -7914
rect 19327 -8111 19493 -7914
rect 20914 -7918 20920 -7884
rect 20954 -7918 20960 -7884
rect 20914 -7957 20960 -7918
rect 20914 -7991 20920 -7957
rect 20954 -7991 20960 -7957
rect 20914 -8030 20960 -7991
rect 20914 -8064 20920 -8030
rect 20954 -8064 20960 -8030
rect 20914 -8103 20960 -8064
rect 16113 -8172 16119 -8138
rect 16153 -8172 16159 -8138
rect 20914 -8137 20920 -8103
rect 20954 -8137 20960 -8103
rect 16113 -8210 16159 -8172
rect 16113 -8244 16119 -8210
rect 16153 -8244 16159 -8210
rect 16113 -8282 16159 -8244
rect 16113 -8316 16119 -8282
rect 16153 -8316 16159 -8282
rect 16113 -8354 16159 -8316
rect 16239 -8343 16389 -8141
rect 18128 -8147 18330 -8141
rect 18128 -8199 18129 -8147
rect 18181 -8199 18203 -8147
rect 18255 -8199 18277 -8147
rect 18329 -8199 18330 -8147
rect 18128 -8216 18330 -8199
rect 18128 -8268 18129 -8216
rect 18181 -8268 18203 -8216
rect 18255 -8268 18277 -8216
rect 18329 -8268 18330 -8216
rect 18128 -8285 18330 -8268
rect 18128 -8337 18129 -8285
rect 18181 -8337 18203 -8285
rect 18255 -8337 18277 -8285
rect 18329 -8337 18330 -8285
rect 18128 -8343 18330 -8337
rect 19994 -8142 20314 -8141
rect 19994 -8194 20000 -8142
rect 20052 -8194 20086 -8142
rect 20138 -8194 20171 -8142
rect 20223 -8194 20256 -8142
rect 20308 -8194 20314 -8142
rect 19994 -8216 20314 -8194
rect 19994 -8268 20000 -8216
rect 20052 -8268 20086 -8216
rect 20138 -8268 20171 -8216
rect 20223 -8268 20256 -8216
rect 20308 -8268 20314 -8216
rect 19994 -8290 20314 -8268
rect 19994 -8342 20000 -8290
rect 20052 -8342 20086 -8290
rect 20138 -8342 20171 -8290
rect 20223 -8342 20256 -8290
rect 20308 -8342 20314 -8290
rect 20914 -8176 20960 -8137
rect 20914 -8210 20920 -8176
rect 20954 -8210 20960 -8176
rect 20914 -8249 20960 -8210
rect 20914 -8283 20920 -8249
rect 20954 -8283 20960 -8249
rect 20914 -8316 20960 -8283
rect 19994 -8343 20314 -8342
rect 20673 -8322 20960 -8316
rect 16113 -8388 16119 -8354
rect 16153 -8388 16159 -8354
rect 20673 -8356 20763 -8322
rect 20797 -8356 20848 -8322
rect 20882 -8356 20960 -8322
rect 20673 -8362 20960 -8356
rect 16113 -8426 16159 -8388
rect 16113 -8460 16119 -8426
rect 16153 -8460 16159 -8426
rect 16113 -8498 16159 -8460
rect 16113 -8532 16119 -8498
rect 16153 -8532 16159 -8498
rect 17697 -8383 17749 -8377
rect 17697 -8447 17749 -8435
rect 17697 -8505 17749 -8499
rect 18682 -8383 18734 -8377
rect 18682 -8447 18734 -8435
rect 18682 -8505 18734 -8499
rect 20673 -8394 20719 -8362
rect 20673 -8428 20679 -8394
rect 20713 -8428 20719 -8394
rect 20673 -8468 20719 -8428
rect 20673 -8502 20679 -8468
rect 20713 -8502 20719 -8468
rect 16113 -8570 16159 -8532
rect 16113 -8604 16119 -8570
rect 16153 -8604 16159 -8570
rect 16113 -8642 16159 -8604
rect 16113 -8676 16119 -8642
rect 16153 -8676 16159 -8642
rect 20673 -8542 20719 -8502
rect 20673 -8576 20679 -8542
rect 20713 -8576 20719 -8542
rect 20673 -8616 20719 -8576
rect 16113 -8714 16159 -8676
rect 16515 -8696 16521 -8644
rect 16573 -8696 16585 -8644
rect 16637 -8696 16643 -8644
rect 17861 -8680 18531 -8674
rect 16113 -8748 16119 -8714
rect 16153 -8748 16159 -8714
rect 17408 -8733 17414 -8681
rect 17466 -8733 17478 -8681
rect 17530 -8733 17536 -8681
rect 17779 -8689 17831 -8683
rect 16113 -8787 16159 -8748
rect 16520 -8786 16526 -8734
rect 16578 -8786 16590 -8734
rect 16642 -8786 16648 -8734
rect 17861 -8714 17873 -8680
rect 17907 -8714 17949 -8680
rect 17983 -8714 18025 -8680
rect 18059 -8714 18101 -8680
rect 18135 -8714 18177 -8680
rect 18211 -8714 18254 -8680
rect 18288 -8714 18331 -8680
rect 18365 -8714 18408 -8680
rect 18442 -8714 18485 -8680
rect 18519 -8714 18531 -8680
rect 17861 -8720 18531 -8714
rect 18910 -8727 18916 -8675
rect 18968 -8727 18981 -8675
rect 19033 -8727 19039 -8675
tri 19039 -8681 19045 -8675 sw
rect 19763 -8696 19769 -8644
rect 19821 -8696 19833 -8644
rect 19885 -8696 19891 -8644
rect 20673 -8650 20679 -8616
rect 20713 -8650 20719 -8616
rect 20673 -8690 20719 -8650
rect 20673 -8724 20679 -8690
rect 20713 -8724 20719 -8690
rect 16113 -8821 16119 -8787
rect 16153 -8821 16159 -8787
rect 16751 -8803 16757 -8751
rect 16809 -8803 16821 -8751
rect 16873 -8803 16879 -8751
rect 17779 -8753 17831 -8741
rect 17779 -8811 17831 -8805
rect 17985 -8811 18438 -8765
rect 19609 -8792 19637 -8764
rect 19824 -8772 19852 -8744
rect 20673 -8764 20719 -8724
rect 20673 -8798 20679 -8764
rect 20713 -8798 20719 -8764
rect 16113 -8860 16159 -8821
rect 16113 -8894 16119 -8860
rect 16153 -8894 16159 -8860
rect 16113 -8933 16159 -8894
rect 16113 -8967 16119 -8933
rect 16153 -8967 16159 -8933
rect 20673 -8838 20719 -8798
rect 20673 -8872 20679 -8838
rect 20713 -8872 20719 -8838
rect 20673 -8912 20719 -8872
rect 20673 -8946 20679 -8912
rect 20713 -8946 20719 -8912
rect 16113 -9006 16159 -8967
rect 16113 -9040 16119 -9006
rect 16153 -9040 16159 -9006
rect 16113 -9079 16159 -9040
rect 16113 -9113 16119 -9079
rect 16153 -9113 16159 -9079
rect 16113 -9152 16159 -9113
rect 16113 -9186 16119 -9152
rect 16153 -9186 16159 -9152
rect 16113 -9225 16159 -9186
rect 16113 -9259 16119 -9225
rect 16153 -9259 16159 -9225
rect 16113 -9298 16159 -9259
rect 16113 -9332 16119 -9298
rect 16153 -9332 16159 -9298
rect 16909 -9003 17061 -8997
rect 16961 -9055 17009 -9003
rect 16909 -9083 17061 -9055
rect 16961 -9135 17009 -9083
rect 16909 -9164 17061 -9135
rect 16961 -9216 17009 -9164
rect 16909 -9245 17061 -9216
rect 16961 -9297 17009 -9245
rect 16909 -9303 17061 -9297
rect 17869 -9003 18071 -8997
rect 17869 -9055 17870 -9003
rect 17922 -9055 17944 -9003
rect 17996 -9055 18018 -9003
rect 18070 -9055 18071 -9003
rect 17869 -9083 18071 -9055
rect 17869 -9135 17870 -9083
rect 17922 -9135 17944 -9083
rect 17996 -9135 18018 -9083
rect 18070 -9135 18071 -9083
rect 17869 -9164 18071 -9135
rect 17869 -9216 17870 -9164
rect 17922 -9216 17944 -9164
rect 17996 -9216 18018 -9164
rect 18070 -9216 18071 -9164
rect 17869 -9245 18071 -9216
rect 17869 -9297 17870 -9245
rect 17922 -9297 17944 -9245
rect 17996 -9297 18018 -9245
rect 18070 -9297 18071 -9245
rect 17869 -9303 18071 -9297
rect 18160 -9178 18263 -8964
rect 20673 -8986 20719 -8946
rect 20673 -9020 20679 -8986
rect 20713 -9020 20719 -8986
rect 18415 -9073 18487 -9045
rect 20673 -9060 20719 -9020
rect 20673 -9094 20679 -9060
rect 20713 -9094 20719 -9060
rect 20673 -9134 20719 -9094
rect 20673 -9168 20679 -9134
rect 20713 -9168 20719 -9134
rect 16113 -9371 16159 -9332
rect 18160 -9336 18396 -9178
rect 18627 -9220 18875 -9219
rect 16113 -9405 16119 -9371
rect 16153 -9405 16159 -9371
rect 16113 -9444 16159 -9405
rect 16113 -9478 16119 -9444
rect 16153 -9478 16159 -9444
rect 16113 -9517 16159 -9478
rect 17779 -9495 17831 -9489
rect 16113 -9551 16119 -9517
rect 16153 -9551 16159 -9517
rect 16113 -9590 16159 -9551
rect 16520 -9565 16526 -9513
rect 16578 -9565 16590 -9513
rect 16642 -9565 16648 -9513
rect 16751 -9548 16757 -9496
rect 16809 -9548 16821 -9496
rect 16873 -9548 16879 -9496
rect 17779 -9559 17831 -9547
rect 16113 -9624 16119 -9590
rect 16153 -9624 16159 -9590
rect 16113 -9663 16159 -9624
rect 16515 -9656 16521 -9604
rect 16573 -9656 16585 -9604
rect 16637 -9656 16643 -9604
rect 17409 -9622 17415 -9570
rect 17467 -9622 17479 -9570
rect 17531 -9622 17537 -9570
rect 17779 -9617 17831 -9611
rect 18230 -9598 18396 -9336
rect 18602 -9225 18875 -9220
rect 18602 -9226 18757 -9225
rect 18654 -9259 18757 -9226
rect 18791 -9259 18829 -9225
rect 18863 -9259 18875 -9225
rect 18654 -9265 18875 -9259
rect 18602 -9290 18654 -9278
rect 18602 -9348 18654 -9342
rect 18763 -9305 18809 -9293
rect 18763 -9339 18769 -9305
rect 18803 -9339 18809 -9305
rect 18763 -9365 18809 -9339
rect 18919 -9305 18965 -9174
rect 18919 -9339 18925 -9305
rect 18959 -9339 18965 -9305
rect 18763 -9371 18815 -9365
rect 18763 -9435 18815 -9423
rect 18763 -9493 18815 -9487
rect 18919 -9377 18965 -9339
rect 18919 -9411 18925 -9377
rect 18959 -9411 18965 -9377
rect 18919 -9449 18965 -9411
rect 18919 -9483 18925 -9449
rect 18959 -9483 18965 -9449
rect 18763 -9495 18809 -9493
rect 18919 -9495 18965 -9483
rect 19075 -9299 19161 -9293
rect 19075 -9305 19109 -9299
rect 19075 -9339 19081 -9305
rect 19075 -9351 19109 -9339
rect 19075 -9368 19161 -9351
rect 19075 -9377 19109 -9368
rect 19075 -9411 19081 -9377
rect 19469 -9335 19515 -9323
rect 19469 -9369 19475 -9335
rect 19509 -9369 19515 -9335
rect 19469 -9393 19515 -9369
rect 19075 -9420 19109 -9411
rect 19075 -9437 19161 -9420
rect 19075 -9449 19109 -9437
rect 19075 -9483 19081 -9449
rect 19075 -9489 19109 -9483
rect 19075 -9495 19161 -9489
rect 19454 -9399 19515 -9393
rect 19506 -9407 19515 -9399
rect 19509 -9441 19515 -9407
rect 19506 -9451 19515 -9441
rect 19454 -9463 19515 -9451
rect 19506 -9479 19515 -9463
rect 19509 -9513 19515 -9479
rect 19506 -9515 19515 -9513
rect 19454 -9521 19515 -9515
rect 19469 -9525 19515 -9521
rect 19625 -9335 19671 -9178
rect 19746 -9221 19752 -9216
rect 19735 -9227 19752 -9221
rect 19735 -9261 19747 -9227
rect 19735 -9267 19752 -9261
rect 19746 -9268 19752 -9267
rect 19804 -9268 19816 -9216
rect 19868 -9268 19874 -9216
rect 19904 -9309 19950 -9178
rect 20673 -9208 20719 -9168
rect 20673 -9242 20679 -9208
rect 20713 -9242 20719 -9208
rect 20673 -9282 20719 -9242
rect 19625 -9369 19631 -9335
rect 19665 -9369 19671 -9335
rect 19625 -9407 19671 -9369
rect 19781 -9335 19827 -9323
rect 19781 -9369 19787 -9335
rect 19821 -9369 19827 -9335
rect 19781 -9393 19827 -9369
rect 19625 -9441 19631 -9407
rect 19665 -9441 19671 -9407
rect 19625 -9479 19671 -9441
rect 19625 -9513 19631 -9479
rect 19665 -9513 19671 -9479
rect 19625 -9525 19671 -9513
rect 19775 -9399 19827 -9393
rect 19904 -9343 19910 -9309
rect 19944 -9343 19950 -9309
rect 19904 -9381 19950 -9343
rect 19904 -9415 19910 -9381
rect 19944 -9415 19950 -9381
rect 19904 -9427 19950 -9415
rect 20045 -9314 20097 -9308
rect 20045 -9384 20097 -9366
rect 20045 -9442 20097 -9436
rect 20673 -9316 20679 -9282
rect 20713 -9316 20719 -9282
rect 20673 -9356 20719 -9316
rect 20673 -9390 20679 -9356
rect 20713 -9390 20719 -9356
rect 20673 -9430 20719 -9390
rect 19775 -9467 19827 -9451
rect 19775 -9525 19827 -9519
rect 20673 -9464 20679 -9430
rect 20713 -9464 20719 -9430
rect 20673 -9504 20719 -9464
rect 20673 -9538 20679 -9504
rect 20713 -9538 20719 -9504
tri 20196 -9550 20208 -9538 se
rect 20208 -9550 20290 -9538
tri 20162 -9584 20196 -9550 se
rect 20196 -9584 20250 -9550
rect 20284 -9584 20290 -9550
rect 20673 -9578 20719 -9538
tri 20153 -9593 20162 -9584 se
rect 20162 -9593 20290 -9584
tri 20148 -9598 20153 -9593 se
rect 20153 -9598 20290 -9593
rect 16113 -9697 16119 -9663
rect 16153 -9697 16159 -9663
rect 16113 -9736 16159 -9697
rect 18230 -9728 18582 -9598
rect 19286 -9728 19410 -9598
rect 19556 -9604 19678 -9598
rect 19608 -9656 19626 -9604
rect 19556 -9670 19678 -9656
rect 19608 -9722 19626 -9670
rect 19556 -9728 19678 -9722
rect 20036 -9622 20290 -9598
rect 20036 -9656 20250 -9622
rect 20284 -9656 20290 -9622
rect 20036 -9728 20290 -9656
rect 20406 -9593 20452 -9581
rect 20406 -9627 20412 -9593
rect 20446 -9627 20452 -9593
rect 20406 -9665 20452 -9627
rect 20322 -9671 20374 -9665
rect 20406 -9699 20412 -9665
rect 20446 -9699 20452 -9665
rect 20406 -9711 20452 -9699
rect 20673 -9612 20679 -9578
rect 20713 -9612 20719 -9578
rect 20673 -9652 20719 -9612
rect 20673 -9686 20679 -9652
rect 20713 -9686 20719 -9652
rect 16113 -9770 16119 -9736
rect 16153 -9770 16159 -9736
rect 20322 -9735 20374 -9723
rect 16113 -9809 16159 -9770
rect 18763 -9766 18815 -9760
rect 16113 -9843 16119 -9809
rect 16153 -9834 16159 -9809
rect 18053 -9800 18125 -9790
tri 18125 -9800 18135 -9790 sw
rect 18053 -9806 18135 -9800
tri 18135 -9806 18141 -9800 sw
tri 16159 -9834 16167 -9826 sw
rect 18053 -9834 18141 -9806
tri 18141 -9834 18169 -9806 sw
rect 18763 -9830 18815 -9818
rect 16153 -9836 16167 -9834
tri 16167 -9836 16169 -9834 sw
rect 18053 -9836 18169 -9834
rect 16153 -9843 16169 -9836
rect 16113 -9861 16169 -9843
tri 16169 -9861 16194 -9836 sw
tri 18116 -9861 18141 -9836 ne
rect 18141 -9861 18169 -9836
tri 18169 -9861 18196 -9834 sw
rect 16113 -9874 16194 -9861
tri 16194 -9874 16207 -9861 sw
tri 18141 -9874 18154 -9861 ne
rect 18154 -9874 18196 -9861
tri 18196 -9874 18209 -9861 sw
rect 16113 -9882 16207 -9874
rect 16113 -9916 16119 -9882
rect 16153 -9908 16207 -9882
tri 16207 -9908 16241 -9874 sw
tri 18154 -9908 18188 -9874 ne
rect 18188 -9888 18209 -9874
tri 18209 -9888 18223 -9874 sw
rect 19109 -9764 19161 -9758
rect 19109 -9828 19161 -9816
rect 18763 -9888 18815 -9882
tri 18899 -9886 18903 -9882 sw
rect 19109 -9886 19161 -9880
rect 19251 -9759 19367 -9758
rect 19251 -9765 19407 -9759
rect 19251 -9817 19355 -9765
rect 19251 -9829 19407 -9817
rect 19251 -9881 19355 -9829
rect 18899 -9888 18903 -9886
tri 18903 -9888 18905 -9886 sw
rect 19251 -9887 19407 -9881
rect 19454 -9766 19506 -9760
rect 19454 -9830 19506 -9818
rect 19251 -9888 19367 -9887
rect 19454 -9888 19506 -9882
rect 19775 -9764 19827 -9758
rect 20322 -9793 20374 -9787
rect 20673 -9726 20719 -9686
rect 20673 -9760 20679 -9726
rect 20713 -9760 20719 -9726
rect 20324 -9795 20370 -9793
rect 19775 -9828 19827 -9816
rect 19775 -9886 19827 -9880
rect 20673 -9800 20719 -9760
rect 20673 -9834 20679 -9800
rect 20713 -9834 20719 -9800
rect 20673 -9874 20719 -9834
rect 18188 -9908 18223 -9888
tri 18223 -9908 18243 -9888 sw
tri 18835 -9908 18853 -9890 se
rect 18853 -9908 18905 -9888
tri 18905 -9908 18925 -9888 sw
rect 16153 -9916 16241 -9908
tri 16241 -9916 16249 -9908 sw
tri 18188 -9916 18196 -9908 ne
rect 18196 -9916 18243 -9908
tri 18243 -9916 18251 -9908 sw
tri 18827 -9916 18835 -9908 se
rect 18835 -9916 18925 -9908
tri 18925 -9916 18933 -9908 sw
rect 19909 -9916 19955 -9888
rect 16113 -9944 16249 -9916
tri 16249 -9944 16277 -9916 sw
tri 18196 -9944 18224 -9916 ne
rect 18224 -9944 19955 -9916
rect 20673 -9908 20679 -9874
rect 20713 -9908 20719 -9874
rect 16113 -9948 16277 -9944
tri 16277 -9948 16281 -9944 sw
rect 20673 -9948 20719 -9908
rect 16113 -9955 16281 -9948
rect 16113 -9989 16119 -9955
rect 16153 -9957 16281 -9955
tri 16281 -9957 16290 -9948 sw
rect 16153 -9989 16389 -9957
rect 16113 -10028 16389 -9989
tri 18155 -9982 18180 -9957 sw
rect 20673 -9982 20679 -9948
rect 20713 -9982 20719 -9948
rect 18155 -9992 18180 -9982
tri 18180 -9992 18190 -9982 sw
rect 16113 -10062 16119 -10028
rect 16153 -10062 16389 -10028
rect 16113 -10101 16389 -10062
rect 16113 -10135 16119 -10101
rect 16153 -10135 16389 -10101
rect 16585 -9998 16637 -9992
rect 18155 -10022 18190 -9992
tri 18190 -10022 18220 -9992 sw
rect 20673 -10022 20719 -9982
rect 18155 -10028 18220 -10022
tri 18220 -10028 18226 -10022 sw
rect 16585 -10062 16637 -10050
rect 17464 -10079 17492 -10051
rect 16585 -10120 16637 -10114
rect 18127 -10080 18133 -10028
rect 18185 -10080 18198 -10028
rect 18250 -10080 18262 -10028
rect 18314 -10040 19410 -10028
rect 18314 -10074 18349 -10040
rect 18383 -10074 19410 -10040
rect 18314 -10080 19410 -10074
rect 18127 -10106 19410 -10080
rect 16113 -10159 16389 -10135
rect 18127 -10158 18133 -10106
rect 18185 -10158 18198 -10106
rect 18250 -10158 18262 -10106
rect 18314 -10112 19410 -10106
rect 18314 -10146 18349 -10112
rect 18383 -10146 19410 -10112
rect 18314 -10158 19410 -10146
rect 19994 -10080 20000 -10028
rect 20052 -10080 20086 -10028
rect 20138 -10080 20171 -10028
rect 20223 -10040 20256 -10028
rect 20223 -10074 20250 -10040
rect 20223 -10080 20256 -10074
rect 20308 -10080 20314 -10028
rect 19994 -10106 20314 -10080
rect 19994 -10158 20000 -10106
rect 20052 -10158 20086 -10106
rect 20138 -10158 20171 -10106
rect 20223 -10112 20256 -10106
rect 20223 -10146 20250 -10112
rect 20223 -10158 20256 -10146
rect 20308 -10158 20314 -10106
rect 20673 -10056 20679 -10022
rect 20713 -10056 20719 -10022
rect 20673 -10096 20719 -10056
rect 20673 -10130 20679 -10096
rect 20713 -10130 20719 -10096
rect 18155 -10159 18343 -10158
tri 18343 -10159 18344 -10158 nw
rect 16113 -10170 16258 -10159
tri 16258 -10170 16269 -10159 nw
rect 20673 -10170 20719 -10130
rect 16113 -10174 16233 -10170
rect 16113 -10208 16119 -10174
rect 16153 -10195 16233 -10174
tri 16233 -10195 16258 -10170 nw
rect 16628 -10193 18067 -10187
rect 16153 -10199 16229 -10195
tri 16229 -10199 16233 -10195 nw
rect 16628 -10199 16936 -10193
rect 16153 -10208 16195 -10199
rect 16113 -10233 16195 -10208
tri 16195 -10233 16229 -10199 nw
rect 16628 -10233 16634 -10199
rect 16668 -10233 16936 -10199
rect 16113 -10243 16185 -10233
tri 16185 -10243 16195 -10233 nw
rect 16628 -10243 16693 -10233
tri 16693 -10243 16703 -10233 nw
tri 16902 -10243 16912 -10233 ne
rect 16912 -10243 16936 -10233
rect 16113 -10247 16181 -10243
tri 16181 -10247 16185 -10243 nw
rect 16113 -10281 16119 -10247
rect 16153 -10281 16159 -10247
tri 16159 -10269 16181 -10247 nw
rect 16113 -10320 16159 -10281
rect 16113 -10354 16119 -10320
rect 16153 -10354 16159 -10320
rect 16113 -10393 16159 -10354
rect 16113 -10427 16119 -10393
rect 16153 -10427 16159 -10393
rect 16113 -10466 16159 -10427
rect 16547 -10279 16593 -10267
rect 16547 -10313 16553 -10279
rect 16587 -10313 16593 -10279
rect 16547 -10351 16593 -10313
rect 16628 -10271 16674 -10243
tri 16674 -10262 16693 -10243 nw
tri 16912 -10262 16931 -10243 ne
rect 16931 -10245 16936 -10243
rect 16988 -10243 17010 -10193
rect 17062 -10195 18067 -10193
rect 17062 -10229 17222 -10195
rect 17256 -10229 17294 -10195
rect 17328 -10208 18067 -10195
rect 19890 -10201 19896 -10195
tri 19186 -10204 19189 -10201 se
rect 19189 -10204 19896 -10201
rect 17328 -10229 17874 -10208
rect 17062 -10243 17874 -10229
rect 16988 -10245 16999 -10243
rect 17062 -10245 17071 -10243
rect 16931 -10262 16999 -10245
tri 16931 -10267 16936 -10262 ne
rect 16628 -10305 16634 -10271
rect 16668 -10305 16674 -10271
rect 16628 -10317 16674 -10305
rect 16709 -10273 16869 -10267
rect 16709 -10279 16817 -10273
rect 16709 -10313 16715 -10279
rect 16749 -10313 16817 -10279
rect 16547 -10385 16553 -10351
rect 16587 -10385 16593 -10351
rect 16547 -10427 16593 -10385
rect 16709 -10325 16817 -10313
rect 16709 -10339 16869 -10325
rect 16709 -10351 16817 -10339
rect 16709 -10385 16715 -10351
rect 16749 -10385 16817 -10351
rect 16709 -10391 16817 -10385
rect 16709 -10397 16869 -10391
rect 16936 -10277 16999 -10262
rect 17033 -10277 17071 -10245
rect 17105 -10260 17874 -10243
rect 17926 -10260 17942 -10208
rect 17994 -10260 18009 -10208
rect 18061 -10260 18067 -10208
tri 19146 -10244 19186 -10204 se
rect 19186 -10244 19896 -10204
tri 19143 -10247 19146 -10244 se
rect 19146 -10247 19896 -10244
rect 19948 -10247 19960 -10195
rect 20012 -10247 20018 -10195
rect 20673 -10204 20679 -10170
rect 20713 -10204 20719 -10170
rect 20673 -10244 20719 -10204
rect 17105 -10277 18067 -10260
tri 19123 -10267 19143 -10247 se
rect 19143 -10267 19189 -10247
tri 19189 -10267 19209 -10247 nw
tri 19121 -10269 19123 -10267 se
rect 19123 -10269 19178 -10267
rect 16936 -10278 18067 -10277
tri 19112 -10278 19121 -10269 se
rect 19121 -10278 19178 -10269
tri 19178 -10278 19189 -10267 nw
rect 20673 -10278 20679 -10244
rect 20713 -10278 20719 -10244
rect 16988 -10330 17010 -10278
rect 17062 -10281 18067 -10278
tri 19109 -10281 19112 -10278 se
rect 19112 -10281 19147 -10278
rect 17062 -10309 17156 -10281
tri 17156 -10309 17184 -10281 nw
tri 19081 -10309 19109 -10281 se
rect 19109 -10309 19147 -10281
tri 19147 -10309 19178 -10278 nw
rect 17062 -10315 17150 -10309
tri 17150 -10315 17156 -10309 nw
rect 17228 -10315 19138 -10309
rect 17062 -10330 17137 -10315
tri 17137 -10328 17150 -10315 nw
rect 16936 -10364 17137 -10330
rect 17228 -10349 17240 -10315
rect 17274 -10349 17327 -10315
rect 17361 -10349 17414 -10315
rect 17448 -10349 18246 -10315
rect 18280 -10349 18318 -10315
rect 18352 -10318 19138 -10315
tri 19138 -10318 19147 -10309 nw
rect 20673 -10318 20719 -10278
rect 18352 -10349 19104 -10318
rect 17228 -10352 19104 -10349
tri 19104 -10352 19138 -10318 nw
rect 20673 -10352 20679 -10318
rect 20713 -10352 20719 -10318
rect 17228 -10354 19102 -10352
tri 19102 -10354 19104 -10352 nw
rect 17228 -10355 18195 -10354
tri 18195 -10355 18196 -10354 nw
tri 18233 -10355 18234 -10354 ne
rect 18234 -10355 18364 -10354
tri 18364 -10355 18365 -10354 nw
rect 16988 -10371 17010 -10364
rect 17062 -10371 17137 -10364
rect 17062 -10405 17063 -10371
rect 17097 -10405 17137 -10371
tri 17323 -10392 17360 -10355 ne
rect 17360 -10392 17406 -10355
tri 17406 -10392 17443 -10355 nw
tri 17360 -10395 17363 -10392 ne
rect 17363 -10395 17403 -10392
tri 17403 -10395 17406 -10392 nw
rect 17535 -10395 17581 -10383
tri 17363 -10401 17369 -10395 ne
rect 16988 -10416 17010 -10405
rect 17062 -10416 17137 -10405
tri 16547 -10429 16549 -10427 ne
rect 16549 -10429 16593 -10427
tri 16593 -10429 16603 -10419 sw
rect 16936 -10429 17137 -10416
tri 17137 -10429 17138 -10428 sw
tri 16549 -10437 16557 -10429 ne
rect 16557 -10437 16603 -10429
rect 16113 -10500 16119 -10466
rect 16153 -10500 16159 -10466
rect 16113 -10539 16159 -10500
rect 16113 -10573 16119 -10539
rect 16153 -10573 16159 -10539
rect 16472 -10449 16518 -10437
tri 16557 -10443 16563 -10437 ne
rect 16563 -10443 16603 -10437
tri 16603 -10443 16617 -10429 sw
rect 16936 -10443 17138 -10429
tri 16563 -10444 16564 -10443 ne
rect 16564 -10444 16617 -10443
tri 16617 -10444 16618 -10443 sw
rect 16472 -10483 16478 -10449
rect 16512 -10483 16518 -10449
tri 16564 -10457 16577 -10444 ne
rect 16577 -10457 16678 -10444
tri 16678 -10457 16691 -10444 sw
rect 16936 -10450 16979 -10443
rect 17013 -10450 17063 -10443
tri 16577 -10472 16592 -10457 ne
rect 16592 -10472 16691 -10457
tri 16662 -10477 16667 -10472 ne
rect 16667 -10477 16691 -10472
tri 16691 -10477 16711 -10457 sw
rect 17062 -10477 17063 -10450
rect 17097 -10444 17138 -10443
tri 17138 -10444 17153 -10429 sw
rect 17097 -10457 17153 -10444
tri 17153 -10457 17166 -10444 sw
rect 17097 -10458 17166 -10457
tri 17166 -10458 17167 -10457 sw
rect 17097 -10462 17167 -10458
tri 17167 -10462 17171 -10458 sw
rect 17097 -10468 17340 -10462
rect 17097 -10477 17222 -10468
rect 16472 -10521 16518 -10483
tri 16667 -10501 16691 -10477 ne
rect 16691 -10501 16711 -10477
tri 16711 -10501 16735 -10477 sw
tri 16691 -10502 16692 -10501 ne
rect 16692 -10502 16735 -10501
tri 16735 -10502 16736 -10501 sw
rect 16988 -10502 17010 -10477
rect 17062 -10502 17222 -10477
rect 17256 -10502 17294 -10468
rect 17328 -10502 17340 -10468
rect 16472 -10555 16478 -10521
rect 16512 -10555 16518 -10521
tri 16692 -10530 16720 -10502 ne
rect 16720 -10519 16736 -10502
tri 16736 -10519 16753 -10502 sw
rect 16936 -10508 17340 -10502
rect 16720 -10530 16753 -10519
tri 16753 -10530 16764 -10519 sw
tri 17358 -10530 17369 -10519 se
rect 17369 -10530 17397 -10395
tri 17397 -10401 17403 -10395 nw
tri 16720 -10538 16728 -10530 ne
rect 16728 -10538 16764 -10530
tri 16764 -10538 16772 -10530 sw
tri 17350 -10538 17358 -10530 se
rect 17358 -10538 17397 -10530
tri 16728 -10545 16735 -10538 ne
rect 16735 -10542 16772 -10538
tri 16772 -10542 16776 -10538 sw
tri 17346 -10542 17350 -10538 se
rect 17350 -10542 17397 -10538
rect 16735 -10545 16776 -10542
tri 16776 -10545 16779 -10542 sw
tri 17343 -10545 17346 -10542 se
rect 17346 -10545 17397 -10542
rect 16472 -10567 16518 -10555
tri 16735 -10563 16753 -10545 ne
rect 16753 -10553 17397 -10545
rect 16753 -10563 17379 -10553
rect 16113 -10612 16159 -10573
rect 16113 -10646 16119 -10612
rect 16153 -10646 16159 -10612
rect 16113 -10685 16159 -10646
rect 16113 -10719 16119 -10685
rect 16153 -10719 16159 -10685
rect 16585 -10569 16675 -10563
rect 16637 -10575 16675 -10569
tri 16753 -10571 16761 -10563 ne
rect 16761 -10571 17379 -10563
tri 17379 -10571 17397 -10553 nw
rect 17535 -10429 17541 -10395
rect 17575 -10429 17581 -10395
rect 20673 -10392 20719 -10352
rect 17535 -10467 17581 -10429
rect 17535 -10501 17541 -10467
rect 17575 -10501 17581 -10467
rect 17535 -10530 17581 -10501
rect 17806 -10424 18133 -10412
rect 17806 -10458 17812 -10424
rect 17846 -10458 18133 -10424
rect 17806 -10464 18133 -10458
rect 18185 -10464 18203 -10412
rect 18255 -10464 18272 -10412
rect 18324 -10424 20000 -10412
rect 18324 -10458 18736 -10424
rect 18770 -10458 20000 -10424
rect 18324 -10464 20000 -10458
rect 20052 -10464 20086 -10412
rect 20138 -10464 20171 -10412
rect 20223 -10464 20256 -10412
rect 20308 -10464 20355 -10412
rect 17806 -10486 20355 -10464
rect 17806 -10496 18133 -10486
tri 17581 -10530 17589 -10522 sw
rect 17806 -10530 17812 -10496
rect 17846 -10530 18133 -10496
rect 17535 -10538 17589 -10530
tri 17589 -10538 17597 -10530 sw
rect 17806 -10538 18133 -10530
rect 18185 -10538 18203 -10486
rect 18255 -10538 18272 -10486
rect 18324 -10490 20355 -10486
rect 18324 -10496 20000 -10490
rect 18324 -10530 18736 -10496
rect 18770 -10530 20000 -10496
rect 18324 -10538 20000 -10530
rect 17535 -10542 17597 -10538
tri 17597 -10542 17601 -10538 sw
rect 17806 -10542 20000 -10538
rect 20052 -10542 20086 -10490
rect 20138 -10542 20171 -10490
rect 20223 -10542 20256 -10490
rect 20308 -10542 20355 -10490
rect 20673 -10426 20679 -10392
rect 20713 -10426 20719 -10392
rect 20673 -10465 20719 -10426
rect 20673 -10499 20679 -10465
rect 20713 -10499 20719 -10465
rect 20673 -10538 20719 -10499
tri 17535 -10571 17564 -10542 ne
rect 17564 -10571 17601 -10542
tri 17601 -10571 17630 -10542 sw
tri 16761 -10572 16762 -10571 ne
rect 16762 -10572 17378 -10571
tri 17378 -10572 17379 -10571 nw
tri 17564 -10572 17565 -10571 ne
rect 17565 -10572 17630 -10571
tri 17630 -10572 17631 -10571 sw
tri 19097 -10572 19098 -10571 se
rect 19098 -10572 19678 -10571
tri 16762 -10573 16763 -10572 ne
rect 16763 -10573 17377 -10572
tri 17377 -10573 17378 -10572 nw
tri 17565 -10573 17566 -10572 ne
rect 17566 -10573 18644 -10572
rect 16669 -10609 16675 -10575
tri 17566 -10578 17571 -10573 ne
rect 17571 -10578 18644 -10573
rect 18696 -10578 18708 -10572
tri 17571 -10588 17581 -10578 ne
rect 17581 -10588 17919 -10578
rect 16637 -10621 16675 -10609
tri 17581 -10612 17605 -10588 ne
rect 17605 -10612 17919 -10588
rect 17953 -10612 17998 -10578
rect 18032 -10612 18077 -10578
rect 18111 -10612 18156 -10578
rect 18190 -10612 18235 -10578
rect 18269 -10612 18314 -10578
rect 18348 -10612 18393 -10578
rect 18427 -10612 18471 -10578
rect 18505 -10612 18549 -10578
rect 18583 -10612 18627 -10578
rect 18696 -10612 18705 -10578
tri 17605 -10618 17611 -10612 ne
rect 17611 -10618 18644 -10612
rect 16585 -10635 16675 -10621
rect 18638 -10624 18644 -10618
rect 18696 -10624 18708 -10612
rect 18760 -10624 18766 -10572
tri 19058 -10611 19097 -10572 se
rect 19097 -10577 19678 -10572
rect 19097 -10611 19556 -10577
tri 19045 -10624 19058 -10611 se
rect 19058 -10624 19556 -10611
rect 16637 -10647 16675 -10635
tri 19024 -10645 19045 -10624 se
rect 19045 -10629 19556 -10624
rect 19608 -10629 19626 -10577
rect 19045 -10643 19678 -10629
rect 19045 -10645 19556 -10643
rect 16669 -10681 16675 -10647
tri 19006 -10663 19024 -10645 se
rect 19024 -10663 19556 -10645
rect 16637 -10687 16675 -10681
rect 16585 -10693 16675 -10687
rect 16794 -10675 16840 -10663
rect 16113 -10758 16159 -10719
rect 16113 -10792 16119 -10758
rect 16153 -10792 16159 -10758
rect 16113 -10831 16159 -10792
rect 16794 -10709 16800 -10675
rect 16834 -10709 16840 -10675
tri 18988 -10681 19006 -10663 se
rect 19006 -10681 19556 -10663
rect 16794 -10747 16840 -10709
rect 16794 -10781 16800 -10747
rect 16834 -10781 16840 -10747
rect 16794 -10793 16840 -10781
rect 18127 -10733 18133 -10681
rect 18185 -10733 18200 -10681
rect 18252 -10733 18258 -10681
tri 18985 -10684 18988 -10681 se
rect 18988 -10684 19556 -10681
tri 18968 -10701 18985 -10684 se
rect 18985 -10695 19556 -10684
rect 19608 -10695 19626 -10643
rect 18985 -10701 19678 -10695
rect 20673 -10572 20679 -10538
rect 20713 -10572 20719 -10538
rect 20673 -10611 20719 -10572
rect 20673 -10645 20679 -10611
rect 20713 -10645 20719 -10611
rect 20673 -10684 20719 -10645
tri 18951 -10718 18968 -10701 se
rect 18968 -10718 19285 -10701
tri 19285 -10718 19302 -10701 nw
rect 20673 -10718 20679 -10684
rect 20713 -10718 20719 -10684
rect 18127 -10745 18258 -10733
tri 18926 -10743 18951 -10718 se
rect 18951 -10738 19260 -10718
rect 18951 -10743 19159 -10738
rect 19236 -10743 19260 -10738
tri 19260 -10743 19285 -10718 nw
rect 18127 -10791 18133 -10745
tri 17385 -10793 17387 -10791 ne
rect 17387 -10793 17419 -10791
tri 17387 -10807 17401 -10793 ne
rect 17401 -10807 17419 -10793
tri 17401 -10825 17419 -10807 ne
rect 17465 -10793 17497 -10791
tri 17497 -10793 17499 -10791 nw
tri 17925 -10793 17927 -10791 ne
rect 17927 -10793 17959 -10791
rect 17465 -10807 17483 -10793
tri 17483 -10807 17497 -10793 nw
tri 17927 -10807 17941 -10793 ne
rect 17941 -10807 17959 -10793
tri 17465 -10825 17483 -10807 nw
tri 17941 -10825 17959 -10807 ne
rect 18005 -10793 18037 -10791
tri 18037 -10793 18039 -10791 nw
tri 18121 -10793 18123 -10791 ne
rect 18123 -10793 18133 -10791
rect 18005 -10797 18033 -10793
tri 18033 -10797 18037 -10793 nw
tri 18123 -10797 18127 -10793 ne
rect 18127 -10797 18133 -10793
rect 18185 -10797 18200 -10745
rect 18252 -10797 18258 -10745
rect 19236 -10757 19246 -10743
tri 19246 -10757 19260 -10743 nw
rect 20673 -10757 20719 -10718
tri 19236 -10767 19246 -10757 nw
rect 20673 -10791 20679 -10757
rect 20713 -10791 20719 -10757
rect 18005 -10807 18023 -10797
tri 18023 -10807 18033 -10797 nw
rect 18005 -10811 18019 -10807
tri 18019 -10811 18023 -10807 nw
tri 18005 -10825 18019 -10811 nw
tri 18277 -10825 18291 -10811 se
tri 18272 -10830 18277 -10825 se
rect 18277 -10830 18291 -10825
rect 16113 -10865 16119 -10831
rect 16153 -10865 16159 -10831
tri 18257 -10845 18272 -10830 se
rect 18272 -10845 18291 -10830
rect 20673 -10830 20719 -10791
rect 16113 -10904 16159 -10865
rect 20673 -10864 20679 -10830
rect 20713 -10864 20719 -10830
tri 18389 -10900 18399 -10890 se
tri 18387 -10902 18389 -10900 se
rect 18389 -10902 18399 -10900
tri 18386 -10903 18387 -10902 se
rect 18387 -10903 18399 -10902
rect 16113 -10938 16119 -10904
rect 16153 -10938 16159 -10904
tri 18365 -10924 18386 -10903 se
rect 18386 -10924 18399 -10903
tri 18445 -10902 18447 -10900 sw
rect 18445 -10903 18447 -10902
tri 18447 -10903 18448 -10902 sw
rect 20673 -10903 20719 -10864
rect 18445 -10924 18448 -10903
tri 18448 -10924 18469 -10903 sw
rect 18445 -10934 18469 -10924
tri 18469 -10934 18479 -10924 sw
rect 16113 -10977 16159 -10938
rect 20673 -10937 20679 -10903
rect 20713 -10937 20719 -10903
tri 18389 -10976 18395 -10970 ne
rect 18395 -10976 18399 -10970
rect 16113 -11011 16119 -10977
rect 16153 -11011 16159 -10977
tri 18395 -10980 18399 -10976 ne
rect 20673 -10976 20719 -10937
tri 17797 -11010 17800 -11007 se
rect 17800 -11010 17801 -11007
rect 17927 -11010 17928 -11007
tri 17928 -11010 17931 -11007 sw
rect 20673 -11010 20679 -10976
rect 20713 -11010 20719 -10976
rect 16113 -11050 16159 -11011
rect 16113 -11084 16119 -11050
rect 16153 -11084 16159 -11050
rect 20673 -11049 20719 -11010
tri 17797 -11059 17800 -11056 ne
tri 17928 -11059 17931 -11056 nw
rect 18759 -11059 18790 -11056
tri 18790 -11059 18793 -11056 nw
rect 18759 -11070 18779 -11059
tri 18779 -11070 18790 -11059 nw
tri 18700 -11083 18713 -11070 se
rect 16113 -11123 16159 -11084
tri 18693 -11090 18700 -11083 se
rect 18700 -11090 18713 -11083
rect 18759 -11083 18766 -11070
tri 18766 -11083 18779 -11070 nw
rect 20673 -11083 20679 -11049
rect 20713 -11083 20719 -11049
tri 18759 -11090 18766 -11083 nw
tri 18680 -11103 18693 -11090 se
rect 18693 -11103 18713 -11090
tri 18679 -11104 18680 -11103 se
rect 18680 -11104 18713 -11103
rect 16113 -11157 16119 -11123
rect 16153 -11157 16159 -11123
rect 20673 -11122 20719 -11083
rect 18834 -11144 18854 -11130
tri 18854 -11144 18868 -11130 nw
tri 18794 -11156 18806 -11144 se
rect 16113 -11196 16159 -11157
tri 18786 -11164 18794 -11156 se
rect 18794 -11164 18806 -11156
rect 18834 -11156 18842 -11144
tri 18842 -11156 18854 -11144 nw
rect 20673 -11156 20679 -11122
rect 20713 -11156 20719 -11122
tri 18834 -11164 18842 -11156 nw
tri 18775 -11175 18786 -11164 se
rect 18786 -11175 18806 -11164
tri 18772 -11178 18775 -11175 se
rect 18775 -11178 18806 -11175
rect 16113 -11230 16119 -11196
rect 16153 -11230 16159 -11196
rect 16113 -11269 16159 -11230
rect 16113 -11303 16119 -11269
rect 16153 -11303 16159 -11269
rect 20673 -11195 20719 -11156
rect 20673 -11229 20679 -11195
rect 20713 -11229 20719 -11195
rect 20673 -11268 20719 -11229
tri 20672 -11302 20673 -11301 se
rect 20673 -11302 20679 -11268
rect 20713 -11302 20719 -11268
rect 16113 -11335 16159 -11303
tri 20642 -11332 20672 -11302 se
rect 20672 -11332 20719 -11302
tri 20093 -11335 20096 -11332 se
rect 20096 -11335 20102 -11332
rect 16113 -11341 20102 -11335
rect 20154 -11341 20180 -11332
rect 20232 -11341 20257 -11332
rect 20309 -11335 20315 -11332
tri 20315 -11335 20318 -11332 sw
tri 20639 -11335 20642 -11332 se
rect 20642 -11335 20719 -11332
rect 20309 -11341 20719 -11335
rect 16113 -11375 16191 -11341
rect 16225 -11375 16263 -11341
rect 16297 -11375 16335 -11341
rect 16369 -11375 16407 -11341
rect 16441 -11375 16479 -11341
rect 16513 -11375 16551 -11341
rect 16585 -11375 16623 -11341
rect 16657 -11375 16695 -11341
rect 16729 -11375 16767 -11341
rect 16801 -11375 16839 -11341
rect 16873 -11375 16911 -11341
rect 16945 -11375 16983 -11341
rect 17017 -11375 17055 -11341
rect 17089 -11375 17127 -11341
rect 17161 -11375 17199 -11341
rect 17233 -11375 17271 -11341
rect 17305 -11375 17343 -11341
rect 17377 -11375 17415 -11341
rect 17449 -11375 17487 -11341
rect 17521 -11375 17559 -11341
rect 17593 -11375 17631 -11341
rect 17665 -11375 17703 -11341
rect 17737 -11375 17775 -11341
rect 17809 -11375 17847 -11341
rect 17881 -11375 17919 -11341
rect 17953 -11375 17991 -11341
rect 18025 -11375 18063 -11341
rect 18097 -11375 18135 -11341
rect 18169 -11375 18207 -11341
rect 18241 -11375 18279 -11341
rect 18313 -11375 18351 -11341
rect 18385 -11375 18423 -11341
rect 18457 -11375 18495 -11341
rect 18529 -11375 18567 -11341
rect 18601 -11375 18639 -11341
rect 18673 -11375 18711 -11341
rect 18745 -11375 18783 -11341
rect 18817 -11375 18855 -11341
rect 18889 -11375 18928 -11341
rect 18962 -11375 19001 -11341
rect 19035 -11375 19074 -11341
rect 19108 -11375 19147 -11341
rect 19181 -11375 19220 -11341
rect 19254 -11375 19293 -11341
rect 19327 -11375 19366 -11341
rect 19400 -11375 19439 -11341
rect 19473 -11375 19512 -11341
rect 19546 -11375 19585 -11341
rect 19619 -11375 19658 -11341
rect 19692 -11375 19731 -11341
rect 19765 -11375 19804 -11341
rect 19838 -11375 19877 -11341
rect 19911 -11375 19950 -11341
rect 19984 -11375 20023 -11341
rect 20057 -11375 20096 -11341
rect 20154 -11375 20169 -11341
rect 20232 -11375 20242 -11341
rect 20309 -11375 20315 -11341
rect 20349 -11375 20388 -11341
rect 20422 -11375 20461 -11341
rect 20495 -11375 20534 -11341
rect 20568 -11375 20607 -11341
rect 20641 -11375 20719 -11341
rect 16113 -11381 20102 -11375
rect 17333 -11384 17404 -11381
tri 17404 -11384 17407 -11381 nw
tri 20093 -11384 20096 -11381 ne
rect 20096 -11384 20102 -11381
rect 20154 -11384 20180 -11375
rect 20232 -11384 20257 -11375
rect 20309 -11381 20719 -11375
rect 20309 -11384 20315 -11381
tri 20315 -11384 20318 -11381 nw
rect 17333 -11409 17379 -11384
tri 17379 -11409 17404 -11384 nw
rect 17333 -11432 17356 -11409
tri 17356 -11432 17379 -11409 nw
rect 17333 -11434 17354 -11432
tri 17354 -11434 17356 -11432 nw
rect 17685 -11461 17691 -11409
rect 17743 -11461 17755 -11409
rect 17807 -11461 19349 -11409
rect 19401 -11461 19413 -11409
rect 19465 -11461 19471 -11409
tri 19617 -11465 19618 -11464 se
rect 17059 -11466 17060 -11465
tri 17060 -11466 17061 -11465 sw
tri 19616 -11466 19617 -11465 se
rect 19617 -11466 19618 -11465
rect 17059 -11489 17061 -11466
tri 17061 -11489 17084 -11466 sw
tri 19593 -11489 19616 -11466 se
rect 19616 -11489 19618 -11466
tri 19746 -11466 19748 -11464 sw
rect 19746 -11489 19748 -11466
tri 19748 -11489 19771 -11466 sw
tri 19990 -11489 19993 -11486 se
rect 19993 -11489 19994 -11486
tri 19989 -11490 19990 -11489 se
rect 19990 -11490 19994 -11489
tri 19972 -11538 19993 -11517 ne
tri 16635 -11564 16636 -11563 sw
rect 16863 -11605 16869 -11553
rect 16921 -11605 16933 -11553
rect 16985 -11559 19827 -11553
rect 16985 -11581 19775 -11559
rect 16985 -11605 16991 -11581
tri 16991 -11604 17014 -11581 nw
tri 19741 -11604 19764 -11581 ne
rect 19764 -11604 19775 -11581
tri 19764 -11605 19765 -11604 ne
rect 19765 -11605 19775 -11604
tri 19765 -11610 19770 -11605 ne
rect 19770 -11610 19775 -11605
rect 16633 -11615 16635 -11610
tri 16635 -11615 16640 -11610 nw
tri 18090 -11615 18095 -11610 se
rect 18095 -11615 18105 -11610
tri 19770 -11615 19775 -11610 ne
tri 18081 -11624 18090 -11615 se
rect 18090 -11624 18105 -11615
rect 19775 -11623 19827 -11611
tri 18084 -11662 18095 -11651 ne
rect 18095 -11662 18101 -11651
rect 18222 -11662 18223 -11648
tri 18223 -11662 18237 -11648 nw
tri 19518 -11662 19532 -11648 ne
rect 19532 -11662 19534 -11648
tri 18355 -11689 18368 -11676 se
rect 18368 -11689 18374 -11676
rect 17473 -11695 17525 -11689
tri 17525 -11699 17535 -11689 sw
tri 18345 -11699 18355 -11689 se
rect 18355 -11699 18374 -11689
rect 17525 -11727 18374 -11699
rect 17525 -11728 17558 -11727
tri 17558 -11728 17559 -11727 nw
tri 18367 -11728 18368 -11727 ne
rect 18368 -11728 18374 -11727
rect 18426 -11728 18438 -11676
rect 18490 -11728 18496 -11676
rect 19775 -11681 19827 -11675
rect 17525 -11747 17530 -11728
rect 17473 -11756 17530 -11747
tri 17530 -11756 17558 -11728 nw
rect 17473 -11759 17525 -11756
tri 17525 -11761 17530 -11756 nw
tri 18479 -11761 18484 -11756 se
rect 18484 -11761 18490 -11756
tri 18478 -11762 18479 -11761 se
rect 18479 -11762 18490 -11761
rect 17473 -11817 17525 -11811
rect 17572 -11814 17578 -11762
rect 17630 -11814 17642 -11762
rect 17694 -11790 18490 -11762
rect 17694 -11808 17706 -11790
tri 17706 -11808 17724 -11790 nw
tri 18466 -11808 18484 -11790 ne
rect 18484 -11808 18490 -11790
rect 18542 -11808 18554 -11756
rect 18606 -11808 18612 -11756
rect 17694 -11814 17700 -11808
tri 17700 -11814 17706 -11808 nw
tri 17795 -11868 17819 -11844 se
rect 20992 -11873 21032 -7531
rect 21072 -11772 21112 -7432
rect 21236 -7710 21288 -7704
rect 21236 -7774 21288 -7762
rect 21147 -7808 21199 -7802
rect 21147 -7872 21199 -7860
rect 21147 -7930 21199 -7924
rect 21236 -7832 21288 -7826
rect 21160 -11715 21188 -7930
rect 21236 -11663 21264 -7832
tri 22737 -8633 22755 -8615 se
rect 22755 -8667 22761 -8615
rect 22813 -8667 22825 -8615
rect 22877 -8639 22883 -8615
tri 22883 -8639 22907 -8615 sw
tri 26749 -8639 26773 -8615 se
rect 26773 -8639 26774 -8615
rect 22877 -8664 25670 -8639
tri 25670 -8664 25695 -8639 sw
tri 26724 -8664 26749 -8639 se
rect 26749 -8664 26774 -8639
rect 22877 -8667 26906 -8664
tri 25585 -8696 25614 -8667 ne
rect 25614 -8696 26906 -8667
rect 23065 -8927 23299 -8904
rect 23065 -8979 23071 -8927
rect 23123 -8979 23156 -8927
rect 23208 -8979 23241 -8927
rect 23293 -8979 23299 -8927
rect 23065 -9002 23299 -8979
tri 23054 -9427 23088 -9393 sw
tri 22876 -9465 22910 -9431 se
rect 23402 -9873 23454 -9867
rect 23402 -9939 23454 -9925
rect 23402 -9997 23454 -9991
rect 23228 -10198 23234 -10146
rect 23286 -10198 23298 -10146
rect 23350 -10198 23356 -10146
tri 23356 -10151 23361 -10146 sw
tri 23356 -10198 23361 -10193 nw
rect 23054 -10259 23236 -10236
rect 23054 -10311 23060 -10259
rect 23112 -10311 23178 -10259
rect 23230 -10311 23236 -10259
rect 23054 -10334 23236 -10311
rect 22403 -10444 23685 -10438
rect 22403 -10478 22415 -10444
rect 22449 -10478 22492 -10444
rect 22526 -10478 22569 -10444
rect 22603 -10478 22646 -10444
rect 22680 -10478 22723 -10444
rect 22757 -10478 22800 -10444
rect 22834 -10478 22877 -10444
rect 22911 -10478 22954 -10444
rect 22988 -10478 23031 -10444
rect 23065 -10478 23108 -10444
rect 23142 -10478 23185 -10444
rect 23219 -10478 23261 -10444
rect 23295 -10478 23337 -10444
rect 23371 -10478 23413 -10444
rect 23447 -10478 23489 -10444
rect 23523 -10478 23565 -10444
rect 23599 -10478 23685 -10444
rect 22403 -10484 23685 -10478
rect 22906 -10546 22934 -10518
rect 22718 -10773 22764 -10761
rect 22718 -10807 22724 -10773
rect 22758 -10807 22764 -10773
rect 22718 -10845 22764 -10807
rect 22718 -10879 22724 -10845
rect 22758 -10879 22764 -10845
rect 22718 -10891 22764 -10879
rect 22899 -10773 22945 -10761
rect 22899 -10807 22905 -10773
rect 22939 -10807 22945 -10773
rect 22899 -10845 22945 -10807
rect 22899 -10879 22905 -10845
rect 22939 -10879 22945 -10845
rect 22899 -10891 22945 -10879
rect 23066 -10830 23112 -10818
rect 23066 -10864 23072 -10830
rect 23106 -10864 23112 -10830
rect 23066 -10902 23112 -10864
rect 23066 -10936 23072 -10902
rect 23106 -10936 23112 -10902
rect 23162 -10888 23466 -10882
rect 23162 -10922 23174 -10888
rect 23208 -10922 23246 -10888
rect 23280 -10922 23466 -10888
rect 23162 -10928 23466 -10922
rect 23066 -10948 23112 -10936
rect 22452 -11069 22498 -11057
rect 22452 -11103 22458 -11069
rect 22492 -11103 22498 -11069
rect 22452 -11141 22498 -11103
rect 22452 -11175 22458 -11141
rect 22492 -11175 22498 -11141
rect 22452 -11187 22498 -11175
rect 22542 -11069 22850 -11057
rect 22542 -11103 22548 -11069
rect 22582 -11103 22810 -11069
rect 22844 -11103 22850 -11069
rect 22542 -11141 22850 -11103
rect 22542 -11175 22548 -11141
rect 22582 -11175 22810 -11141
rect 22844 -11175 22850 -11141
rect 22542 -11187 22850 -11175
rect 22898 -11062 22944 -11050
rect 22898 -11096 22904 -11062
rect 22938 -11096 22944 -11062
rect 22898 -11134 22944 -11096
rect 22898 -11168 22904 -11134
rect 22938 -11168 22944 -11134
rect 22898 -11180 22944 -11168
rect 23063 -11064 23294 -11052
rect 23063 -11098 23069 -11064
rect 23103 -11098 23254 -11064
rect 23288 -11098 23294 -11064
rect 23063 -11136 23294 -11098
rect 23063 -11170 23069 -11136
rect 23103 -11170 23254 -11136
rect 23288 -11170 23294 -11136
rect 23063 -11182 23294 -11170
rect 23420 -11069 23466 -10928
rect 23420 -11103 23426 -11069
rect 23460 -11103 23466 -11069
rect 23420 -11141 23466 -11103
rect 23420 -11175 23426 -11141
rect 23460 -11175 23466 -11141
rect 23420 -11187 23466 -11175
rect 23508 -11069 23554 -11057
rect 23508 -11103 23514 -11069
rect 23548 -11103 23554 -11069
rect 23508 -11141 23554 -11103
rect 23508 -11175 23514 -11141
rect 23548 -11175 23554 -11141
rect 23508 -11187 23554 -11175
rect 23137 -11269 23253 -11263
rect 23189 -11321 23201 -11269
rect 22961 -11349 22989 -11321
rect 23137 -11344 23253 -11321
rect 23189 -11396 23201 -11344
rect 23137 -11420 23253 -11396
rect 22482 -11432 23137 -11426
rect 22482 -11466 22494 -11432
rect 22528 -11466 22567 -11432
rect 22601 -11466 22640 -11432
rect 22674 -11466 22713 -11432
rect 22747 -11466 22786 -11432
rect 22820 -11466 22859 -11432
rect 22893 -11466 22932 -11432
rect 22966 -11466 23005 -11432
rect 23039 -11466 23078 -11432
rect 23112 -11466 23137 -11432
rect 22482 -11472 23137 -11466
rect 23189 -11472 23201 -11420
rect 23253 -11432 26295 -11426
rect 23258 -11466 23297 -11432
rect 23331 -11466 23369 -11432
rect 23403 -11466 23441 -11432
rect 23475 -11466 23513 -11432
rect 23547 -11466 23585 -11432
rect 23619 -11466 23657 -11432
rect 23691 -11466 23729 -11432
rect 23763 -11466 23801 -11432
rect 23835 -11466 23873 -11432
rect 23907 -11466 23945 -11432
rect 23979 -11466 24017 -11432
rect 24051 -11466 24089 -11432
rect 24123 -11466 24161 -11432
rect 24195 -11466 24233 -11432
rect 24267 -11466 24305 -11432
rect 24339 -11466 24377 -11432
rect 24411 -11466 24449 -11432
rect 24483 -11466 24521 -11432
rect 24555 -11466 24593 -11432
rect 24627 -11466 24665 -11432
rect 24699 -11466 24737 -11432
rect 24771 -11466 24809 -11432
rect 24843 -11466 24881 -11432
rect 24915 -11466 24953 -11432
rect 24987 -11466 25025 -11432
rect 25059 -11466 25097 -11432
rect 25131 -11466 25169 -11432
rect 25203 -11466 25241 -11432
rect 25275 -11466 25313 -11432
rect 25347 -11466 25385 -11432
rect 25419 -11466 25457 -11432
rect 25491 -11466 25529 -11432
rect 25563 -11466 25601 -11432
rect 25635 -11466 25673 -11432
rect 25707 -11466 25745 -11432
rect 25779 -11466 25817 -11432
rect 25851 -11466 25889 -11432
rect 25923 -11466 25961 -11432
rect 25995 -11466 26033 -11432
rect 26067 -11466 26105 -11432
rect 26139 -11466 26177 -11432
rect 26211 -11466 26249 -11432
rect 26283 -11466 26295 -11432
rect 23253 -11472 26295 -11466
rect 23137 -11478 23253 -11472
rect 22966 -11558 22972 -11506
rect 23024 -11558 23036 -11506
rect 23088 -11558 23094 -11506
rect 23401 -11569 23407 -11517
rect 23459 -11569 23471 -11517
rect 23523 -11545 28144 -11517
rect 23523 -11569 23529 -11545
rect 23249 -11651 23255 -11599
rect 23307 -11651 23319 -11599
rect 23371 -11622 23377 -11599
rect 23772 -11601 28263 -11573
rect 23772 -11622 23800 -11601
rect 23371 -11650 23800 -11622
rect 23371 -11651 23377 -11650
tri 21264 -11663 21274 -11653 sw
rect 21236 -11687 21274 -11663
tri 21274 -11687 21298 -11663 sw
rect 23829 -11687 24088 -11663
rect 21236 -11691 24088 -11687
tri 21188 -11715 21193 -11710 sw
rect 21236 -11715 23857 -11691
rect 24082 -11715 24088 -11691
rect 24140 -11715 24152 -11663
rect 24204 -11715 24210 -11663
rect 21160 -11720 21193 -11715
tri 21193 -11720 21198 -11715 sw
rect 21160 -11744 21198 -11720
tri 21198 -11744 21222 -11720 sw
rect 23909 -11744 23915 -11720
tri 21112 -11772 21118 -11766 sw
rect 21160 -11772 23915 -11744
rect 23967 -11772 23979 -11720
rect 24031 -11772 24037 -11720
rect 21072 -11800 21118 -11772
tri 21118 -11800 21146 -11772 sw
tri 24112 -11800 24138 -11774 se
rect 24138 -11800 24145 -11774
rect 21072 -11824 24145 -11800
tri 21072 -11839 21087 -11824 ne
rect 21087 -11826 24145 -11824
rect 24197 -11826 24209 -11774
rect 24261 -11826 24267 -11774
rect 21087 -11839 24129 -11826
tri 24129 -11839 24142 -11826 nw
rect 24471 -11831 24667 -11629
rect 26433 -11831 26459 -11629
rect 28008 -11681 28014 -11629
rect 28066 -11681 28091 -11629
rect 28143 -11681 28167 -11629
rect 28219 -11681 28225 -11629
rect 26764 -11721 26792 -11693
rect 28008 -11703 28225 -11681
rect 28008 -11755 28014 -11703
rect 28066 -11755 28091 -11703
rect 28143 -11755 28167 -11703
rect 28219 -11755 28225 -11703
rect 28008 -11777 28225 -11755
rect 28008 -11829 28014 -11777
rect 28066 -11829 28091 -11777
rect 28143 -11829 28167 -11777
rect 28219 -11829 28225 -11777
tri 24145 -11867 24158 -11854 se
rect 24158 -11867 24164 -11854
tri 22784 -11873 22790 -11867 se
rect 22790 -11873 22796 -11867
rect 20992 -11913 22796 -11873
tri 22784 -11919 22790 -11913 ne
rect 22790 -11919 22796 -11913
rect 22848 -11919 22860 -11867
rect 22912 -11873 22918 -11867
tri 22918 -11873 22924 -11867 sw
tri 24139 -11873 24145 -11867 se
rect 24145 -11873 24164 -11867
rect 22912 -11906 24164 -11873
rect 24216 -11906 24228 -11854
rect 24280 -11906 24286 -11854
rect 22912 -11913 22924 -11906
tri 22924 -11913 22931 -11906 nw
rect 22912 -11919 22918 -11913
tri 22918 -11919 22924 -11913 nw
tri 19639 -11947 19663 -11923 se
rect 19663 -11947 19669 -11923
rect 16407 -11953 19669 -11947
rect 16459 -11975 19669 -11953
rect 19721 -11975 19733 -11923
rect 19785 -11934 19791 -11923
tri 19791 -11934 19802 -11923 sw
rect 19785 -11947 19802 -11934
tri 19802 -11947 19815 -11934 sw
rect 24140 -11947 24146 -11934
rect 19785 -11975 24146 -11947
rect 16459 -11986 16482 -11975
tri 16482 -11986 16493 -11975 nw
rect 24140 -11986 24146 -11975
rect 24198 -11986 24210 -11934
rect 24262 -11986 24268 -11934
rect 16459 -11996 16472 -11986
tri 16472 -11996 16482 -11986 nw
rect 16459 -12003 16465 -11996
tri 16465 -12003 16472 -11996 nw
rect 16407 -12017 16459 -12005
tri 16459 -12009 16465 -12003 nw
rect 16919 -12055 16925 -12003
rect 16977 -12055 16989 -12003
rect 17041 -12016 17047 -12003
tri 17047 -12016 17060 -12003 sw
rect 24298 -12016 24304 -11996
rect 17041 -12046 24304 -12016
rect 17041 -12055 17047 -12046
tri 17047 -12055 17056 -12046 nw
rect 24298 -12048 24304 -12046
rect 24356 -12048 24368 -11996
rect 24420 -12048 24426 -11996
tri 24466 -12048 24471 -12043 se
rect 24471 -12048 24601 -11831
tri 24601 -11897 24667 -11831 nw
rect 24696 -11919 24702 -11867
rect 24754 -11919 24766 -11867
rect 24818 -11919 24824 -11867
rect 25603 -11917 25609 -11865
rect 25661 -11917 25673 -11865
rect 25725 -11917 25731 -11865
tri 24459 -12055 24466 -12048 se
rect 24466 -12055 24601 -12048
rect 16407 -12075 16459 -12069
tri 24439 -12075 24459 -12055 se
rect 24459 -12075 24601 -12055
tri 24438 -12076 24439 -12075 se
rect 24439 -12076 24601 -12075
tri 17457 -12126 17481 -12102 nw
tri 16789 -12170 16823 -12136 sw
tri 16696 -12206 16705 -12197 sw
rect 24360 -12206 24601 -12076
rect 26678 -12103 26684 -12051
rect 26736 -12103 26748 -12051
rect 26800 -12103 26806 -12051
rect 24810 -12157 24816 -12105
rect 24868 -12157 24880 -12105
rect 24932 -12157 24938 -12105
rect 16696 -12221 16705 -12206
tri 16705 -12221 16720 -12206 sw
rect 25663 -12221 25669 -12169
rect 25721 -12221 25733 -12169
rect 25785 -12221 25791 -12169
rect 27110 -12221 27116 -12169
rect 27168 -12221 27180 -12169
rect 27232 -12221 27238 -12169
rect 27954 -12190 27960 -12138
rect 28012 -12190 28028 -12138
rect 28080 -12190 28086 -12138
rect 16696 -12225 16720 -12221
tri 16720 -12225 16724 -12221 sw
rect 16696 -12226 16724 -12225
tri 16724 -12226 16725 -12225 sw
rect 24849 -12241 24877 -12232
rect 16691 -12255 16696 -12251
tri 16696 -12255 16700 -12251 nw
tri 16576 -12271 16588 -12259 sw
rect 16576 -12293 16588 -12271
tri 16588 -12293 16610 -12271 sw
tri 23721 -12323 23727 -12317 ne
rect 23727 -12323 23733 -12271
rect 23785 -12323 23797 -12271
rect 23849 -12323 23855 -12271
rect 23993 -12315 24065 -12272
rect 24796 -12293 24802 -12241
rect 24854 -12293 24868 -12241
rect 24920 -12293 24926 -12241
rect 25049 -12293 25055 -12241
rect 25107 -12293 25119 -12241
rect 25171 -12293 25177 -12241
rect 26333 -12299 26559 -12253
rect 26629 -12291 26657 -12263
rect 27730 -12295 27736 -12243
rect 27788 -12295 27800 -12243
rect 27852 -12295 27858 -12243
rect 27966 -12277 27972 -12225
rect 28024 -12277 28036 -12225
rect 28088 -12277 28094 -12225
tri 23855 -12323 23861 -12317 nw
rect 22632 -12352 22684 -12349
rect 17572 -12404 17578 -12352
rect 17630 -12404 17642 -12352
rect 17694 -12370 20823 -12352
rect 21084 -12355 22684 -12352
rect 21084 -12370 22632 -12355
rect 17694 -12382 22632 -12370
rect 17694 -12400 17704 -12382
tri 17704 -12400 17722 -12382 nw
rect 20793 -12400 21114 -12382
rect 17694 -12404 17700 -12400
tri 17700 -12404 17704 -12400 nw
rect 23175 -12352 23227 -12346
tri 17993 -12506 18089 -12410 se
rect 18089 -12462 18429 -12410
rect 18481 -12462 18508 -12410
rect 18560 -12462 18586 -12410
rect 18638 -12462 18664 -12410
rect 18716 -12462 18742 -12410
rect 18794 -12462 18800 -12410
rect 18089 -12506 18800 -12462
rect 22632 -12419 22684 -12407
rect 22734 -12422 22762 -12394
rect 23095 -12422 23123 -12394
tri 24281 -12392 24288 -12385 se
rect 23175 -12419 23227 -12404
rect 22632 -12477 22684 -12471
rect 24288 -12437 24294 -12385
rect 24346 -12437 24358 -12385
rect 24410 -12437 24416 -12385
tri 24674 -12425 24693 -12406 se
tri 24662 -12437 24674 -12425 se
rect 24674 -12437 24693 -12425
rect 23175 -12477 23227 -12471
tri 24622 -12477 24662 -12437 se
rect 24662 -12477 24693 -12437
tri 24614 -12485 24622 -12477 se
rect 24622 -12485 24693 -12477
tri 24760 -12452 24787 -12425 sw
rect 24760 -12477 24787 -12452
tri 24787 -12477 24812 -12452 sw
rect 24760 -12485 24812 -12477
tri 24812 -12485 24820 -12477 sw
tri 24593 -12506 24614 -12485 se
rect 24614 -12506 24693 -12485
tri 17950 -12549 17993 -12506 se
rect 17993 -12516 18800 -12506
rect 17993 -12549 18429 -12516
rect 18009 -12568 18429 -12549
rect 18481 -12568 18508 -12516
rect 18560 -12568 18586 -12516
rect 18638 -12568 18664 -12516
rect 18716 -12568 18742 -12516
rect 18794 -12568 18800 -12516
rect 18009 -12569 18800 -12568
rect 23066 -12558 23072 -12506
rect 23124 -12558 23166 -12506
rect 23218 -12558 23259 -12506
rect 23311 -12558 23317 -12506
rect 18009 -12636 18090 -12569
tri 18090 -12636 18157 -12569 nw
rect 23066 -12584 23317 -12558
rect 23066 -12636 23072 -12584
rect 23124 -12636 23166 -12584
rect 23218 -12636 23259 -12584
rect 23311 -12636 23317 -12584
rect 24360 -12507 24693 -12506
rect 24360 -12636 24647 -12507
rect 18009 -12649 18077 -12636
tri 18077 -12649 18090 -12636 nw
tri 24617 -12649 24630 -12636 ne
rect 24630 -12649 24647 -12636
rect 17217 -12677 17245 -12649
rect 18009 -12677 18049 -12649
tri 18049 -12677 18077 -12649 nw
tri 24630 -12666 24647 -12649 ne
rect 26438 -12666 26454 -12452
rect 28182 -12531 28210 -12503
tri 18009 -12717 18049 -12677 nw
tri 17408 -12785 17414 -12779 se
rect 17414 -12831 17420 -12779
rect 17472 -12831 17484 -12779
rect 17536 -12831 17639 -12779
rect 17562 -12978 17614 -12972
rect 16960 -13013 17012 -13007
rect 16382 -13106 16388 -13054
rect 16440 -13106 16452 -13054
rect 16504 -13106 16514 -13054
tri 17524 -13055 17562 -13017 ne
rect 17562 -13042 17614 -13030
tri 16942 -13089 16960 -13071 se
rect 16960 -13077 17012 -13065
tri 16775 -13135 16788 -13122 ne
rect 16788 -13135 16809 -13122
tri 17012 -13090 17041 -13061 sw
tri 17614 -13051 17648 -13017 nw
rect 17562 -13100 17614 -13094
rect 17899 -13097 17951 -13091
rect 16960 -13135 17012 -13129
tri 16788 -13142 16795 -13135 ne
rect 16795 -13142 16809 -13135
rect 16372 -13194 16380 -13142
rect 16432 -13194 16444 -13142
rect 16496 -13194 16502 -13142
tri 16795 -13156 16809 -13142 ne
tri 17882 -13156 17899 -13139 se
rect 17899 -13156 17951 -13149
tri 17876 -13162 17882 -13156 se
rect 17882 -13161 17951 -13156
rect 17882 -13162 17899 -13161
rect 16605 -13214 16613 -13162
rect 16665 -13214 16677 -13162
rect 16729 -13214 16735 -13162
tri 17865 -13173 17876 -13162 se
rect 17876 -13173 17899 -13162
rect 17759 -13207 17787 -13179
rect 17899 -13219 17951 -13213
tri 16634 -13286 16668 -13252 sw
tri 16223 -13372 16267 -13328 se
rect 16634 -13346 16654 -13332
tri 16654 -13346 16668 -13332 nw
tri 16338 -13372 16364 -13346 sw
tri 16634 -13366 16654 -13346 nw
rect 16338 -13405 16364 -13372
tri 16364 -13405 16397 -13372 sw
tri 16482 -13405 16502 -13385 se
tri 16548 -13405 16568 -13385 sw
rect 17060 -13513 17088 -13485
<< via1 >>
rect 17004 -6668 17056 -6616
rect 16250 -6698 16302 -6686
rect 16250 -6732 16271 -6698
rect 16271 -6732 16302 -6698
rect 16250 -6738 16302 -6732
rect 16314 -6738 16366 -6686
rect 17004 -6732 17056 -6680
rect 20221 -7018 20273 -6966
rect 18469 -7089 18521 -7037
rect 18533 -7089 18585 -7037
rect 20221 -7082 20273 -7030
rect 18581 -7261 18633 -7209
rect 18645 -7261 18697 -7209
rect 20071 -7261 20123 -7209
rect 20135 -7261 20187 -7209
rect 18343 -7344 18395 -7292
rect 18343 -7408 18395 -7356
rect 18543 -7368 18595 -7316
rect 18543 -7432 18595 -7380
rect 20410 -7359 20462 -7307
rect 20474 -7359 20526 -7307
rect 20057 -7454 20109 -7402
rect 20121 -7454 20173 -7402
rect 21068 -7362 21120 -7310
rect 20988 -7461 21040 -7409
rect 21068 -7426 21120 -7374
rect 20988 -7525 21040 -7473
rect 17583 -7718 17635 -7666
rect 17647 -7718 17699 -7666
rect 18909 -7718 18961 -7666
rect 18973 -7718 19025 -7666
rect 20593 -7773 20645 -7721
rect 20657 -7773 20709 -7721
rect 16678 -7857 16730 -7805
rect 16678 -7921 16730 -7869
rect 16778 -7860 16830 -7808
rect 16778 -7924 16830 -7872
rect 19725 -7885 19777 -7833
rect 19789 -7885 19841 -7833
rect 20593 -7854 20645 -7802
rect 20657 -7854 20709 -7802
rect 16453 -8043 16505 -7991
rect 16453 -8107 16505 -8055
rect 16922 -7974 16974 -7922
rect 17008 -7974 17060 -7922
rect 16922 -8039 16974 -7987
rect 17008 -8039 17060 -7987
rect 16922 -8104 16974 -8052
rect 17008 -8104 17060 -8052
rect 17874 -7970 17926 -7918
rect 17944 -7970 17996 -7918
rect 18013 -7970 18065 -7918
rect 17874 -8040 17926 -7988
rect 17944 -8040 17996 -7988
rect 18013 -8040 18065 -7988
rect 17874 -8110 17926 -8058
rect 17944 -8110 17996 -8058
rect 18013 -8110 18065 -8058
rect 18129 -8199 18181 -8147
rect 18203 -8199 18255 -8147
rect 18277 -8199 18329 -8147
rect 18129 -8268 18181 -8216
rect 18203 -8268 18255 -8216
rect 18277 -8268 18329 -8216
rect 18129 -8337 18181 -8285
rect 18203 -8337 18255 -8285
rect 18277 -8337 18329 -8285
rect 20000 -8194 20052 -8142
rect 20086 -8194 20138 -8142
rect 20171 -8194 20223 -8142
rect 20256 -8194 20308 -8142
rect 20000 -8268 20052 -8216
rect 20086 -8268 20138 -8216
rect 20171 -8268 20223 -8216
rect 20256 -8268 20308 -8216
rect 20000 -8342 20052 -8290
rect 20086 -8342 20138 -8290
rect 20171 -8342 20223 -8290
rect 20256 -8342 20308 -8290
rect 17697 -8435 17749 -8383
rect 17697 -8499 17749 -8447
rect 18682 -8435 18734 -8383
rect 18682 -8499 18734 -8447
rect 16521 -8696 16573 -8644
rect 16585 -8696 16637 -8644
rect 17414 -8733 17466 -8681
rect 17478 -8733 17530 -8681
rect 16526 -8786 16578 -8734
rect 16590 -8786 16642 -8734
rect 17779 -8741 17831 -8689
rect 18916 -8727 18968 -8675
rect 18981 -8727 19033 -8675
rect 19769 -8696 19821 -8644
rect 19833 -8696 19885 -8644
rect 16757 -8803 16809 -8751
rect 16821 -8803 16873 -8751
rect 17779 -8805 17831 -8753
rect 16909 -9055 16961 -9003
rect 17009 -9055 17061 -9003
rect 16909 -9135 16961 -9083
rect 17009 -9135 17061 -9083
rect 16909 -9216 16961 -9164
rect 17009 -9216 17061 -9164
rect 16909 -9297 16961 -9245
rect 17009 -9297 17061 -9245
rect 17870 -9055 17922 -9003
rect 17944 -9055 17996 -9003
rect 18018 -9055 18070 -9003
rect 17870 -9135 17922 -9083
rect 17944 -9135 17996 -9083
rect 18018 -9135 18070 -9083
rect 17870 -9216 17922 -9164
rect 17944 -9216 17996 -9164
rect 18018 -9216 18070 -9164
rect 17870 -9297 17922 -9245
rect 17944 -9297 17996 -9245
rect 18018 -9297 18070 -9245
rect 16526 -9565 16578 -9513
rect 16590 -9565 16642 -9513
rect 16757 -9548 16809 -9496
rect 16821 -9548 16873 -9496
rect 17779 -9547 17831 -9495
rect 16521 -9656 16573 -9604
rect 16585 -9656 16637 -9604
rect 17415 -9622 17467 -9570
rect 17479 -9622 17531 -9570
rect 17779 -9611 17831 -9559
rect 18602 -9278 18654 -9226
rect 18602 -9342 18654 -9290
rect 18763 -9377 18815 -9371
rect 18763 -9411 18769 -9377
rect 18769 -9411 18803 -9377
rect 18803 -9411 18815 -9377
rect 18763 -9423 18815 -9411
rect 18763 -9449 18815 -9435
rect 18763 -9483 18769 -9449
rect 18769 -9483 18803 -9449
rect 18803 -9483 18815 -9449
rect 18763 -9487 18815 -9483
rect 19109 -9305 19161 -9299
rect 19109 -9339 19115 -9305
rect 19115 -9339 19161 -9305
rect 19109 -9351 19161 -9339
rect 19109 -9377 19161 -9368
rect 19109 -9411 19115 -9377
rect 19115 -9411 19161 -9377
rect 19109 -9420 19161 -9411
rect 19109 -9449 19161 -9437
rect 19109 -9483 19115 -9449
rect 19115 -9483 19161 -9449
rect 19109 -9489 19161 -9483
rect 19454 -9407 19506 -9399
rect 19454 -9441 19475 -9407
rect 19475 -9441 19506 -9407
rect 19454 -9451 19506 -9441
rect 19454 -9479 19506 -9463
rect 19454 -9513 19475 -9479
rect 19475 -9513 19506 -9479
rect 19454 -9515 19506 -9513
rect 19752 -9227 19804 -9216
rect 19752 -9261 19781 -9227
rect 19781 -9261 19804 -9227
rect 19752 -9268 19804 -9261
rect 19816 -9227 19868 -9216
rect 19816 -9261 19819 -9227
rect 19819 -9261 19853 -9227
rect 19853 -9261 19868 -9227
rect 19816 -9268 19868 -9261
rect 19775 -9407 19827 -9399
rect 19775 -9441 19787 -9407
rect 19787 -9441 19821 -9407
rect 19821 -9441 19827 -9407
rect 20045 -9324 20097 -9314
rect 20045 -9358 20054 -9324
rect 20054 -9358 20088 -9324
rect 20088 -9358 20097 -9324
rect 20045 -9366 20097 -9358
rect 20045 -9396 20097 -9384
rect 19775 -9451 19827 -9441
rect 20045 -9430 20054 -9396
rect 20054 -9430 20088 -9396
rect 20088 -9430 20097 -9396
rect 20045 -9436 20097 -9430
rect 19775 -9479 19827 -9467
rect 19775 -9513 19787 -9479
rect 19787 -9513 19821 -9479
rect 19821 -9513 19827 -9479
rect 19775 -9519 19827 -9513
rect 19556 -9656 19608 -9604
rect 19626 -9656 19678 -9604
rect 19556 -9722 19608 -9670
rect 19626 -9722 19678 -9670
rect 20322 -9677 20374 -9671
rect 20322 -9711 20330 -9677
rect 20330 -9711 20364 -9677
rect 20364 -9711 20374 -9677
rect 20322 -9723 20374 -9711
rect 20322 -9749 20374 -9735
rect 18763 -9818 18815 -9766
rect 18763 -9882 18815 -9830
rect 19109 -9816 19161 -9764
rect 19109 -9880 19161 -9828
rect 19355 -9817 19407 -9765
rect 19355 -9881 19407 -9829
rect 19454 -9818 19506 -9766
rect 19454 -9882 19506 -9830
rect 19775 -9816 19827 -9764
rect 20322 -9783 20330 -9749
rect 20330 -9783 20364 -9749
rect 20364 -9783 20374 -9749
rect 20322 -9787 20374 -9783
rect 19775 -9880 19827 -9828
rect 16585 -10050 16637 -9998
rect 16585 -10114 16637 -10062
rect 18133 -10080 18185 -10028
rect 18198 -10080 18250 -10028
rect 18262 -10080 18314 -10028
rect 18133 -10158 18185 -10106
rect 18198 -10158 18250 -10106
rect 18262 -10158 18314 -10106
rect 20000 -10080 20052 -10028
rect 20086 -10080 20138 -10028
rect 20171 -10080 20223 -10028
rect 20256 -10040 20308 -10028
rect 20256 -10074 20284 -10040
rect 20284 -10074 20308 -10040
rect 20256 -10080 20308 -10074
rect 20000 -10158 20052 -10106
rect 20086 -10158 20138 -10106
rect 20171 -10158 20223 -10106
rect 20256 -10112 20308 -10106
rect 20256 -10146 20284 -10112
rect 20284 -10146 20308 -10112
rect 20256 -10158 20308 -10146
rect 16936 -10245 16988 -10193
rect 17010 -10243 17062 -10193
rect 17010 -10245 17033 -10243
rect 17033 -10245 17062 -10243
rect 16817 -10325 16869 -10273
rect 16817 -10391 16869 -10339
rect 17874 -10260 17926 -10208
rect 17942 -10260 17994 -10208
rect 18009 -10260 18061 -10208
rect 19896 -10247 19948 -10195
rect 19960 -10247 20012 -10195
rect 16936 -10330 16988 -10278
rect 17010 -10330 17062 -10278
rect 16936 -10371 16988 -10364
rect 17010 -10371 17062 -10364
rect 16936 -10405 16979 -10371
rect 16979 -10405 16988 -10371
rect 17010 -10405 17013 -10371
rect 17013 -10405 17062 -10371
rect 16936 -10416 16988 -10405
rect 17010 -10416 17062 -10405
rect 16936 -10477 16979 -10450
rect 16979 -10477 16988 -10450
rect 17010 -10477 17013 -10450
rect 17013 -10477 17062 -10450
rect 16936 -10502 16988 -10477
rect 17010 -10502 17062 -10477
rect 16585 -10575 16637 -10569
rect 18133 -10464 18185 -10412
rect 18203 -10464 18255 -10412
rect 18272 -10464 18324 -10412
rect 20000 -10464 20052 -10412
rect 20086 -10464 20138 -10412
rect 20171 -10464 20223 -10412
rect 20256 -10464 20308 -10412
rect 18133 -10538 18185 -10486
rect 18203 -10538 18255 -10486
rect 18272 -10538 18324 -10486
rect 20000 -10542 20052 -10490
rect 20086 -10542 20138 -10490
rect 20171 -10542 20223 -10490
rect 20256 -10542 20308 -10490
rect 16585 -10609 16635 -10575
rect 16635 -10609 16637 -10575
rect 18644 -10578 18696 -10572
rect 18708 -10578 18760 -10572
rect 16585 -10621 16637 -10609
rect 18644 -10612 18661 -10578
rect 18661 -10612 18696 -10578
rect 18708 -10612 18739 -10578
rect 18739 -10612 18760 -10578
rect 18644 -10624 18696 -10612
rect 18708 -10624 18760 -10612
rect 16585 -10647 16637 -10635
rect 19556 -10629 19608 -10577
rect 19626 -10629 19678 -10577
rect 16585 -10681 16635 -10647
rect 16635 -10681 16637 -10647
rect 16585 -10687 16637 -10681
rect 18133 -10733 18185 -10681
rect 18200 -10733 18252 -10681
rect 19556 -10695 19608 -10643
rect 19626 -10695 19678 -10643
rect 18133 -10797 18185 -10745
rect 18200 -10797 18252 -10745
rect 20102 -11341 20154 -11332
rect 20180 -11341 20232 -11332
rect 20257 -11341 20309 -11332
rect 20102 -11375 20130 -11341
rect 20130 -11375 20154 -11341
rect 20180 -11375 20203 -11341
rect 20203 -11375 20232 -11341
rect 20257 -11375 20276 -11341
rect 20276 -11375 20309 -11341
rect 20102 -11384 20154 -11375
rect 20180 -11384 20232 -11375
rect 20257 -11384 20309 -11375
rect 17691 -11461 17743 -11409
rect 17755 -11461 17807 -11409
rect 19349 -11461 19401 -11409
rect 19413 -11461 19465 -11409
rect 16869 -11605 16921 -11553
rect 16933 -11605 16985 -11553
rect 19775 -11611 19827 -11559
rect 19775 -11675 19827 -11623
rect 17473 -11747 17525 -11695
rect 18374 -11728 18426 -11676
rect 18438 -11728 18490 -11676
rect 17473 -11811 17525 -11759
rect 17578 -11814 17630 -11762
rect 17642 -11814 17694 -11762
rect 18490 -11808 18542 -11756
rect 18554 -11808 18606 -11756
rect 21236 -7762 21288 -7710
rect 21147 -7860 21199 -7808
rect 21147 -7924 21199 -7872
rect 21236 -7826 21288 -7774
rect 22761 -8667 22813 -8615
rect 22825 -8667 22877 -8615
rect 23071 -8979 23123 -8927
rect 23156 -8979 23208 -8927
rect 23241 -8979 23293 -8927
rect 23402 -9925 23454 -9873
rect 23402 -9991 23454 -9939
rect 23234 -10198 23286 -10146
rect 23298 -10198 23350 -10146
rect 23060 -10311 23112 -10259
rect 23178 -10311 23230 -10259
rect 23137 -11321 23189 -11269
rect 23201 -11321 23253 -11269
rect 23137 -11396 23189 -11344
rect 23201 -11396 23253 -11344
rect 23137 -11432 23189 -11420
rect 23137 -11466 23151 -11432
rect 23151 -11466 23185 -11432
rect 23185 -11466 23189 -11432
rect 23137 -11472 23189 -11466
rect 23201 -11432 23253 -11420
rect 23201 -11466 23224 -11432
rect 23224 -11466 23253 -11432
rect 23201 -11472 23253 -11466
rect 22972 -11558 23024 -11506
rect 23036 -11558 23088 -11506
rect 23407 -11569 23459 -11517
rect 23471 -11569 23523 -11517
rect 23255 -11651 23307 -11599
rect 23319 -11651 23371 -11599
rect 24088 -11715 24140 -11663
rect 24152 -11715 24204 -11663
rect 23915 -11772 23967 -11720
rect 23979 -11772 24031 -11720
rect 24145 -11826 24197 -11774
rect 24209 -11826 24261 -11774
rect 28014 -11681 28066 -11629
rect 28091 -11681 28143 -11629
rect 28167 -11681 28219 -11629
rect 28014 -11755 28066 -11703
rect 28091 -11755 28143 -11703
rect 28167 -11755 28219 -11703
rect 28014 -11829 28066 -11777
rect 28091 -11829 28143 -11777
rect 28167 -11829 28219 -11777
rect 22796 -11919 22848 -11867
rect 22860 -11919 22912 -11867
rect 24164 -11906 24216 -11854
rect 24228 -11906 24280 -11854
rect 16407 -12005 16459 -11953
rect 19669 -11975 19721 -11923
rect 19733 -11975 19785 -11923
rect 24146 -11986 24198 -11934
rect 24210 -11986 24262 -11934
rect 16407 -12069 16459 -12017
rect 16925 -12055 16977 -12003
rect 16989 -12055 17041 -12003
rect 24304 -12048 24356 -11996
rect 24368 -12048 24420 -11996
rect 24702 -11919 24754 -11867
rect 24766 -11919 24818 -11867
rect 25609 -11917 25661 -11865
rect 25673 -11917 25725 -11865
rect 26684 -12103 26736 -12051
rect 26748 -12103 26800 -12051
rect 24816 -12157 24868 -12105
rect 24880 -12157 24932 -12105
rect 25669 -12221 25721 -12169
rect 25733 -12221 25785 -12169
rect 27116 -12221 27168 -12169
rect 27180 -12221 27232 -12169
rect 27960 -12190 28012 -12138
rect 28028 -12190 28080 -12138
rect 23733 -12323 23785 -12271
rect 23797 -12323 23849 -12271
rect 24802 -12293 24854 -12241
rect 24868 -12293 24920 -12241
rect 25055 -12293 25107 -12241
rect 25119 -12293 25171 -12241
rect 27736 -12295 27788 -12243
rect 27800 -12295 27852 -12243
rect 27972 -12277 28024 -12225
rect 28036 -12277 28088 -12225
rect 17578 -12404 17630 -12352
rect 17642 -12404 17694 -12352
rect 22632 -12407 22684 -12355
rect 18429 -12462 18481 -12410
rect 18508 -12462 18560 -12410
rect 18586 -12462 18638 -12410
rect 18664 -12462 18716 -12410
rect 18742 -12462 18794 -12410
rect 22632 -12471 22684 -12419
rect 23175 -12404 23227 -12352
rect 23175 -12471 23227 -12419
rect 24294 -12437 24346 -12385
rect 24358 -12437 24410 -12385
rect 18429 -12568 18481 -12516
rect 18508 -12568 18560 -12516
rect 18586 -12568 18638 -12516
rect 18664 -12568 18716 -12516
rect 18742 -12568 18794 -12516
rect 23072 -12558 23124 -12506
rect 23166 -12558 23218 -12506
rect 23259 -12558 23311 -12506
rect 23072 -12636 23124 -12584
rect 23166 -12636 23218 -12584
rect 23259 -12636 23311 -12584
rect 17420 -12831 17472 -12779
rect 17484 -12831 17536 -12779
rect 16388 -13106 16440 -13054
rect 16452 -13106 16504 -13054
rect 16960 -13065 17012 -13013
rect 17562 -13030 17614 -12978
rect 16960 -13129 17012 -13077
rect 17562 -13094 17614 -13042
rect 16380 -13194 16432 -13142
rect 16444 -13194 16496 -13142
rect 17899 -13149 17951 -13097
rect 16613 -13214 16665 -13162
rect 16677 -13214 16729 -13162
rect 17899 -13213 17951 -13161
<< metal2 >>
rect 17004 -6616 17056 -6610
tri 16988 -6668 17004 -6652 se
tri 16976 -6680 16988 -6668 se
rect 16988 -6680 17056 -6668
tri 16970 -6686 16976 -6680 se
rect 16976 -6686 17004 -6680
rect 16244 -6738 16250 -6686
rect 16302 -6738 16314 -6686
rect 16366 -6732 17004 -6686
rect 16366 -6738 17056 -6732
rect 18462 -6966 20273 -6960
rect 18462 -7018 20221 -6966
rect 18462 -7030 20273 -7018
rect 18462 -7037 20221 -7030
rect 18462 -7089 18469 -7037
rect 18521 -7089 18533 -7037
rect 18585 -7082 20221 -7037
rect 18585 -7088 20273 -7082
rect 18585 -7089 20265 -7088
rect 18575 -7261 18581 -7209
rect 18633 -7261 18645 -7209
rect 18697 -7261 20071 -7209
rect 20123 -7261 20135 -7209
rect 20187 -7261 20193 -7209
rect 18343 -7292 18395 -7286
rect 18343 -7356 18395 -7344
rect 18343 -7414 18395 -7408
rect 18543 -7316 18595 -7310
rect 18543 -7380 18595 -7368
rect 18357 -7473 18385 -7414
rect 18543 -7438 18595 -7432
tri 18385 -7473 18386 -7472 sw
rect 18357 -7479 18386 -7473
tri 18386 -7479 18392 -7473 sw
rect 18357 -7496 18392 -7479
tri 18357 -7525 18386 -7496 ne
rect 18386 -7525 18392 -7496
tri 18392 -7525 18438 -7479 sw
tri 18386 -7531 18392 -7525 ne
rect 18392 -7531 18438 -7525
tri 18438 -7531 18444 -7525 sw
tri 18392 -7583 18444 -7531 ne
tri 18444 -7583 18496 -7531 sw
tri 18444 -7607 18468 -7583 ne
rect 17577 -7718 17583 -7666
rect 17635 -7718 17647 -7666
rect 17699 -7718 17705 -7666
rect 17577 -7721 17702 -7718
tri 17702 -7721 17705 -7718 nw
rect 17577 -7773 17650 -7721
tri 17650 -7773 17702 -7721 nw
rect 17577 -7774 17649 -7773
tri 17649 -7774 17650 -7773 nw
rect 16678 -7805 16730 -7799
rect 17577 -7802 17621 -7774
tri 17621 -7802 17649 -7774 nw
rect 16678 -7869 16730 -7857
rect 16678 -7927 16730 -7921
rect 16777 -7808 16830 -7802
rect 16777 -7860 16778 -7808
rect 16777 -7872 16830 -7860
rect 16777 -7924 16778 -7872
rect 16453 -7991 16505 -7985
rect 16453 -8055 16505 -8043
rect 16453 -8113 16505 -8107
rect 16453 -8644 16481 -8113
rect 16453 -8696 16521 -8644
rect 16573 -8696 16585 -8644
rect 16637 -8696 16643 -8644
tri 16696 -8696 16697 -8695 se
rect 16697 -8696 16725 -7927
rect 16453 -9604 16481 -8696
tri 16659 -8733 16696 -8696 se
rect 16696 -8725 16725 -8696
rect 16696 -8733 16717 -8725
tri 16717 -8733 16725 -8725 nw
rect 16777 -7930 16830 -7924
rect 16909 -7922 17062 -7905
tri 16658 -8734 16659 -8733 se
rect 16659 -8734 16716 -8733
tri 16716 -8734 16717 -8733 nw
rect 16520 -8786 16526 -8734
rect 16578 -8786 16590 -8734
rect 16642 -8741 16709 -8734
tri 16709 -8741 16716 -8734 nw
rect 16642 -8751 16699 -8741
tri 16699 -8751 16709 -8741 nw
rect 16777 -8751 16805 -7930
rect 16909 -7974 16922 -7922
rect 16974 -7974 17008 -7922
rect 17060 -7974 17062 -7922
tri 17525 -7970 17577 -7918 se
rect 17577 -7934 17615 -7802
tri 17615 -7808 17621 -7802 nw
rect 17577 -7970 17579 -7934
tri 17579 -7970 17615 -7934 nw
rect 17868 -7918 18071 -7913
rect 17868 -7925 17874 -7918
tri 17523 -7972 17525 -7970 se
rect 17525 -7972 17577 -7970
tri 17577 -7972 17579 -7970 nw
rect 16909 -7987 17062 -7974
rect 16909 -8039 16922 -7987
rect 16974 -8039 17008 -7987
rect 17060 -8039 17062 -7987
tri 17507 -7988 17523 -7972 se
rect 17523 -7988 17561 -7972
tri 17561 -7988 17577 -7972 nw
rect 17868 -7981 17870 -7925
rect 17926 -7970 17944 -7918
rect 17996 -7925 18013 -7918
rect 17996 -7970 18008 -7925
rect 18065 -7970 18071 -7918
rect 17926 -7981 18008 -7970
rect 18064 -7981 18071 -7970
rect 17868 -7988 18071 -7981
rect 16909 -8052 17062 -8039
rect 16909 -8104 16922 -8052
rect 16974 -8104 17008 -8052
rect 17060 -8104 17062 -8052
rect 16642 -8786 16664 -8751
tri 16664 -8786 16699 -8751 nw
rect 16751 -8803 16757 -8751
rect 16809 -8803 16821 -8751
rect 16873 -8803 16879 -8751
rect 16909 -9003 17062 -8104
tri 17498 -7997 17507 -7988 se
rect 17507 -7997 17552 -7988
tri 17552 -7997 17561 -7988 nw
rect 17498 -8681 17536 -7997
tri 17536 -8013 17552 -7997 nw
rect 17868 -8010 17874 -7988
rect 17868 -8066 17870 -8010
rect 17926 -8040 17944 -7988
rect 17996 -8010 18013 -7988
rect 17996 -8040 18008 -8010
rect 18065 -8040 18071 -7988
rect 17926 -8058 18008 -8040
rect 18064 -8058 18071 -8040
rect 17868 -8095 17874 -8066
rect 17868 -8151 17870 -8095
rect 17926 -8110 17944 -8058
rect 17996 -8066 18008 -8058
rect 17996 -8095 18013 -8066
rect 17996 -8110 18008 -8095
rect 18065 -8110 18071 -8058
rect 17926 -8151 18008 -8110
rect 18064 -8151 18071 -8110
rect 17868 -8180 18071 -8151
rect 17868 -8236 17870 -8180
rect 17926 -8236 18008 -8180
rect 18064 -8236 18071 -8180
rect 17868 -8265 18071 -8236
rect 17868 -8321 17870 -8265
rect 17926 -8321 18008 -8265
rect 18064 -8321 18071 -8265
rect 17868 -8350 18071 -8321
rect 17408 -8733 17414 -8681
rect 17466 -8733 17478 -8681
rect 17530 -8733 17536 -8681
rect 17697 -8383 17749 -8377
rect 17697 -8447 17749 -8435
rect 16961 -9055 17009 -9003
rect 17061 -9055 17062 -9003
rect 16909 -9083 17062 -9055
rect 16961 -9135 17009 -9083
rect 17061 -9135 17062 -9083
rect 16909 -9164 17062 -9135
rect 16961 -9216 17009 -9164
rect 17061 -9216 17062 -9164
rect 16909 -9245 17062 -9216
rect 16961 -9297 17009 -9245
rect 17061 -9297 17062 -9245
rect 16520 -9565 16526 -9513
rect 16578 -9565 16590 -9513
rect 16642 -9548 16673 -9513
tri 16673 -9548 16708 -9513 sw
rect 16747 -9548 16757 -9496
rect 16809 -9548 16821 -9496
rect 16873 -9548 16879 -9496
rect 16642 -9557 16708 -9548
tri 16708 -9557 16717 -9548 sw
rect 16642 -9565 16717 -9557
tri 16659 -9570 16664 -9565 ne
rect 16664 -9570 16717 -9565
tri 16664 -9595 16689 -9570 ne
rect 16453 -9656 16521 -9604
rect 16573 -9656 16585 -9604
rect 16637 -9656 16643 -9604
tri 16684 -9735 16689 -9730 se
rect 16689 -9735 16717 -9570
tri 16668 -9751 16684 -9735 se
rect 16684 -9751 16717 -9735
rect 16668 -9764 16717 -9751
rect 16668 -9766 16715 -9764
tri 16715 -9766 16717 -9764 nw
rect 16747 -9559 16798 -9548
tri 16798 -9559 16809 -9548 nw
rect 16747 -9570 16787 -9559
tri 16787 -9570 16798 -9559 nw
rect 16585 -9998 16637 -9992
rect 16585 -10062 16637 -10050
rect 16585 -10569 16637 -10114
rect 16585 -10635 16637 -10621
rect 16585 -10693 16637 -10687
tri 16539 -11002 16573 -10968 ne
tri 16539 -11154 16573 -11120 se
tri 16610 -11154 16640 -11124 sw
tri 16478 -11164 16484 -11158 nw
tri 16539 -11240 16573 -11206 ne
tri 16610 -11236 16640 -11206 nw
tri 16549 -11553 16573 -11529 se
tri 16539 -11563 16549 -11553 se
rect 16549 -11563 16573 -11553
tri 16613 -11553 16625 -11541 sw
rect 16613 -11563 16625 -11553
tri 16625 -11563 16635 -11553 sw
tri 16473 -11654 16484 -11643 sw
tri 16340 -11711 16352 -11699 se
tri 16276 -11747 16279 -11744 sw
rect 16276 -11756 16279 -11747
tri 16279 -11756 16288 -11747 sw
rect 16276 -11759 16288 -11756
tri 16288 -11759 16291 -11756 sw
rect 16276 -11768 16291 -11759
tri 16291 -11768 16300 -11759 sw
rect 16407 -11953 16459 -11947
rect 16407 -12017 16459 -12005
rect 16407 -12075 16459 -12069
tri 16407 -12099 16431 -12075 ne
rect 16431 -13054 16459 -12075
tri 16666 -12105 16668 -12103 se
rect 16668 -12105 16696 -9766
tri 16696 -9785 16715 -9766 nw
tri 16644 -12127 16666 -12105 se
rect 16666 -12127 16696 -12105
rect 16668 -12255 16696 -12127
tri 16644 -12271 16660 -12255 ne
rect 16660 -12271 16696 -12255
tri 16660 -12279 16668 -12271 ne
tri 16658 -13013 16668 -13003 se
rect 16668 -13013 16696 -12271
tri 16625 -13046 16658 -13013 se
rect 16658 -13018 16696 -13013
rect 16658 -13046 16668 -13018
tri 16668 -13046 16696 -13018 nw
tri 16617 -13054 16625 -13046 se
rect 16625 -13054 16649 -13046
rect 16382 -13106 16388 -13054
rect 16440 -13106 16452 -13054
rect 16504 -13106 16510 -13054
tri 16606 -13065 16617 -13054 se
rect 16617 -13065 16649 -13054
tri 16649 -13065 16668 -13046 nw
tri 16594 -13077 16606 -13065 se
rect 16606 -13077 16637 -13065
tri 16637 -13077 16649 -13065 nw
tri 16582 -13089 16594 -13077 se
rect 16594 -13089 16625 -13077
tri 16625 -13089 16637 -13077 nw
tri 16565 -13106 16582 -13089 se
rect 16582 -13106 16585 -13089
tri 16542 -13129 16565 -13106 se
rect 16565 -13129 16585 -13106
tri 16585 -13129 16625 -13089 nw
tri 16539 -13132 16542 -13129 se
rect 16542 -13132 16582 -13129
tri 16582 -13132 16585 -13129 nw
tri 16537 -13134 16539 -13132 se
rect 16539 -13134 16580 -13132
tri 16580 -13134 16582 -13132 nw
tri 16529 -13142 16537 -13134 se
rect 16537 -13142 16572 -13134
tri 16572 -13142 16580 -13134 nw
tri 16739 -13142 16747 -13134 se
rect 16747 -13142 16775 -9570
tri 16775 -9582 16787 -9570 nw
rect 16909 -10193 17062 -9297
rect 17440 -9570 17492 -8733
rect 17409 -9622 17415 -9570
rect 17467 -9622 17479 -9570
rect 17531 -9622 17537 -9570
rect 16909 -10245 16936 -10193
rect 16988 -10245 17010 -10193
rect 16817 -10273 16869 -10267
rect 16817 -10339 16869 -10325
rect 16817 -11605 16869 -10391
rect 16909 -10278 17062 -10245
rect 16909 -10330 16936 -10278
rect 16988 -10330 17010 -10278
rect 16909 -10364 17062 -10330
rect 16909 -10416 16936 -10364
rect 16988 -10416 17010 -10364
rect 16909 -10450 17062 -10416
rect 16909 -10502 16936 -10450
rect 16988 -10502 17010 -10450
rect 16909 -10508 17062 -10502
rect 17697 -11409 17749 -8499
rect 17868 -8406 17870 -8350
rect 17926 -8406 18008 -8350
rect 18064 -8406 18071 -8350
rect 17868 -8435 18071 -8406
rect 17868 -8491 17870 -8435
rect 17926 -8491 18008 -8435
rect 18064 -8491 18071 -8435
rect 17868 -8520 18071 -8491
rect 17868 -8576 17870 -8520
rect 17926 -8576 18008 -8520
rect 18064 -8576 18071 -8520
rect 17868 -8606 18071 -8576
rect 17868 -8662 17870 -8606
rect 17926 -8662 18008 -8606
rect 18064 -8662 18071 -8606
rect 17779 -8689 17831 -8683
rect 17779 -8753 17831 -8741
rect 17779 -9495 17831 -8805
rect 17779 -9559 17831 -9547
rect 17779 -10890 17831 -9611
rect 17868 -9003 18071 -8662
rect 17868 -9055 17870 -9003
rect 17922 -9055 17944 -9003
rect 17996 -9055 18018 -9003
rect 18070 -9055 18071 -9003
rect 17868 -9083 18071 -9055
rect 17868 -9135 17870 -9083
rect 17922 -9087 17944 -9083
rect 17996 -9087 18018 -9083
rect 17927 -9135 17944 -9087
rect 18070 -9135 18071 -9083
rect 17868 -9143 17871 -9135
rect 17927 -9143 17977 -9135
rect 18033 -9143 18071 -9135
rect 17868 -9164 18071 -9143
rect 17868 -9216 17870 -9164
rect 17922 -9169 17944 -9164
rect 17996 -9169 18018 -9164
rect 17927 -9216 17944 -9169
rect 18070 -9216 18071 -9164
rect 17868 -9225 17871 -9216
rect 17927 -9225 17977 -9216
rect 18033 -9225 18071 -9216
rect 17868 -9245 18071 -9225
rect 17868 -9297 17870 -9245
rect 17922 -9251 17944 -9245
rect 17996 -9251 18018 -9245
rect 17927 -9297 17944 -9251
rect 18070 -9297 18071 -9245
rect 17868 -9307 17871 -9297
rect 17927 -9307 17977 -9297
rect 18033 -9307 18071 -9297
rect 17868 -9333 18071 -9307
rect 17868 -9389 17871 -9333
rect 17927 -9389 17977 -9333
rect 18033 -9389 18071 -9333
rect 17868 -9415 18071 -9389
rect 17868 -9471 17871 -9415
rect 17927 -9471 17977 -9415
rect 18033 -9471 18071 -9415
rect 17868 -9497 18071 -9471
rect 17868 -9553 17871 -9497
rect 17927 -9553 17977 -9497
rect 18033 -9553 18071 -9497
rect 17868 -9579 18071 -9553
rect 17868 -9635 17871 -9579
rect 17927 -9635 17977 -9579
rect 18033 -9635 18071 -9579
rect 17868 -9661 18071 -9635
rect 17868 -9717 17871 -9661
rect 17927 -9717 17977 -9661
rect 18033 -9717 18071 -9661
rect 17868 -9743 18071 -9717
rect 17868 -9799 17871 -9743
rect 17927 -9799 17977 -9743
rect 18033 -9799 18071 -9743
rect 17868 -9825 18071 -9799
rect 17868 -9881 17871 -9825
rect 17927 -9881 17977 -9825
rect 18033 -9881 18071 -9825
rect 17868 -9907 18071 -9881
rect 17868 -9963 17871 -9907
rect 17927 -9963 17977 -9907
rect 18033 -9963 18071 -9907
rect 17868 -9989 18071 -9963
rect 17868 -10045 17871 -9989
rect 17927 -10045 17977 -9989
rect 18033 -10045 18071 -9989
rect 17868 -10071 18071 -10045
rect 17868 -10127 17871 -10071
rect 17927 -10127 17977 -10071
rect 18033 -10127 18071 -10071
rect 17868 -10153 18071 -10127
rect 17868 -10209 17871 -10153
rect 17927 -10208 17977 -10153
rect 18033 -10208 18071 -10153
rect 17927 -10209 17942 -10208
rect 17868 -10235 17874 -10209
rect 17926 -10235 17942 -10209
rect 17994 -10235 18009 -10209
rect 17868 -10291 17871 -10235
rect 17927 -10260 17942 -10235
rect 18061 -10260 18071 -10208
rect 17927 -10291 17977 -10260
rect 18033 -10291 18071 -10260
rect 17868 -10318 18071 -10291
rect 17868 -10374 17871 -10318
rect 17927 -10374 17977 -10318
rect 18033 -10374 18071 -10318
rect 17868 -10401 18071 -10374
rect 17868 -10457 17871 -10401
rect 17927 -10457 17977 -10401
rect 18033 -10457 18071 -10401
rect 17868 -10470 18071 -10457
rect 18127 -8147 18330 -8141
rect 18127 -8199 18129 -8147
rect 18181 -8199 18203 -8147
rect 18255 -8199 18277 -8147
rect 18329 -8199 18330 -8147
rect 18127 -8216 18330 -8199
rect 18127 -8268 18129 -8216
rect 18181 -8268 18203 -8216
rect 18255 -8268 18277 -8216
rect 18329 -8268 18330 -8216
rect 18127 -8285 18330 -8268
rect 18127 -8337 18129 -8285
rect 18181 -8337 18203 -8285
rect 18255 -8337 18277 -8285
rect 18329 -8337 18330 -8285
rect 18127 -10028 18330 -8337
rect 18127 -10080 18133 -10028
rect 18185 -10080 18198 -10028
rect 18250 -10080 18262 -10028
rect 18314 -10080 18330 -10028
rect 18127 -10106 18330 -10080
rect 18127 -10158 18133 -10106
rect 18185 -10158 18198 -10106
rect 18250 -10158 18262 -10106
rect 18314 -10158 18330 -10106
rect 18127 -10412 18330 -10158
rect 18127 -10464 18133 -10412
rect 18185 -10464 18203 -10412
rect 18255 -10464 18272 -10412
rect 18324 -10464 18330 -10412
rect 18127 -10486 18330 -10464
rect 18127 -10538 18133 -10486
rect 18185 -10538 18203 -10486
rect 18255 -10538 18272 -10486
rect 18324 -10538 18330 -10486
rect 18127 -10554 18330 -10538
rect 18127 -10572 18312 -10554
tri 18312 -10572 18330 -10554 nw
rect 18127 -10624 18260 -10572
tri 18260 -10624 18312 -10572 nw
rect 18127 -10681 18258 -10624
tri 18258 -10626 18260 -10624 nw
rect 18127 -10733 18133 -10681
rect 18185 -10733 18200 -10681
rect 18252 -10733 18258 -10681
rect 18127 -10745 18258 -10733
rect 18127 -10797 18133 -10745
rect 18185 -10797 18200 -10745
rect 18252 -10797 18258 -10745
tri 17779 -10895 17784 -10890 ne
rect 17784 -10895 17831 -10890
tri 17831 -10895 17858 -10868 sw
tri 17784 -10942 17831 -10895 ne
rect 17831 -10942 17961 -10895
tri 17831 -10947 17836 -10942 ne
rect 17836 -10947 17961 -10942
tri 17939 -10948 17940 -10947 ne
rect 17940 -10948 17961 -10947
tri 17961 -10948 18014 -10895 sw
tri 17940 -10969 17961 -10948 ne
rect 17961 -10969 18014 -10948
tri 17961 -10990 17982 -10969 ne
rect 17685 -11461 17691 -11409
rect 17743 -11461 17755 -11409
rect 17807 -11461 17813 -11409
rect 16921 -11605 16933 -11553
rect 16985 -11605 16991 -11553
rect 17473 -11695 17525 -11689
rect 17473 -11759 17525 -11747
rect 17473 -11817 17525 -11811
tri 17473 -11826 17482 -11817 ne
rect 17482 -11826 17525 -11817
tri 17482 -11829 17485 -11826 ne
rect 17485 -11829 17525 -11826
tri 17485 -11841 17497 -11829 ne
rect 16919 -12055 16925 -12003
rect 16977 -12055 16989 -12003
rect 17041 -12055 17047 -12003
tri 17371 -12043 17374 -12040 se
tri 17366 -12048 17371 -12043 se
rect 17371 -12048 17374 -12043
tri 17363 -12051 17366 -12048 se
rect 17366 -12051 17374 -12048
tri 17359 -12055 17363 -12051 se
rect 17363 -12055 17374 -12051
rect 16982 -13007 17012 -12055
tri 17340 -12074 17359 -12055 se
rect 17359 -12074 17374 -12055
tri 17426 -12048 17431 -12043 sw
rect 17426 -12051 17431 -12048
tri 17431 -12051 17434 -12048 sw
rect 17426 -12055 17434 -12051
tri 17434 -12055 17438 -12051 sw
rect 17426 -12074 17438 -12055
tri 17438 -12074 17457 -12055 sw
tri 17464 -12779 17497 -12746 se
rect 17497 -12779 17525 -11829
rect 17572 -11814 17578 -11762
rect 17630 -11814 17642 -11762
rect 17694 -11814 17700 -11762
rect 17982 -11808 18014 -10969
rect 18468 -11676 18496 -7583
rect 18368 -11728 18374 -11676
rect 18426 -11728 18438 -11676
rect 18490 -11728 18496 -11676
tri 18540 -11728 18546 -11722 se
rect 18546 -11728 18574 -7438
rect 18626 -9220 18654 -7261
rect 21068 -7307 21120 -7304
rect 20404 -7359 20410 -7307
rect 20462 -7359 20474 -7307
rect 20526 -7310 21120 -7307
rect 20526 -7359 21068 -7310
rect 21068 -7374 21120 -7362
rect 20051 -7454 20057 -7402
rect 20109 -7454 20121 -7402
rect 20173 -7403 20179 -7402
rect 20173 -7409 21040 -7403
rect 20173 -7454 20988 -7409
rect 21068 -7432 21120 -7426
rect 20988 -7473 21040 -7461
rect 20988 -7531 21040 -7525
rect 18903 -7718 18909 -7666
rect 18961 -7718 18973 -7666
rect 19025 -7718 19031 -7666
tri 18903 -7721 18906 -7718 ne
rect 18906 -7721 19028 -7718
tri 19028 -7721 19031 -7718 nw
rect 21236 -7710 21288 -7704
tri 18906 -7755 18940 -7721 ne
rect 18602 -9226 18654 -9220
rect 18602 -9290 18654 -9278
rect 18602 -9348 18654 -9342
rect 18682 -8383 18734 -8377
rect 18682 -8447 18734 -8435
rect 18682 -10572 18734 -8499
rect 18940 -8644 18984 -7721
tri 18984 -7765 19028 -7721 nw
rect 20587 -7773 20593 -7721
rect 20645 -7773 20657 -7721
rect 20709 -7762 21236 -7721
rect 20709 -7773 21288 -7762
rect 21236 -7774 21288 -7773
rect 19719 -7885 19725 -7833
rect 19777 -7885 19789 -7833
rect 19841 -7885 19847 -7833
rect 20587 -7854 20593 -7802
rect 20645 -7854 20657 -7802
rect 20709 -7808 21199 -7802
rect 20709 -7854 21147 -7808
tri 18984 -8644 19008 -8620 sw
rect 19819 -8644 19847 -7885
rect 21236 -7832 21288 -7826
rect 21147 -7872 21199 -7860
rect 21147 -7930 21199 -7924
rect 19994 -8142 20003 -8141
rect 20059 -8142 20126 -8141
rect 20182 -8142 20249 -8141
rect 20305 -8142 20314 -8141
rect 19994 -8194 20000 -8142
rect 20059 -8194 20086 -8142
rect 20223 -8194 20249 -8142
rect 20308 -8194 20314 -8142
rect 19994 -8197 20003 -8194
rect 20059 -8197 20126 -8194
rect 20182 -8197 20249 -8194
rect 20305 -8197 20314 -8194
rect 19994 -8216 20314 -8197
rect 19994 -8268 20000 -8216
rect 20052 -8268 20086 -8216
rect 20138 -8268 20171 -8216
rect 20223 -8268 20256 -8216
rect 20308 -8268 20314 -8216
rect 19994 -8287 20314 -8268
rect 19994 -8290 20003 -8287
rect 20059 -8290 20126 -8287
rect 20182 -8290 20249 -8287
rect 20305 -8290 20314 -8287
rect 19994 -8342 20000 -8290
rect 20059 -8342 20086 -8290
rect 20223 -8342 20249 -8290
rect 20308 -8342 20314 -8290
rect 19994 -8343 20003 -8342
rect 20059 -8343 20126 -8342
rect 20182 -8343 20249 -8342
rect 20305 -8343 20314 -8342
tri 18910 -8675 18940 -8645 se
rect 18940 -8660 19008 -8644
tri 19008 -8660 19024 -8644 sw
rect 18940 -8667 19024 -8660
tri 19024 -8667 19031 -8660 sw
rect 18940 -8675 19031 -8667
tri 19031 -8675 19039 -8667 sw
rect 18910 -8727 18916 -8675
rect 18968 -8727 18981 -8675
rect 19033 -8727 19039 -8675
rect 19763 -8696 19769 -8644
rect 19821 -8696 19833 -8644
rect 19885 -8696 19891 -8644
rect 22755 -8667 22761 -8615
rect 22813 -8667 22825 -8615
rect 22877 -8667 22883 -8615
rect 19454 -9144 20370 -9116
rect 19109 -9299 19161 -9293
rect 18763 -9371 18815 -9365
rect 18763 -9435 18815 -9423
rect 18763 -9766 18815 -9487
rect 18763 -9830 18815 -9818
rect 18763 -9888 18815 -9882
rect 19109 -9368 19161 -9351
rect 19109 -9437 19161 -9420
rect 19109 -9764 19161 -9489
rect 19454 -9399 19506 -9144
tri 19506 -9178 19540 -9144 nw
tri 20290 -9178 20324 -9144 ne
rect 19454 -9463 19506 -9451
rect 19109 -9828 19161 -9816
rect 19109 -9886 19161 -9880
rect 19355 -9765 19407 -9759
rect 19355 -9829 19407 -9817
rect 19355 -10028 19407 -9881
rect 19454 -9766 19506 -9515
rect 19718 -9268 19752 -9216
rect 19804 -9268 19816 -9216
rect 19868 -9268 19874 -9216
rect 19454 -9830 19506 -9818
rect 19454 -9893 19506 -9882
rect 19556 -9604 19684 -9598
rect 19608 -9656 19626 -9604
rect 19678 -9656 19684 -9604
rect 19556 -9670 19684 -9656
rect 19608 -9722 19626 -9670
rect 19678 -9722 19684 -9670
tri 19407 -10028 19425 -10010 sw
rect 19355 -10032 19425 -10028
tri 19355 -10060 19383 -10032 ne
rect 19383 -10060 19425 -10032
tri 19425 -10060 19457 -10028 sw
tri 19383 -10080 19403 -10060 ne
rect 19403 -10080 19457 -10060
tri 19403 -10082 19405 -10080 ne
rect 18638 -10624 18644 -10572
rect 18696 -10624 18708 -10572
rect 18760 -10624 18766 -10572
tri 19396 -11384 19405 -11375 se
rect 19405 -11384 19457 -10080
rect 19556 -10577 19684 -9722
rect 19608 -10629 19626 -10577
rect 19678 -10629 19684 -10577
rect 19556 -10643 19684 -10629
rect 19608 -10695 19626 -10643
rect 19678 -10695 19684 -10643
rect 19556 -10701 19684 -10695
tri 19384 -11396 19396 -11384 se
rect 19396 -11396 19457 -11384
tri 19457 -11396 19458 -11395 sw
tri 19371 -11409 19384 -11396 se
rect 19384 -11409 19458 -11396
tri 19458 -11409 19471 -11396 sw
rect 19343 -11461 19349 -11409
rect 19401 -11461 19413 -11409
rect 19465 -11461 19471 -11409
tri 19687 -11461 19718 -11430 se
rect 19718 -11461 19746 -9268
tri 19746 -9302 19780 -9268 nw
rect 20045 -9314 20097 -9308
rect 20045 -9384 20097 -9366
tri 19684 -11464 19687 -11461 se
rect 19687 -11464 19746 -11461
tri 19684 -11550 19718 -11516 ne
tri 19572 -11607 19603 -11576 sw
tri 19532 -11610 19535 -11607 se
rect 19572 -11610 19603 -11607
tri 19603 -11610 19606 -11607 sw
tri 18512 -11756 18540 -11728 se
rect 18540 -11756 18574 -11728
tri 18574 -11756 18608 -11722 sw
tri 18014 -11808 18020 -11802 sw
rect 18484 -11808 18490 -11756
rect 18542 -11808 18554 -11756
rect 18606 -11808 18612 -11756
tri 17871 -11814 17875 -11810 se
rect 17572 -11826 17622 -11814
tri 17622 -11826 17634 -11814 nw
tri 17859 -11826 17871 -11814 se
rect 17871 -11826 17875 -11814
rect 17572 -11829 17619 -11826
tri 17619 -11829 17622 -11826 nw
tri 17856 -11829 17859 -11826 se
rect 17859 -11829 17875 -11826
rect 17572 -11844 17604 -11829
tri 17604 -11844 17619 -11829 nw
tri 17841 -11844 17856 -11829 se
rect 17856 -11844 17875 -11829
tri 17903 -11826 17919 -11810 sw
rect 17982 -11826 18020 -11808
tri 18020 -11826 18038 -11808 sw
rect 17903 -11829 17919 -11826
tri 17919 -11829 17922 -11826 sw
rect 17982 -11829 18038 -11826
tri 18038 -11829 18041 -11826 sw
rect 17903 -11844 17922 -11829
tri 17922 -11844 17937 -11829 sw
rect 17982 -11836 18041 -11829
tri 18041 -11836 18048 -11829 sw
rect 17572 -12323 17600 -11844
tri 17600 -11848 17604 -11844 nw
rect 17982 -11888 18014 -11836
tri 19698 -11888 19718 -11868 se
rect 19718 -11888 19746 -11464
rect 19775 -9399 19827 -9393
tri 20002 -9436 20045 -9393 se
tri 19996 -9442 20002 -9436 se
rect 20002 -9442 20097 -9436
rect 19775 -9467 19827 -9451
tri 19982 -9456 19996 -9442 se
rect 19996 -9456 20048 -9442
tri 20048 -9456 20062 -9442 nw
rect 19775 -9764 19827 -9519
tri 19916 -9522 19982 -9456 se
tri 19982 -9522 20048 -9456 nw
rect 19775 -9828 19827 -9816
rect 19775 -11559 19827 -9880
tri 19890 -9548 19916 -9522 se
rect 19916 -9548 19956 -9522
tri 19956 -9548 19982 -9522 nw
rect 19890 -10164 19936 -9548
tri 19936 -9568 19956 -9548 nw
rect 20324 -9665 20370 -9144
rect 20322 -9671 20374 -9665
rect 22787 -9694 22839 -8667
rect 23065 -8923 23299 -8904
rect 23065 -8927 23074 -8923
rect 23065 -8979 23071 -8927
rect 23130 -8979 23154 -8923
rect 23210 -8979 23234 -8923
rect 23290 -8927 23299 -8923
rect 23293 -8979 23299 -8927
rect 23065 -9002 23299 -8979
rect 20322 -9735 20374 -9723
rect 20322 -9793 20374 -9787
rect 22776 -9746 22839 -9694
rect 19990 -10084 19999 -10028
rect 20055 -10084 20084 -10028
rect 20140 -10084 20169 -10028
rect 20225 -10084 20253 -10028
rect 20309 -10084 20318 -10028
rect 19990 -10106 20318 -10084
rect 19990 -10108 20000 -10106
rect 20052 -10108 20086 -10106
rect 20138 -10108 20171 -10106
rect 20223 -10108 20256 -10106
rect 20308 -10108 20318 -10106
tri 19936 -10164 19939 -10161 sw
rect 19990 -10164 19999 -10108
rect 20055 -10164 20084 -10108
rect 20140 -10164 20169 -10108
rect 20225 -10164 20253 -10108
rect 20309 -10164 20318 -10108
rect 22776 -10046 22821 -9746
rect 23402 -9873 23454 -9867
rect 23402 -9939 23454 -9925
tri 22821 -10046 22839 -10028 sw
rect 22776 -10098 22839 -10046
tri 22776 -10109 22787 -10098 ne
rect 19890 -10195 19939 -10164
tri 19939 -10195 19970 -10164 sw
rect 19890 -10247 19896 -10195
rect 19948 -10247 19960 -10195
rect 20012 -10247 20018 -10195
rect 19990 -10468 19999 -10412
rect 20055 -10468 20084 -10412
rect 20140 -10468 20169 -10412
rect 20225 -10468 20253 -10412
rect 20309 -10468 20318 -10412
rect 19990 -10490 20318 -10468
rect 19990 -10492 20000 -10490
rect 20052 -10492 20086 -10490
rect 20138 -10492 20171 -10490
rect 20223 -10492 20256 -10490
rect 20308 -10492 20318 -10490
rect 19990 -10548 19999 -10492
rect 20055 -10548 20084 -10492
rect 20140 -10548 20169 -10492
rect 20225 -10548 20253 -10492
rect 20309 -10548 20318 -10492
rect 22787 -10518 22839 -10098
rect 23228 -10198 23234 -10146
rect 23286 -10198 23298 -10146
rect 23350 -10198 23356 -10146
tri 23269 -10232 23303 -10198 ne
rect 23303 -10200 23356 -10198
rect 23054 -10257 23236 -10236
rect 23054 -10259 23079 -10257
rect 23054 -10311 23060 -10259
rect 23054 -10313 23079 -10311
rect 23135 -10313 23159 -10257
rect 23215 -10259 23236 -10257
rect 23230 -10311 23236 -10259
rect 23215 -10313 23236 -10311
rect 23054 -10334 23236 -10313
rect 22787 -10570 23094 -10518
rect 20082 -11386 20091 -11330
rect 20147 -11332 20172 -11330
rect 20228 -11332 20253 -11330
rect 20154 -11384 20172 -11332
rect 20232 -11384 20253 -11332
rect 20147 -11386 20172 -11384
rect 20228 -11386 20253 -11384
rect 20309 -11386 20318 -11330
tri 20051 -11456 20055 -11452 sw
tri 20007 -11472 20023 -11456 se
tri 19993 -11486 20007 -11472 se
rect 20007 -11486 20023 -11472
rect 20051 -11472 20055 -11456
tri 20055 -11472 20071 -11456 sw
rect 20051 -11486 20071 -11472
tri 20071 -11486 20085 -11472 sw
rect 23042 -11506 23094 -10570
rect 23127 -11269 23263 -11263
rect 23127 -11272 23137 -11269
rect 23189 -11321 23201 -11269
rect 23253 -11272 23263 -11269
rect 23183 -11328 23207 -11321
rect 23127 -11344 23263 -11328
rect 23127 -11396 23137 -11344
rect 23189 -11396 23201 -11344
rect 23253 -11396 23263 -11344
rect 23127 -11413 23263 -11396
rect 23183 -11420 23207 -11413
rect 23127 -11472 23137 -11469
rect 23189 -11472 23201 -11420
rect 23253 -11472 23263 -11469
rect 23127 -11478 23263 -11472
rect 22966 -11558 22972 -11506
rect 23024 -11558 23036 -11506
rect 23088 -11558 23094 -11506
rect 19775 -11623 19827 -11611
rect 19775 -11681 19827 -11675
rect 23042 -11760 23094 -11558
rect 23303 -11599 23355 -10200
tri 23355 -10201 23356 -10200 nw
rect 23402 -11517 23454 -9991
rect 27137 -11276 27146 -11220
rect 27202 -11276 27252 -11220
rect 27308 -11276 27358 -11220
rect 27414 -11276 27423 -11220
rect 27137 -11344 27423 -11276
rect 27137 -11400 27146 -11344
rect 27202 -11400 27252 -11344
rect 27308 -11400 27358 -11344
rect 27414 -11400 27423 -11344
rect 23401 -11569 23407 -11517
rect 23459 -11569 23471 -11517
rect 23523 -11569 23529 -11517
rect 23249 -11651 23255 -11599
rect 23307 -11651 23319 -11599
rect 23371 -11651 23377 -11599
rect 24082 -11715 24088 -11663
rect 24140 -11715 24152 -11663
rect 24204 -11715 24210 -11663
rect 28005 -11682 28014 -11626
rect 28070 -11629 28095 -11626
rect 28151 -11629 28175 -11626
rect 28070 -11681 28091 -11629
rect 28151 -11681 28167 -11629
rect 28070 -11682 28095 -11681
rect 28151 -11682 28175 -11681
rect 28231 -11682 28240 -11626
rect 28005 -11703 28240 -11682
rect 23042 -11797 23809 -11760
rect 23909 -11772 23915 -11720
rect 23967 -11772 23979 -11720
rect 24031 -11772 24037 -11720
tri 23042 -11808 23053 -11797 ne
rect 23053 -11808 23809 -11797
tri 23053 -11812 23057 -11808 ne
rect 23057 -11812 23809 -11808
rect 17982 -11919 18017 -11888
tri 18017 -11919 18048 -11888 nw
tri 19667 -11919 19698 -11888 se
rect 19698 -11919 19746 -11888
tri 19746 -11919 19787 -11878 sw
tri 20912 -11919 20939 -11892 ne
rect 20939 -11919 20946 -11892
rect 22790 -11919 22796 -11867
rect 22848 -11919 22860 -11867
rect 22912 -11919 22918 -11867
tri 17600 -12323 17605 -12318 sw
rect 17572 -12352 17605 -12323
tri 17605 -12352 17634 -12323 sw
rect 17572 -12404 17578 -12352
rect 17630 -12404 17642 -12352
rect 17694 -12404 17700 -12352
rect 17572 -12407 17631 -12404
tri 17631 -12407 17634 -12404 nw
rect 17572 -12410 17628 -12407
tri 17628 -12410 17631 -12407 nw
tri 17525 -12779 17542 -12762 sw
rect 17414 -12831 17420 -12779
rect 17472 -12831 17484 -12779
rect 17536 -12831 17542 -12779
rect 17572 -12972 17600 -12410
tri 17600 -12438 17628 -12410 nw
tri 17936 -12887 17982 -12841 se
rect 17982 -12855 18014 -11919
tri 18014 -11922 18017 -11919 nw
tri 19664 -11922 19667 -11919 se
rect 19667 -11922 19787 -11919
tri 19663 -11923 19664 -11922 se
rect 19664 -11923 19787 -11922
tri 19787 -11923 19791 -11919 sw
tri 20939 -11923 20943 -11919 ne
rect 20943 -11923 20946 -11919
tri 22835 -11923 22839 -11919 ne
rect 22839 -11923 22918 -11919
rect 19663 -11975 19669 -11923
rect 19721 -11975 19733 -11923
rect 19785 -11975 19791 -11923
tri 20943 -11926 20946 -11923 ne
tri 22839 -11926 22842 -11923 ne
rect 22842 -11926 22918 -11923
tri 22842 -11928 22844 -11926 ne
rect 22844 -11928 22918 -11926
tri 22844 -11934 22850 -11928 ne
rect 22850 -11934 22918 -11928
tri 22918 -11934 22924 -11928 sw
tri 22850 -11941 22857 -11934 ne
rect 22857 -11941 22924 -11934
tri 22924 -11941 22931 -11934 sw
tri 22857 -11975 22891 -11941 ne
rect 22891 -11975 22931 -11941
tri 22931 -11975 22965 -11941 sw
tri 22891 -11986 22902 -11975 ne
rect 22902 -11986 22965 -11975
tri 22965 -11986 22976 -11975 sw
tri 22902 -11996 22912 -11986 ne
rect 22912 -11996 22976 -11986
tri 22976 -11996 22986 -11986 sw
tri 22912 -12002 22918 -11996 ne
rect 22918 -12002 22986 -11996
tri 22918 -12015 22931 -12002 ne
rect 22931 -12015 22986 -12002
tri 22986 -12015 23005 -11996 sw
tri 22931 -12048 22964 -12015 ne
rect 22964 -12048 23005 -12015
tri 23005 -12048 23038 -12015 sw
tri 22964 -12051 22967 -12048 ne
rect 22967 -12051 23038 -12048
tri 23038 -12051 23041 -12048 sw
tri 22967 -12089 23005 -12051 ne
rect 23005 -12089 23041 -12051
tri 23041 -12089 23079 -12051 sw
tri 23005 -12103 23019 -12089 ne
rect 23019 -12103 23079 -12089
tri 23079 -12103 23093 -12089 sw
tri 23019 -12105 23021 -12103 ne
rect 23021 -12105 23093 -12103
tri 23093 -12105 23095 -12103 sw
tri 23021 -12157 23073 -12105 ne
rect 23073 -12157 23095 -12105
tri 23095 -12157 23147 -12105 sw
tri 23073 -12163 23079 -12157 ne
rect 23079 -12163 23147 -12157
tri 23147 -12163 23153 -12157 sw
tri 23079 -12169 23085 -12163 ne
rect 23085 -12169 23153 -12163
tri 23153 -12169 23159 -12163 sw
tri 23085 -12221 23137 -12169 ne
rect 23137 -12221 23159 -12169
tri 23159 -12221 23211 -12169 sw
tri 23137 -12225 23141 -12221 ne
rect 23141 -12225 23211 -12221
tri 23211 -12225 23215 -12221 sw
tri 23141 -12237 23153 -12225 ne
rect 23153 -12237 23215 -12225
tri 23215 -12237 23227 -12225 sw
tri 23153 -12241 23157 -12237 ne
rect 23157 -12241 23227 -12237
tri 23157 -12259 23175 -12241 ne
rect 22632 -12355 22684 -12349
rect 18423 -12462 18429 -12410
rect 18481 -12411 18508 -12410
rect 18560 -12411 18586 -12410
rect 18638 -12411 18664 -12410
rect 18716 -12411 18742 -12410
rect 18492 -12462 18508 -12411
rect 18716 -12462 18730 -12411
rect 18794 -12462 18800 -12410
rect 18423 -12467 18436 -12462
rect 18492 -12467 18534 -12462
rect 18590 -12467 18632 -12462
rect 18688 -12467 18730 -12462
rect 18786 -12467 18800 -12462
rect 18423 -12503 18800 -12467
rect 22632 -12419 22684 -12407
rect 22632 -12477 22684 -12471
rect 23175 -12352 23227 -12241
rect 23757 -12271 23809 -11812
rect 23980 -12141 24008 -11772
rect 24082 -12071 24110 -11715
rect 28005 -11755 28014 -11703
rect 28066 -11755 28091 -11703
rect 28143 -11755 28167 -11703
rect 28219 -11755 28240 -11703
rect 24139 -11826 24145 -11774
rect 24197 -11826 24209 -11774
rect 24261 -11777 25445 -11774
tri 25445 -11777 25448 -11774 sw
rect 28005 -11776 28240 -11755
rect 24261 -11826 25448 -11777
tri 25448 -11826 25497 -11777 sw
tri 25439 -11829 25442 -11826 ne
rect 25442 -11829 25497 -11826
tri 25497 -11829 25500 -11826 sw
tri 25442 -11834 25447 -11829 ne
rect 25447 -11834 25500 -11829
tri 25500 -11834 25505 -11829 sw
rect 28005 -11832 28014 -11776
rect 28070 -11777 28095 -11776
rect 28151 -11777 28175 -11776
rect 28070 -11829 28091 -11777
rect 28151 -11829 28167 -11777
rect 28070 -11832 28095 -11829
rect 28151 -11832 28175 -11829
rect 28231 -11832 28240 -11776
tri 25447 -11854 25467 -11834 ne
rect 25467 -11854 25505 -11834
rect 24158 -11906 24164 -11854
rect 24216 -11906 24228 -11854
rect 24280 -11873 24286 -11854
tri 25467 -11862 25475 -11854 ne
rect 25475 -11862 25505 -11854
tri 25505 -11862 25533 -11834 sw
tri 26098 -11862 26126 -11834 se
rect 26126 -11862 27734 -11834
tri 27734 -11862 27762 -11834 sw
tri 25475 -11865 25478 -11862 ne
rect 25478 -11865 25533 -11862
tri 25533 -11865 25536 -11862 sw
tri 26095 -11865 26098 -11862 se
rect 26098 -11865 26128 -11862
tri 25478 -11867 25480 -11865 ne
rect 25480 -11867 25609 -11865
rect 24696 -11873 24702 -11867
rect 24280 -11906 24702 -11873
rect 24696 -11919 24702 -11906
rect 24754 -11919 24766 -11867
rect 24818 -11919 24824 -11867
tri 25480 -11884 25497 -11867 ne
rect 25497 -11884 25609 -11867
tri 25497 -11890 25503 -11884 ne
rect 25503 -11890 25609 -11884
tri 25503 -11917 25530 -11890 ne
rect 25530 -11917 25609 -11890
rect 25661 -11917 25673 -11865
rect 25725 -11917 25731 -11865
tri 26070 -11890 26095 -11865 se
rect 26095 -11890 26128 -11865
tri 26128 -11890 26156 -11862 nw
tri 27710 -11890 27738 -11862 ne
rect 27738 -11890 27762 -11862
tri 26043 -11917 26070 -11890 se
rect 26070 -11917 26084 -11890
tri 26041 -11919 26043 -11917 se
rect 26043 -11919 26084 -11917
tri 26026 -11934 26041 -11919 se
rect 26041 -11934 26084 -11919
tri 26084 -11934 26128 -11890 nw
tri 27738 -11914 27762 -11890 ne
tri 27762 -11914 27814 -11862 sw
tri 27762 -11934 27782 -11914 ne
rect 27782 -11934 27814 -11914
rect 24140 -11986 24146 -11934
rect 24198 -11986 24210 -11934
rect 24262 -11949 24581 -11934
tri 24581 -11949 24596 -11934 sw
tri 26012 -11948 26026 -11934 se
rect 26026 -11948 26070 -11934
tri 26070 -11948 26084 -11934 nw
tri 27782 -11948 27796 -11934 ne
rect 27796 -11948 27814 -11934
tri 26011 -11949 26012 -11948 se
rect 26012 -11949 26069 -11948
tri 26069 -11949 26070 -11948 nw
tri 27796 -11949 27797 -11948 ne
rect 27797 -11949 27814 -11948
rect 24262 -11962 24596 -11949
rect 24262 -11986 24268 -11962
tri 24557 -11986 24581 -11962 ne
rect 24581 -11986 24596 -11962
tri 24581 -11996 24591 -11986 ne
rect 24591 -11996 24596 -11986
rect 24298 -12048 24304 -11996
rect 24356 -12048 24368 -11996
rect 24420 -12001 24529 -11996
tri 24529 -12001 24534 -11996 sw
tri 24591 -12001 24596 -11996 ne
tri 24596 -12001 24648 -11949 sw
tri 25982 -11978 26011 -11949 se
rect 26011 -11966 26052 -11949
tri 26052 -11966 26069 -11949 nw
tri 27797 -11966 27814 -11949 ne
tri 27814 -11966 27866 -11914 sw
rect 26011 -11973 26045 -11966
tri 26045 -11973 26052 -11966 nw
tri 26118 -11973 26125 -11966 se
rect 26125 -11973 27119 -11966
tri 27119 -11973 27126 -11966 sw
tri 27814 -11973 27821 -11966 ne
rect 27821 -11973 27866 -11966
rect 26011 -11978 26017 -11973
tri 25434 -12001 25457 -11978 se
rect 25457 -12001 26017 -11978
tri 26017 -12001 26045 -11973 nw
tri 26090 -12001 26118 -11973 se
rect 26118 -11994 27126 -11973
rect 26118 -12001 26129 -11994
rect 24420 -12035 24534 -12001
tri 24534 -12035 24568 -12001 sw
tri 24596 -12035 24630 -12001 ne
rect 24630 -12035 24648 -12001
rect 24420 -12048 24568 -12035
tri 24531 -12051 24534 -12048 ne
rect 24534 -12051 24568 -12048
tri 24568 -12051 24584 -12035 sw
tri 24630 -12051 24646 -12035 ne
rect 24646 -12051 24648 -12035
tri 24648 -12051 24698 -12001 sw
tri 25429 -12006 25434 -12001 se
rect 25434 -12006 26012 -12001
tri 26012 -12006 26017 -12001 nw
tri 26085 -12006 26090 -12001 se
rect 26090 -12006 26129 -12001
tri 25384 -12051 25429 -12006 se
rect 25429 -12022 25464 -12006
tri 25464 -12022 25480 -12006 nw
tri 26069 -12022 26085 -12006 se
rect 26085 -12022 26129 -12006
tri 26129 -12022 26157 -11994 nw
tri 27098 -12022 27126 -11994 ne
tri 27126 -12001 27154 -11973 sw
tri 27821 -12001 27849 -11973 ne
rect 27849 -12001 27866 -11973
rect 27126 -12022 27154 -12001
tri 27154 -12022 27175 -12001 sw
tri 27849 -12018 27866 -12001 ne
tri 27866 -12018 27918 -11966 sw
rect 25429 -12026 25460 -12022
tri 25460 -12026 25464 -12022 nw
tri 26065 -12026 26069 -12022 se
rect 26069 -12026 26125 -12022
tri 26125 -12026 26129 -12022 nw
tri 27126 -12026 27130 -12022 ne
rect 27130 -12026 27175 -12022
rect 25429 -12051 25435 -12026
tri 25435 -12051 25460 -12026 nw
tri 26040 -12051 26065 -12026 se
rect 26065 -12051 26100 -12026
tri 26100 -12051 26125 -12026 nw
tri 27130 -12043 27147 -12026 ne
tri 24534 -12053 24536 -12051 ne
rect 24536 -12053 24584 -12051
tri 24584 -12053 24586 -12051 sw
tri 24646 -12053 24648 -12051 ne
rect 24648 -12053 24698 -12051
tri 24698 -12053 24700 -12051 sw
tri 25382 -12053 25384 -12051 se
rect 25384 -12053 25433 -12051
tri 25433 -12053 25435 -12051 nw
tri 26038 -12053 26040 -12051 se
rect 26040 -12053 26065 -12051
tri 24082 -12089 24100 -12071 ne
rect 24100 -12089 24110 -12071
tri 24110 -12089 24146 -12053 sw
tri 24536 -12085 24568 -12053 ne
rect 24568 -12085 24586 -12053
tri 24586 -12085 24618 -12053 sw
tri 24648 -12085 24680 -12053 ne
rect 24680 -12085 24700 -12053
tri 24568 -12089 24572 -12085 ne
rect 24572 -12089 24618 -12085
tri 24618 -12089 24622 -12085 sw
tri 24680 -12089 24684 -12085 ne
rect 24684 -12089 24700 -12085
tri 24100 -12099 24110 -12089 ne
rect 24110 -12099 24488 -12089
tri 24110 -12103 24114 -12099 ne
rect 24114 -12103 24488 -12099
tri 24488 -12103 24502 -12089 sw
tri 24572 -12103 24586 -12089 ne
rect 24586 -12103 24622 -12089
tri 24622 -12103 24636 -12089 sw
tri 24684 -12103 24698 -12089 ne
rect 24698 -12103 24700 -12089
tri 24700 -12103 24750 -12053 sw
tri 25380 -12055 25382 -12053 se
rect 25382 -12055 25431 -12053
tri 25431 -12055 25433 -12053 nw
tri 26036 -12055 26038 -12053 se
rect 26038 -12055 26065 -12053
tri 25332 -12103 25380 -12055 se
rect 25380 -12086 25400 -12055
tri 25400 -12086 25431 -12055 nw
tri 26005 -12086 26036 -12055 se
rect 26036 -12086 26065 -12055
tri 26065 -12086 26100 -12051 nw
tri 26486 -12086 26521 -12051 se
rect 26521 -12086 26684 -12051
rect 25380 -12103 25383 -12086
tri 25383 -12103 25400 -12086 nw
tri 25988 -12103 26005 -12086 se
rect 26005 -12103 26048 -12086
tri 26048 -12103 26065 -12086 nw
tri 26469 -12103 26486 -12086 se
rect 26486 -12103 26684 -12086
rect 26736 -12103 26748 -12051
rect 26800 -12103 26806 -12051
tri 24114 -12105 24116 -12103 ne
rect 24116 -12105 24502 -12103
tri 24502 -12105 24504 -12103 sw
tri 24586 -12105 24588 -12103 ne
rect 24588 -12105 24636 -12103
tri 24636 -12105 24638 -12103 sw
tri 24698 -12105 24700 -12103 ne
rect 24700 -12105 24750 -12103
tri 24750 -12105 24752 -12103 sw
tri 25330 -12105 25332 -12103 se
rect 25332 -12105 25381 -12103
tri 25381 -12105 25383 -12103 nw
tri 25986 -12105 25988 -12103 se
rect 25988 -12105 26013 -12103
tri 24116 -12117 24128 -12105 ne
rect 24128 -12117 24504 -12105
tri 24462 -12130 24475 -12117 ne
rect 24475 -12130 24504 -12117
tri 24504 -12130 24529 -12105 sw
tri 24588 -12130 24613 -12105 ne
rect 24613 -12130 24638 -12105
tri 24638 -12130 24663 -12105 sw
tri 24700 -12130 24725 -12105 ne
rect 24725 -12130 24816 -12105
tri 24008 -12141 24019 -12130 sw
tri 24475 -12133 24478 -12130 ne
rect 24478 -12133 24529 -12130
tri 24529 -12133 24532 -12130 sw
tri 24613 -12133 24616 -12130 ne
rect 24616 -12133 24663 -12130
tri 24663 -12133 24666 -12130 sw
tri 24725 -12133 24728 -12130 ne
rect 24728 -12133 24816 -12130
tri 24478 -12141 24486 -12133 ne
rect 24486 -12141 24532 -12133
tri 24532 -12141 24540 -12133 sw
tri 24616 -12135 24618 -12133 ne
rect 24618 -12135 24666 -12133
tri 24666 -12135 24668 -12133 sw
tri 24728 -12135 24730 -12133 ne
rect 24730 -12135 24816 -12133
tri 24618 -12141 24624 -12135 ne
rect 24624 -12141 24668 -12135
tri 24668 -12141 24674 -12135 sw
tri 24730 -12141 24736 -12135 ne
rect 24736 -12141 24816 -12135
rect 23980 -12153 24019 -12141
tri 23980 -12157 23984 -12153 ne
rect 23984 -12157 24019 -12153
tri 24019 -12157 24035 -12141 sw
tri 24486 -12143 24488 -12141 ne
rect 24488 -12143 24540 -12141
tri 24488 -12157 24502 -12143 ne
rect 24502 -12156 24540 -12143
tri 24540 -12156 24555 -12141 sw
tri 24624 -12156 24639 -12141 ne
rect 24639 -12156 24674 -12141
tri 24674 -12156 24689 -12141 sw
tri 24736 -12156 24751 -12141 ne
rect 24502 -12157 24555 -12156
tri 24555 -12157 24556 -12156 sw
tri 24639 -12157 24640 -12156 ne
rect 24640 -12157 24689 -12156
tri 24689 -12157 24690 -12156 sw
rect 24751 -12157 24816 -12141
rect 24868 -12157 24880 -12105
rect 24932 -12129 24938 -12105
tri 25329 -12106 25330 -12105 se
rect 25330 -12106 25380 -12105
tri 25380 -12106 25381 -12105 nw
tri 25985 -12106 25986 -12105 se
rect 25986 -12106 26013 -12105
tri 25306 -12129 25329 -12106 se
rect 25329 -12129 25357 -12106
tri 25357 -12129 25380 -12106 nw
tri 25962 -12129 25985 -12106 se
rect 25985 -12129 26013 -12106
rect 24932 -12138 25348 -12129
tri 25348 -12138 25357 -12129 nw
tri 25953 -12138 25962 -12129 se
rect 25962 -12138 26013 -12129
tri 26013 -12138 26048 -12103 nw
tri 26434 -12138 26469 -12103 se
rect 26469 -12138 26484 -12103
tri 26484 -12138 26519 -12103 nw
rect 24932 -12146 25340 -12138
tri 25340 -12146 25348 -12138 nw
tri 25945 -12146 25953 -12138 se
rect 25953 -12146 26005 -12138
tri 26005 -12146 26013 -12138 nw
tri 26426 -12146 26434 -12138 se
rect 26434 -12146 26476 -12138
tri 26476 -12146 26484 -12138 nw
rect 24932 -12157 25329 -12146
tri 25329 -12157 25340 -12146 nw
tri 25934 -12157 25945 -12146 se
rect 25945 -12157 25982 -12146
tri 23984 -12169 23996 -12157 ne
rect 23996 -12169 24035 -12157
tri 24035 -12169 24047 -12157 sw
tri 24502 -12169 24514 -12157 ne
rect 24514 -12169 24556 -12157
tri 24556 -12169 24568 -12157 sw
tri 24640 -12169 24652 -12157 ne
rect 24652 -12169 24690 -12157
tri 24690 -12169 24702 -12157 sw
tri 25922 -12169 25934 -12157 se
rect 25934 -12169 25982 -12157
tri 25982 -12169 26005 -12146 nw
tri 26419 -12153 26426 -12146 se
rect 26426 -12153 26469 -12146
tri 26469 -12153 26476 -12146 nw
tri 26403 -12169 26419 -12153 se
rect 26419 -12169 26453 -12153
tri 26453 -12169 26469 -12153 nw
rect 27147 -12169 27175 -12026
tri 27866 -12070 27918 -12018 ne
tri 27918 -12054 27954 -12018 sw
rect 27918 -12070 27954 -12054
tri 27954 -12070 27970 -12054 sw
tri 27918 -12106 27954 -12070 ne
rect 27954 -12082 27970 -12070
tri 27970 -12082 27982 -12070 sw
rect 27954 -12138 27982 -12082
tri 23996 -12192 24019 -12169 ne
rect 24019 -12192 24047 -12169
tri 24047 -12192 24070 -12169 sw
tri 24514 -12187 24532 -12169 ne
rect 24532 -12187 24568 -12169
tri 24568 -12187 24586 -12169 sw
tri 24652 -12185 24668 -12169 ne
rect 24668 -12179 24702 -12169
tri 24702 -12179 24712 -12169 sw
rect 25663 -12179 25669 -12169
rect 24668 -12185 24712 -12179
tri 24712 -12185 24718 -12179 sw
tri 25460 -12185 25466 -12179 se
rect 25466 -12185 25669 -12179
tri 24668 -12187 24670 -12185 ne
rect 24670 -12187 25669 -12185
tri 24532 -12192 24537 -12187 ne
rect 24537 -12192 24586 -12187
tri 24586 -12192 24591 -12187 sw
tri 24670 -12192 24675 -12187 ne
rect 24675 -12192 25669 -12187
tri 24019 -12220 24047 -12192 ne
rect 24047 -12220 24446 -12192
tri 24424 -12221 24425 -12220 ne
rect 24425 -12221 24446 -12220
tri 24446 -12221 24475 -12192 sw
tri 24537 -12221 24566 -12192 ne
rect 24566 -12221 24591 -12192
tri 24591 -12221 24620 -12192 sw
tri 24675 -12213 24696 -12192 ne
rect 24696 -12207 25669 -12192
rect 24696 -12213 25484 -12207
tri 25484 -12213 25490 -12207 nw
rect 25663 -12221 25669 -12207
rect 25721 -12221 25733 -12169
rect 25785 -12179 25972 -12169
tri 25972 -12179 25982 -12169 nw
tri 26393 -12179 26403 -12169 se
rect 26403 -12179 26443 -12169
tri 26443 -12179 26453 -12169 nw
rect 25785 -12207 25944 -12179
tri 25944 -12207 25972 -12179 nw
tri 26369 -12203 26393 -12179 se
rect 26393 -12203 26419 -12179
tri 26419 -12203 26443 -12179 nw
tri 26365 -12207 26369 -12203 se
rect 26369 -12207 26415 -12203
tri 26415 -12207 26419 -12203 nw
rect 25785 -12213 25938 -12207
tri 25938 -12213 25944 -12207 nw
tri 26359 -12213 26365 -12207 se
rect 26365 -12213 26409 -12207
tri 26409 -12213 26415 -12207 nw
rect 25785 -12221 25930 -12213
tri 25930 -12221 25938 -12213 nw
tri 26351 -12221 26359 -12213 se
rect 26359 -12221 26401 -12213
tri 26401 -12221 26409 -12213 nw
rect 27110 -12221 27116 -12169
rect 27168 -12221 27180 -12169
rect 27232 -12221 27238 -12169
rect 27954 -12190 27960 -12138
rect 28012 -12190 28028 -12138
rect 28080 -12190 28086 -12138
tri 24425 -12225 24429 -12221 ne
rect 24429 -12225 24475 -12221
tri 24475 -12225 24479 -12221 sw
tri 24566 -12225 24570 -12221 ne
rect 24570 -12225 24620 -12221
tri 24620 -12225 24624 -12221 sw
tri 26347 -12225 26351 -12221 se
rect 26351 -12225 26397 -12221
tri 26397 -12225 26401 -12221 nw
tri 24429 -12231 24435 -12225 ne
rect 24435 -12231 24479 -12225
tri 24479 -12231 24485 -12225 sw
tri 24570 -12231 24576 -12225 ne
rect 24576 -12231 24624 -12225
tri 24624 -12231 24630 -12225 sw
tri 26341 -12231 26347 -12225 se
rect 26347 -12231 26391 -12225
tri 26391 -12231 26397 -12225 nw
tri 24435 -12241 24445 -12231 ne
rect 24445 -12241 24485 -12231
tri 24485 -12241 24495 -12231 sw
tri 24576 -12241 24586 -12231 ne
rect 24586 -12241 24630 -12231
tri 24630 -12241 24640 -12231 sw
tri 26331 -12241 26341 -12231 se
rect 26341 -12241 26381 -12231
tri 26381 -12241 26391 -12231 nw
tri 24445 -12242 24446 -12241 ne
rect 24446 -12242 24495 -12241
tri 24446 -12271 24475 -12242 ne
rect 24475 -12249 24495 -12242
tri 24495 -12249 24503 -12241 sw
tri 24586 -12249 24594 -12241 ne
rect 24594 -12249 24802 -12241
rect 24475 -12271 24503 -12249
rect 23727 -12323 23733 -12271
rect 23785 -12323 23797 -12271
rect 23849 -12323 23855 -12271
tri 24475 -12281 24485 -12271 ne
rect 24485 -12281 24503 -12271
tri 24503 -12281 24535 -12249 sw
tri 24594 -12269 24614 -12249 ne
rect 24614 -12269 24802 -12249
tri 24485 -12293 24497 -12281 ne
rect 24497 -12293 24535 -12281
tri 24535 -12293 24547 -12281 sw
rect 24796 -12293 24802 -12269
rect 24854 -12293 24868 -12241
rect 24920 -12293 24926 -12241
tri 25005 -12293 25049 -12249 se
rect 25049 -12293 25055 -12241
rect 25107 -12293 25119 -12241
rect 25171 -12293 25177 -12241
tri 26329 -12243 26331 -12241 se
rect 26331 -12243 26379 -12241
tri 26379 -12243 26381 -12241 nw
tri 26323 -12249 26329 -12243 se
rect 26329 -12249 26373 -12243
tri 26373 -12249 26379 -12243 nw
tri 26319 -12253 26323 -12249 se
rect 26323 -12253 26369 -12249
tri 26369 -12253 26373 -12249 nw
tri 26279 -12293 26319 -12253 se
rect 26319 -12293 26329 -12253
tri 26329 -12293 26369 -12253 nw
tri 24497 -12295 24499 -12293 ne
rect 24499 -12295 24547 -12293
tri 24547 -12295 24549 -12293 sw
tri 25003 -12295 25005 -12293 se
rect 25005 -12295 25049 -12293
tri 25049 -12295 25051 -12293 nw
tri 26277 -12295 26279 -12293 se
rect 26279 -12295 26327 -12293
tri 26327 -12295 26329 -12293 nw
rect 27730 -12295 27736 -12243
rect 27788 -12295 27800 -12243
rect 27852 -12295 27858 -12243
rect 27966 -12277 27972 -12225
rect 28024 -12277 28036 -12225
rect 28088 -12277 28094 -12225
tri 24499 -12323 24527 -12295 ne
rect 24527 -12323 24549 -12295
tri 24527 -12331 24535 -12323 ne
rect 24535 -12331 24549 -12323
tri 24549 -12331 24585 -12295 sw
tri 24967 -12331 25003 -12295 se
rect 25003 -12331 25013 -12295
tri 25013 -12331 25049 -12295 nw
tri 26269 -12303 26277 -12295 se
rect 26277 -12303 26319 -12295
tri 26319 -12303 26327 -12295 nw
tri 26241 -12331 26269 -12303 se
rect 26269 -12331 26291 -12303
tri 26291 -12331 26319 -12303 nw
tri 24535 -12359 24563 -12331 ne
rect 24563 -12359 24985 -12331
tri 24985 -12359 25013 -12331 nw
tri 26219 -12353 26241 -12331 se
rect 26241 -12353 26269 -12331
tri 26269 -12353 26291 -12331 nw
tri 26213 -12359 26219 -12353 se
rect 26219 -12359 26263 -12353
tri 26263 -12359 26269 -12353 nw
tri 26187 -12385 26213 -12359 se
rect 26213 -12385 26219 -12359
rect 23175 -12419 23227 -12404
rect 24288 -12437 24294 -12385
rect 24346 -12437 24358 -12385
rect 24410 -12392 24523 -12385
tri 24523 -12392 24530 -12385 sw
tri 26180 -12392 26187 -12385 se
rect 26187 -12392 26219 -12385
rect 24410 -12403 26219 -12392
tri 26219 -12403 26263 -12359 nw
rect 24410 -12420 26202 -12403
tri 26202 -12420 26219 -12403 nw
rect 24410 -12437 24416 -12420
tri 24416 -12437 24433 -12420 nw
rect 23175 -12477 23227 -12471
rect 18423 -12516 18436 -12503
rect 18492 -12516 18534 -12503
rect 18590 -12516 18632 -12503
rect 18688 -12516 18730 -12503
rect 18786 -12516 18800 -12503
rect 18423 -12568 18429 -12516
rect 18492 -12559 18508 -12516
rect 18716 -12559 18730 -12516
rect 18481 -12568 18508 -12559
rect 18560 -12568 18586 -12559
rect 18638 -12568 18664 -12559
rect 18716 -12568 18742 -12559
rect 18794 -12568 18800 -12516
rect 23066 -12558 23072 -12506
rect 23066 -12562 23075 -12558
rect 23131 -12562 23164 -12506
rect 23220 -12562 23252 -12506
rect 23311 -12558 23317 -12506
rect 23308 -12562 23317 -12558
rect 23066 -12584 23317 -12562
rect 23066 -12636 23072 -12584
rect 23124 -12586 23166 -12584
rect 23218 -12586 23259 -12584
rect 23066 -12642 23075 -12636
rect 23131 -12642 23164 -12586
rect 23220 -12642 23252 -12586
rect 23311 -12636 23317 -12584
rect 23308 -12642 23317 -12636
tri 17982 -12887 18014 -12855 nw
tri 17899 -12924 17936 -12887 se
rect 17936 -12924 17951 -12887
tri 17951 -12918 17982 -12887 nw
rect 16960 -13013 17012 -13007
rect 16960 -13077 17012 -13065
rect 17562 -12978 17614 -12972
rect 17562 -13042 17614 -13030
rect 17562 -13100 17614 -13094
rect 17899 -13097 17951 -12924
rect 16960 -13135 17012 -13129
rect 16374 -13194 16380 -13142
rect 16432 -13194 16444 -13142
rect 16496 -13149 16565 -13142
tri 16565 -13149 16572 -13142 nw
tri 16732 -13149 16739 -13142 se
rect 16739 -13149 16775 -13142
rect 16496 -13161 16553 -13149
tri 16553 -13161 16565 -13149 nw
tri 16720 -13161 16732 -13149 se
rect 16732 -13161 16775 -13149
rect 16496 -13162 16552 -13161
tri 16552 -13162 16553 -13161 nw
tri 16719 -13162 16720 -13161 se
rect 16720 -13162 16775 -13161
rect 16496 -13194 16520 -13162
tri 16520 -13194 16552 -13162 nw
rect 16607 -13214 16613 -13162
rect 16665 -13214 16677 -13162
rect 16729 -13214 16775 -13162
rect 17899 -13161 17951 -13149
rect 17899 -13219 17951 -13213
<< via2 >>
rect 17870 -7970 17874 -7925
rect 17874 -7970 17926 -7925
rect 18008 -7970 18013 -7925
rect 18013 -7970 18064 -7925
rect 17870 -7981 17926 -7970
rect 18008 -7981 18064 -7970
rect 17870 -8040 17874 -8010
rect 17874 -8040 17926 -8010
rect 18008 -8040 18013 -8010
rect 18013 -8040 18064 -8010
rect 17870 -8058 17926 -8040
rect 18008 -8058 18064 -8040
rect 17870 -8066 17874 -8058
rect 17874 -8066 17926 -8058
rect 17870 -8110 17874 -8095
rect 17874 -8110 17926 -8095
rect 18008 -8066 18013 -8058
rect 18013 -8066 18064 -8058
rect 18008 -8110 18013 -8095
rect 18013 -8110 18064 -8095
rect 17870 -8151 17926 -8110
rect 18008 -8151 18064 -8110
rect 17870 -8236 17926 -8180
rect 18008 -8236 18064 -8180
rect 17870 -8321 17926 -8265
rect 18008 -8321 18064 -8265
rect 17870 -8406 17926 -8350
rect 18008 -8406 18064 -8350
rect 17870 -8491 17926 -8435
rect 18008 -8491 18064 -8435
rect 17870 -8576 17926 -8520
rect 18008 -8576 18064 -8520
rect 17870 -8662 17926 -8606
rect 18008 -8662 18064 -8606
rect 17871 -9135 17922 -9087
rect 17922 -9135 17927 -9087
rect 17977 -9135 17996 -9087
rect 17996 -9135 18018 -9087
rect 18018 -9135 18033 -9087
rect 17871 -9143 17927 -9135
rect 17977 -9143 18033 -9135
rect 17871 -9216 17922 -9169
rect 17922 -9216 17927 -9169
rect 17977 -9216 17996 -9169
rect 17996 -9216 18018 -9169
rect 18018 -9216 18033 -9169
rect 17871 -9225 17927 -9216
rect 17977 -9225 18033 -9216
rect 17871 -9297 17922 -9251
rect 17922 -9297 17927 -9251
rect 17977 -9297 17996 -9251
rect 17996 -9297 18018 -9251
rect 18018 -9297 18033 -9251
rect 17871 -9307 17927 -9297
rect 17977 -9307 18033 -9297
rect 17871 -9389 17927 -9333
rect 17977 -9389 18033 -9333
rect 17871 -9471 17927 -9415
rect 17977 -9471 18033 -9415
rect 17871 -9553 17927 -9497
rect 17977 -9553 18033 -9497
rect 17871 -9635 17927 -9579
rect 17977 -9635 18033 -9579
rect 17871 -9717 17927 -9661
rect 17977 -9717 18033 -9661
rect 17871 -9799 17927 -9743
rect 17977 -9799 18033 -9743
rect 17871 -9881 17927 -9825
rect 17977 -9881 18033 -9825
rect 17871 -9963 17927 -9907
rect 17977 -9963 18033 -9907
rect 17871 -10045 17927 -9989
rect 17977 -10045 18033 -9989
rect 17871 -10127 17927 -10071
rect 17977 -10127 18033 -10071
rect 17871 -10208 17927 -10153
rect 17977 -10208 18033 -10153
rect 17871 -10209 17874 -10208
rect 17874 -10209 17926 -10208
rect 17926 -10209 17927 -10208
rect 17977 -10209 17994 -10208
rect 17994 -10209 18009 -10208
rect 18009 -10209 18033 -10208
rect 17871 -10260 17874 -10235
rect 17874 -10260 17926 -10235
rect 17926 -10260 17927 -10235
rect 17977 -10260 17994 -10235
rect 17994 -10260 18009 -10235
rect 18009 -10260 18033 -10235
rect 17871 -10291 17927 -10260
rect 17977 -10291 18033 -10260
rect 17871 -10374 17927 -10318
rect 17977 -10374 18033 -10318
rect 17871 -10457 17927 -10401
rect 17977 -10457 18033 -10401
rect 20003 -8142 20059 -8141
rect 20126 -8142 20182 -8141
rect 20249 -8142 20305 -8141
rect 20003 -8194 20052 -8142
rect 20052 -8194 20059 -8142
rect 20126 -8194 20138 -8142
rect 20138 -8194 20171 -8142
rect 20171 -8194 20182 -8142
rect 20249 -8194 20256 -8142
rect 20256 -8194 20305 -8142
rect 20003 -8197 20059 -8194
rect 20126 -8197 20182 -8194
rect 20249 -8197 20305 -8194
rect 20003 -8290 20059 -8287
rect 20126 -8290 20182 -8287
rect 20249 -8290 20305 -8287
rect 20003 -8342 20052 -8290
rect 20052 -8342 20059 -8290
rect 20126 -8342 20138 -8290
rect 20138 -8342 20171 -8290
rect 20171 -8342 20182 -8290
rect 20249 -8342 20256 -8290
rect 20256 -8342 20305 -8290
rect 20003 -8343 20059 -8342
rect 20126 -8343 20182 -8342
rect 20249 -8343 20305 -8342
rect 23074 -8927 23130 -8923
rect 23074 -8979 23123 -8927
rect 23123 -8979 23130 -8927
rect 23154 -8927 23210 -8923
rect 23154 -8979 23156 -8927
rect 23156 -8979 23208 -8927
rect 23208 -8979 23210 -8927
rect 23234 -8927 23290 -8923
rect 23234 -8979 23241 -8927
rect 23241 -8979 23290 -8927
rect 19999 -10080 20000 -10028
rect 20000 -10080 20052 -10028
rect 20052 -10080 20055 -10028
rect 19999 -10084 20055 -10080
rect 20084 -10080 20086 -10028
rect 20086 -10080 20138 -10028
rect 20138 -10080 20140 -10028
rect 20084 -10084 20140 -10080
rect 20169 -10080 20171 -10028
rect 20171 -10080 20223 -10028
rect 20223 -10080 20225 -10028
rect 20169 -10084 20225 -10080
rect 20253 -10080 20256 -10028
rect 20256 -10080 20308 -10028
rect 20308 -10080 20309 -10028
rect 20253 -10084 20309 -10080
rect 19999 -10158 20000 -10108
rect 20000 -10158 20052 -10108
rect 20052 -10158 20055 -10108
rect 19999 -10164 20055 -10158
rect 20084 -10158 20086 -10108
rect 20086 -10158 20138 -10108
rect 20138 -10158 20140 -10108
rect 20084 -10164 20140 -10158
rect 20169 -10158 20171 -10108
rect 20171 -10158 20223 -10108
rect 20223 -10158 20225 -10108
rect 20169 -10164 20225 -10158
rect 20253 -10158 20256 -10108
rect 20256 -10158 20308 -10108
rect 20308 -10158 20309 -10108
rect 20253 -10164 20309 -10158
rect 19999 -10464 20000 -10412
rect 20000 -10464 20052 -10412
rect 20052 -10464 20055 -10412
rect 19999 -10468 20055 -10464
rect 20084 -10464 20086 -10412
rect 20086 -10464 20138 -10412
rect 20138 -10464 20140 -10412
rect 20084 -10468 20140 -10464
rect 20169 -10464 20171 -10412
rect 20171 -10464 20223 -10412
rect 20223 -10464 20225 -10412
rect 20169 -10468 20225 -10464
rect 20253 -10464 20256 -10412
rect 20256 -10464 20308 -10412
rect 20308 -10464 20309 -10412
rect 20253 -10468 20309 -10464
rect 19999 -10542 20000 -10492
rect 20000 -10542 20052 -10492
rect 20052 -10542 20055 -10492
rect 19999 -10548 20055 -10542
rect 20084 -10542 20086 -10492
rect 20086 -10542 20138 -10492
rect 20138 -10542 20140 -10492
rect 20084 -10548 20140 -10542
rect 20169 -10542 20171 -10492
rect 20171 -10542 20223 -10492
rect 20223 -10542 20225 -10492
rect 20169 -10548 20225 -10542
rect 20253 -10542 20256 -10492
rect 20256 -10542 20308 -10492
rect 20308 -10542 20309 -10492
rect 20253 -10548 20309 -10542
rect 23079 -10259 23135 -10257
rect 23079 -10311 23112 -10259
rect 23112 -10311 23135 -10259
rect 23079 -10313 23135 -10311
rect 23159 -10259 23215 -10257
rect 23159 -10311 23178 -10259
rect 23178 -10311 23215 -10259
rect 23159 -10313 23215 -10311
rect 20091 -11332 20147 -11330
rect 20172 -11332 20228 -11330
rect 20253 -11332 20309 -11330
rect 20091 -11384 20102 -11332
rect 20102 -11384 20147 -11332
rect 20172 -11384 20180 -11332
rect 20180 -11384 20228 -11332
rect 20253 -11384 20257 -11332
rect 20257 -11384 20309 -11332
rect 20091 -11386 20147 -11384
rect 20172 -11386 20228 -11384
rect 20253 -11386 20309 -11384
rect 23127 -11321 23137 -11272
rect 23137 -11321 23183 -11272
rect 23207 -11321 23253 -11272
rect 23253 -11321 23263 -11272
rect 23127 -11328 23183 -11321
rect 23207 -11328 23263 -11321
rect 23127 -11420 23183 -11413
rect 23207 -11420 23263 -11413
rect 23127 -11469 23137 -11420
rect 23137 -11469 23183 -11420
rect 23207 -11469 23253 -11420
rect 23253 -11469 23263 -11420
rect 27146 -11276 27202 -11220
rect 27252 -11276 27308 -11220
rect 27358 -11276 27414 -11220
rect 27146 -11400 27202 -11344
rect 27252 -11400 27308 -11344
rect 27358 -11400 27414 -11344
rect 28014 -11629 28070 -11626
rect 28095 -11629 28151 -11626
rect 28175 -11629 28231 -11626
rect 28014 -11681 28066 -11629
rect 28066 -11681 28070 -11629
rect 28095 -11681 28143 -11629
rect 28143 -11681 28151 -11629
rect 28175 -11681 28219 -11629
rect 28219 -11681 28231 -11629
rect 28014 -11682 28070 -11681
rect 28095 -11682 28151 -11681
rect 28175 -11682 28231 -11681
rect 18436 -12462 18481 -12411
rect 18481 -12462 18492 -12411
rect 18534 -12462 18560 -12411
rect 18560 -12462 18586 -12411
rect 18586 -12462 18590 -12411
rect 18632 -12462 18638 -12411
rect 18638 -12462 18664 -12411
rect 18664 -12462 18688 -12411
rect 18730 -12462 18742 -12411
rect 18742 -12462 18786 -12411
rect 18436 -12467 18492 -12462
rect 18534 -12467 18590 -12462
rect 18632 -12467 18688 -12462
rect 18730 -12467 18786 -12462
rect 28014 -11777 28070 -11776
rect 28095 -11777 28151 -11776
rect 28175 -11777 28231 -11776
rect 28014 -11829 28066 -11777
rect 28066 -11829 28070 -11777
rect 28095 -11829 28143 -11777
rect 28143 -11829 28151 -11777
rect 28175 -11829 28219 -11777
rect 28219 -11829 28231 -11777
rect 28014 -11832 28070 -11829
rect 28095 -11832 28151 -11829
rect 28175 -11832 28231 -11829
rect 18436 -12516 18492 -12503
rect 18534 -12516 18590 -12503
rect 18632 -12516 18688 -12503
rect 18730 -12516 18786 -12503
rect 18436 -12559 18481 -12516
rect 18481 -12559 18492 -12516
rect 18534 -12559 18560 -12516
rect 18560 -12559 18586 -12516
rect 18586 -12559 18590 -12516
rect 18632 -12559 18638 -12516
rect 18638 -12559 18664 -12516
rect 18664 -12559 18688 -12516
rect 18730 -12559 18742 -12516
rect 18742 -12559 18786 -12516
rect 23075 -12558 23124 -12506
rect 23124 -12558 23131 -12506
rect 23075 -12562 23131 -12558
rect 23164 -12558 23166 -12506
rect 23166 -12558 23218 -12506
rect 23218 -12558 23220 -12506
rect 23164 -12562 23220 -12558
rect 23252 -12558 23259 -12506
rect 23259 -12558 23308 -12506
rect 23252 -12562 23308 -12558
rect 23075 -12636 23124 -12586
rect 23124 -12636 23131 -12586
rect 23075 -12642 23131 -12636
rect 23164 -12636 23166 -12586
rect 23166 -12636 23218 -12586
rect 23218 -12636 23220 -12586
rect 23164 -12642 23220 -12636
rect 23252 -12636 23259 -12586
rect 23259 -12636 23308 -12586
rect 23252 -12642 23308 -12636
<< metal3 >>
rect 17844 -7925 18073 -7911
rect 17844 -7981 17870 -7925
rect 17926 -7981 18008 -7925
rect 18064 -7981 18073 -7925
rect 17844 -8010 18073 -7981
rect 17844 -8066 17870 -8010
rect 17926 -8066 18008 -8010
rect 18064 -8066 18073 -8010
rect 17844 -8095 18073 -8066
rect 17844 -8151 17870 -8095
rect 17926 -8151 18008 -8095
rect 18064 -8151 18073 -8095
rect 17844 -8180 18073 -8151
rect 17844 -8236 17870 -8180
rect 17926 -8236 18008 -8180
rect 18064 -8236 18073 -8180
rect 17844 -8265 18073 -8236
rect 17844 -8321 17870 -8265
rect 17926 -8321 18008 -8265
rect 18064 -8321 18073 -8265
rect 17844 -8350 18073 -8321
rect 19998 -8141 20310 -8136
rect 19998 -8197 20003 -8141
rect 20059 -8197 20126 -8141
rect 20182 -8197 20249 -8141
rect 20305 -8197 20310 -8141
rect 19998 -8287 20310 -8197
rect 19998 -8343 20003 -8287
rect 20059 -8343 20126 -8287
rect 20182 -8343 20249 -8287
rect 20305 -8343 20310 -8287
rect 19998 -8348 20310 -8343
rect 17844 -8406 17870 -8350
rect 17926 -8406 18008 -8350
rect 18064 -8406 18073 -8350
rect 17844 -8435 18073 -8406
rect 17844 -8491 17870 -8435
rect 17926 -8491 18008 -8435
rect 18064 -8491 18073 -8435
rect 17844 -8520 18073 -8491
tri 17828 -8576 17844 -8560 se
rect 17844 -8576 17870 -8520
rect 17926 -8576 18008 -8520
rect 18064 -8576 18073 -8520
tri 17798 -8606 17828 -8576 se
rect 17828 -8606 18073 -8576
tri 17742 -8662 17798 -8606 se
rect 17798 -8662 17870 -8606
rect 17926 -8662 18008 -8606
rect 18064 -8662 18073 -8606
tri 17727 -8677 17742 -8662 se
rect 17742 -8677 18073 -8662
tri 17694 -8710 17727 -8677 se
rect 17727 -8710 17962 -8677
rect 17694 -9077 17962 -8710
tri 17962 -8788 18073 -8677 nw
rect 23051 -8923 23318 -8902
rect 23051 -8979 23074 -8923
rect 23130 -8979 23154 -8923
rect 23210 -8979 23234 -8923
rect 23290 -8979 23318 -8923
tri 17962 -9077 18038 -9001 sw
rect 17694 -9079 18038 -9077
tri 17694 -9087 17702 -9079 ne
rect 17702 -9087 18038 -9079
tri 17702 -9143 17758 -9087 ne
rect 17758 -9143 17871 -9087
rect 17927 -9143 17977 -9087
rect 18033 -9143 18038 -9087
tri 17758 -9169 17784 -9143 ne
rect 17784 -9169 18038 -9143
tri 17784 -9179 17794 -9169 ne
rect 17794 -9225 17871 -9169
rect 17927 -9225 17977 -9169
rect 18033 -9225 18038 -9169
rect 17794 -9251 18038 -9225
rect 17794 -9307 17871 -9251
rect 17927 -9307 17977 -9251
rect 18033 -9307 18038 -9251
rect 17794 -9333 18038 -9307
rect 17794 -9389 17871 -9333
rect 17927 -9389 17977 -9333
rect 18033 -9389 18038 -9333
rect 17794 -9415 18038 -9389
rect 17794 -9471 17871 -9415
rect 17927 -9471 17977 -9415
rect 18033 -9471 18038 -9415
rect 17794 -9497 18038 -9471
rect 17794 -9553 17871 -9497
rect 17927 -9553 17977 -9497
rect 18033 -9553 18038 -9497
rect 17794 -9579 18038 -9553
rect 17794 -9635 17871 -9579
rect 17927 -9635 17977 -9579
rect 18033 -9635 18038 -9579
rect 17794 -9661 18038 -9635
rect 17794 -9717 17871 -9661
rect 17927 -9717 17977 -9661
rect 18033 -9717 18038 -9661
rect 17794 -9743 18038 -9717
rect 17794 -9799 17871 -9743
rect 17927 -9799 17977 -9743
rect 18033 -9799 18038 -9743
rect 17794 -9825 18038 -9799
rect 17794 -9881 17871 -9825
rect 17927 -9881 17977 -9825
rect 18033 -9881 18038 -9825
rect 17794 -9907 18038 -9881
rect 17794 -9963 17871 -9907
rect 17927 -9963 17977 -9907
rect 18033 -9963 18038 -9907
rect 17794 -9989 18038 -9963
rect 17794 -10045 17871 -9989
rect 17927 -10045 17977 -9989
rect 18033 -10045 18038 -9989
rect 17794 -10071 18038 -10045
rect 17794 -10127 17871 -10071
rect 17927 -10127 17977 -10071
rect 18033 -10127 18038 -10071
rect 17794 -10153 18038 -10127
rect 17794 -10209 17871 -10153
rect 17927 -10209 17977 -10153
rect 18033 -10209 18038 -10153
rect 17794 -10235 18038 -10209
rect 17794 -10291 17871 -10235
rect 17927 -10291 17977 -10235
rect 18033 -10291 18038 -10235
rect 17794 -10318 18038 -10291
rect 17794 -10374 17871 -10318
rect 17927 -10374 17977 -10318
rect 18033 -10374 18038 -10318
rect 17794 -10401 18038 -10374
rect 17794 -10457 17871 -10401
rect 17927 -10457 17977 -10401
rect 18033 -10457 18038 -10401
tri 17536 -13573 17794 -13315 se
rect 17794 -13417 18038 -10457
rect 18423 -12411 18800 -9996
rect 19994 -10028 20314 -10023
rect 19994 -10084 19999 -10028
rect 20055 -10084 20084 -10028
rect 20140 -10084 20169 -10028
rect 20225 -10084 20253 -10028
rect 20309 -10084 20314 -10028
rect 19994 -10108 20314 -10084
rect 19994 -10164 19999 -10108
rect 20055 -10164 20084 -10108
rect 20140 -10164 20169 -10108
rect 20225 -10164 20253 -10108
rect 20309 -10164 20314 -10108
rect 19994 -10169 20314 -10164
rect 23051 -10257 23318 -8979
rect 23051 -10313 23079 -10257
rect 23135 -10313 23159 -10257
rect 23215 -10313 23318 -10257
rect 19994 -10412 20314 -10407
rect 19994 -10468 19999 -10412
rect 20055 -10468 20084 -10412
rect 20140 -10468 20169 -10412
rect 20225 -10468 20253 -10412
rect 20309 -10468 20314 -10412
rect 19994 -10492 20314 -10468
rect 19994 -10548 19999 -10492
rect 20055 -10548 20084 -10492
rect 20140 -10548 20169 -10492
rect 20225 -10548 20253 -10492
rect 20309 -10548 20314 -10492
rect 19994 -10553 20314 -10548
rect 23051 -11272 23318 -10313
rect 28003 -9119 28325 -9113
rect 28067 -9183 28089 -9119
rect 28153 -9183 28175 -9119
rect 28239 -9183 28261 -9119
rect 28003 -9199 28325 -9183
rect 28067 -9263 28089 -9199
rect 28153 -9263 28175 -9199
rect 28239 -9263 28261 -9199
rect 28003 -9279 28325 -9263
rect 28067 -9343 28089 -9279
rect 28153 -9343 28175 -9279
rect 28239 -9343 28261 -9279
rect 28003 -9359 28325 -9343
rect 28067 -9423 28089 -9359
rect 28153 -9423 28175 -9359
rect 28239 -9423 28261 -9359
rect 28003 -9439 28325 -9423
rect 28067 -9503 28089 -9439
rect 28153 -9503 28175 -9439
rect 28239 -9503 28261 -9439
rect 28003 -9519 28325 -9503
rect 28067 -9583 28089 -9519
rect 28153 -9583 28175 -9519
rect 28239 -9583 28261 -9519
rect 28003 -9599 28325 -9583
rect 28067 -9663 28089 -9599
rect 28153 -9663 28175 -9599
rect 28239 -9663 28261 -9599
rect 28003 -9679 28325 -9663
rect 28067 -9743 28089 -9679
rect 28153 -9743 28175 -9679
rect 28239 -9743 28261 -9679
rect 28003 -9760 28325 -9743
rect 28067 -9824 28089 -9760
rect 28153 -9824 28175 -9760
rect 28239 -9824 28261 -9760
rect 28003 -9841 28325 -9824
rect 28067 -9905 28089 -9841
rect 28153 -9905 28175 -9841
rect 28239 -9905 28261 -9841
rect 28003 -9922 28325 -9905
rect 28067 -9986 28089 -9922
rect 28153 -9986 28175 -9922
rect 28239 -9986 28261 -9922
rect 20086 -11330 20314 -11325
rect 20086 -11386 20091 -11330
rect 20147 -11386 20172 -11330
rect 20228 -11386 20253 -11330
rect 20309 -11386 20314 -11330
rect 20086 -11391 20314 -11386
rect 23051 -11328 23127 -11272
rect 23183 -11328 23207 -11272
rect 23263 -11328 23318 -11272
rect 18423 -12467 18436 -12411
rect 18492 -12467 18534 -12411
rect 18590 -12467 18632 -12411
rect 18688 -12467 18730 -12411
rect 18786 -12467 18800 -12411
rect 18423 -12503 18800 -12467
rect 23051 -11413 23318 -11328
rect 23051 -11469 23127 -11413
rect 23183 -11469 23207 -11413
rect 23263 -11469 23318 -11413
rect 23051 -12490 23318 -11469
rect 27137 -11220 27423 -11215
rect 27137 -11276 27146 -11220
rect 27202 -11276 27252 -11220
rect 27308 -11276 27358 -11220
rect 27414 -11276 27423 -11220
rect 27137 -11344 27423 -11276
rect 27137 -11400 27146 -11344
rect 27202 -11400 27252 -11344
rect 27308 -11400 27358 -11344
rect 27414 -11400 27423 -11344
rect 18423 -12559 18436 -12503
rect 18492 -12559 18534 -12503
rect 18590 -12559 18632 -12503
rect 18688 -12559 18730 -12503
rect 18786 -12559 18800 -12503
rect 18423 -12565 18800 -12559
rect 23070 -12506 23313 -12501
rect 23070 -12562 23075 -12506
rect 23131 -12562 23164 -12506
rect 23220 -12562 23252 -12506
rect 23308 -12562 23313 -12506
rect 23070 -12586 23313 -12562
rect 23070 -12642 23075 -12586
rect 23131 -12642 23164 -12586
rect 23220 -12642 23252 -12586
rect 23308 -12642 23313 -12586
rect 23070 -12647 23313 -12642
rect 17794 -13573 17882 -13417
tri 17882 -13573 18038 -13417 nw
tri 26847 -13573 27137 -13283 se
rect 27137 -13403 27423 -11400
rect 28003 -11626 28325 -9986
rect 28003 -11682 28014 -11626
rect 28070 -11682 28095 -11626
rect 28151 -11682 28175 -11626
rect 28231 -11682 28325 -11626
rect 28003 -11776 28325 -11682
rect 28003 -11832 28014 -11776
rect 28070 -11832 28095 -11776
rect 28151 -11832 28175 -11776
rect 28231 -11832 28325 -11776
rect 28003 -11837 28325 -11832
rect 27137 -13573 27299 -13403
tri 27299 -13527 27423 -13403 nw
tri 17448 -13661 17536 -13573 se
rect 17536 -13661 17794 -13573
tri 17794 -13661 17882 -13573 nw
tri 17220 -13889 17448 -13661 se
rect 17448 -13889 17566 -13661
tri 17566 -13889 17794 -13661 nw
rect 17220 -14793 17464 -13889
tri 17464 -13991 17566 -13889 nw
rect 17220 -14857 17223 -14793
rect 17287 -14857 17309 -14793
rect 17373 -14857 17395 -14793
rect 17459 -14857 17464 -14793
rect 17220 -14886 17464 -14857
rect 17220 -14950 17223 -14886
rect 17287 -14950 17309 -14886
rect 17373 -14950 17395 -14886
rect 17459 -14950 17464 -14886
rect 17220 -14980 17464 -14950
rect 17220 -15044 17223 -14980
rect 17287 -15044 17309 -14980
rect 17373 -15044 17395 -14980
rect 17459 -15044 17464 -14980
rect 17220 -15074 17464 -15044
rect 17220 -15138 17223 -15074
rect 17287 -15138 17309 -15074
rect 17373 -15138 17395 -15074
rect 17459 -15138 17464 -15074
rect 17220 -15168 17464 -15138
rect 17220 -15232 17223 -15168
rect 17287 -15232 17309 -15168
rect 17373 -15232 17395 -15168
rect 17459 -15232 17464 -15168
rect 17220 -15244 17464 -15232
<< via3 >>
rect 28003 -9183 28067 -9119
rect 28089 -9183 28153 -9119
rect 28175 -9183 28239 -9119
rect 28261 -9183 28325 -9119
rect 28003 -9263 28067 -9199
rect 28089 -9263 28153 -9199
rect 28175 -9263 28239 -9199
rect 28261 -9263 28325 -9199
rect 28003 -9343 28067 -9279
rect 28089 -9343 28153 -9279
rect 28175 -9343 28239 -9279
rect 28261 -9343 28325 -9279
rect 28003 -9423 28067 -9359
rect 28089 -9423 28153 -9359
rect 28175 -9423 28239 -9359
rect 28261 -9423 28325 -9359
rect 28003 -9503 28067 -9439
rect 28089 -9503 28153 -9439
rect 28175 -9503 28239 -9439
rect 28261 -9503 28325 -9439
rect 28003 -9583 28067 -9519
rect 28089 -9583 28153 -9519
rect 28175 -9583 28239 -9519
rect 28261 -9583 28325 -9519
rect 28003 -9663 28067 -9599
rect 28089 -9663 28153 -9599
rect 28175 -9663 28239 -9599
rect 28261 -9663 28325 -9599
rect 28003 -9743 28067 -9679
rect 28089 -9743 28153 -9679
rect 28175 -9743 28239 -9679
rect 28261 -9743 28325 -9679
rect 28003 -9824 28067 -9760
rect 28089 -9824 28153 -9760
rect 28175 -9824 28239 -9760
rect 28261 -9824 28325 -9760
rect 28003 -9905 28067 -9841
rect 28089 -9905 28153 -9841
rect 28175 -9905 28239 -9841
rect 28261 -9905 28325 -9841
rect 28003 -9986 28067 -9922
rect 28089 -9986 28153 -9922
rect 28175 -9986 28239 -9922
rect 28261 -9986 28325 -9922
rect 17223 -14857 17287 -14793
rect 17309 -14857 17373 -14793
rect 17395 -14857 17459 -14793
rect 17223 -14950 17287 -14886
rect 17309 -14950 17373 -14886
rect 17395 -14950 17459 -14886
rect 17223 -15044 17287 -14980
rect 17309 -15044 17373 -14980
rect 17395 -15044 17459 -14980
rect 17223 -15138 17287 -15074
rect 17309 -15138 17373 -15074
rect 17395 -15138 17459 -15074
rect 17223 -15232 17287 -15168
rect 17309 -15232 17373 -15168
rect 17395 -15232 17459 -15168
<< metal4 >>
rect 28002 -9119 28326 -9118
rect 28002 -9183 28003 -9119
rect 28067 -9183 28089 -9119
rect 28153 -9183 28175 -9119
rect 28239 -9183 28261 -9119
rect 28325 -9183 28326 -9119
rect 28002 -9199 28326 -9183
rect 28002 -9263 28003 -9199
rect 28067 -9263 28089 -9199
rect 28153 -9263 28175 -9199
rect 28239 -9263 28261 -9199
rect 28325 -9263 28326 -9199
rect 28002 -9279 28326 -9263
rect 28002 -9343 28003 -9279
rect 28067 -9343 28089 -9279
rect 28153 -9343 28175 -9279
rect 28239 -9343 28261 -9279
rect 28325 -9343 28326 -9279
rect 28002 -9359 28326 -9343
rect 28002 -9423 28003 -9359
rect 28067 -9423 28089 -9359
rect 28153 -9423 28175 -9359
rect 28239 -9423 28261 -9359
rect 28325 -9423 28326 -9359
rect 28002 -9439 28326 -9423
rect 28002 -9503 28003 -9439
rect 28067 -9503 28089 -9439
rect 28153 -9503 28175 -9439
rect 28239 -9503 28261 -9439
rect 28325 -9503 28326 -9439
rect 28002 -9519 28326 -9503
rect 28002 -9583 28003 -9519
rect 28067 -9583 28089 -9519
rect 28153 -9583 28175 -9519
rect 28239 -9583 28261 -9519
rect 28325 -9583 28326 -9519
rect 28002 -9599 28326 -9583
rect 28002 -9663 28003 -9599
rect 28067 -9663 28089 -9599
rect 28153 -9663 28175 -9599
rect 28239 -9663 28261 -9599
rect 28325 -9663 28326 -9599
rect 28002 -9679 28326 -9663
rect 28002 -9743 28003 -9679
rect 28067 -9743 28089 -9679
rect 28153 -9743 28175 -9679
rect 28239 -9743 28261 -9679
rect 28325 -9743 28326 -9679
rect 28002 -9760 28326 -9743
rect 28002 -9824 28003 -9760
rect 28067 -9824 28089 -9760
rect 28153 -9824 28175 -9760
rect 28239 -9824 28261 -9760
rect 28325 -9824 28326 -9760
rect 28002 -9841 28326 -9824
rect 28002 -9905 28003 -9841
rect 28067 -9905 28089 -9841
rect 28153 -9905 28175 -9841
rect 28239 -9905 28261 -9841
rect 28325 -9905 28326 -9841
rect 28002 -9922 28326 -9905
rect 28002 -9986 28003 -9922
rect 28067 -9986 28089 -9922
rect 28153 -9986 28175 -9922
rect 28239 -9986 28261 -9922
rect 28325 -9986 28326 -9922
rect 28002 -9987 28326 -9986
rect 17221 -14793 17461 -14792
rect 17221 -14857 17223 -14793
rect 17287 -14857 17309 -14793
rect 17373 -14857 17395 -14793
rect 17459 -14857 17461 -14793
rect 17221 -14886 17461 -14857
rect 17221 -14950 17223 -14886
rect 17287 -14950 17309 -14886
rect 17373 -14950 17395 -14886
rect 17459 -14950 17461 -14886
rect 17221 -14980 17461 -14950
rect 17221 -15044 17223 -14980
rect 17287 -15044 17309 -14980
rect 17373 -15044 17395 -14980
rect 17459 -15044 17461 -14980
rect 17221 -15074 17461 -15044
rect 17221 -15138 17223 -15074
rect 17287 -15138 17309 -15074
rect 17373 -15138 17395 -15074
rect 17459 -15138 17461 -15074
rect 17221 -15168 17461 -15138
rect 17221 -15232 17223 -15168
rect 17287 -15232 17309 -15168
rect 17373 -15232 17395 -15168
rect 17459 -15232 17461 -15168
rect 17221 -15233 17461 -15232
use sky130_fd_io__amx_inv1  sky130_fd_io__amx_inv1_0
timestamp 1666464484
transform -1 0 16742 0 -1 -10035
box 0 10 338 748
use sky130_fd_io__amx_inv1  sky130_fd_io__amx_inv1_1
timestamp 1666464484
transform 1 0 20176 0 -1 -9456
box 0 10 338 748
use sky130_fd_io__amx_inv1  sky130_fd_io__amx_inv1_2
timestamp 1666464484
transform 1 0 16560 0 -1 -10035
box 0 10 338 748
use sky130_fd_io__gpiov2_amux_drvr_ls  sky130_fd_io__gpiov2_amux_drvr_ls_0
timestamp 1666464484
transform 1 0 16331 0 1 -9217
box 38 24 1860 1138
use sky130_fd_io__gpiov2_amux_drvr_ls  sky130_fd_io__gpiov2_amux_drvr_ls_1
timestamp 1666464484
transform 1 0 24609 0 1 -12705
box 38 24 1860 1138
use sky130_fd_io__gpiov2_amux_drvr_ls  sky130_fd_io__gpiov2_amux_drvr_ls_2
timestamp 1666464484
transform -1 0 20092 0 1 -9217
box 38 24 1860 1138
use sky130_fd_io__gpiov2_amux_drvr_ls  sky130_fd_io__gpiov2_amux_drvr_ls_3
timestamp 1666464484
transform 1 0 16331 0 -1 -9083
box 38 24 1860 1138
use sky130_fd_io__gpiov2_amux_drvr_ls  sky130_fd_io__gpiov2_amux_drvr_ls_4
timestamp 1666464484
transform 1 0 16185 0 1 -13625
box 38 24 1860 1138
use sky130_fd_io__gpiov2_amux_drvr_ls  sky130_fd_io__gpiov2_amux_drvr_ls_5
timestamp 1666464484
transform -1 0 28283 0 1 -12705
box 38 24 1860 1138
use sky130_fd_io__gpiov2_amux_drvr_lshv2hv2  sky130_fd_io__gpiov2_amux_drvr_lshv2hv2_0
timestamp 1666464484
transform -1 0 21030 0 1 -8115
box 279 -16 4943 3838
use sky130_fd_io__gpiov2_amux_drvr_lshv2hv  sky130_fd_io__gpiov2_amux_drvr_lshv2hv_0
timestamp 1666464484
transform 1 0 17744 0 1 -8115
box -1543 -16 1692 3442
use sky130_fd_io__gpiov2_amx_inv4  sky130_fd_io__gpiov2_amx_inv4_0
timestamp 1666464484
transform 1 0 19218 0 -1 -9588
box 0 10 534 616
use sky130_fd_io__gpiov2_amx_inv4  sky130_fd_io__gpiov2_amx_inv4_1
timestamp 1666464484
transform -1 0 19400 0 -1 -9588
box 0 10 534 616
use sky130_fd_io__gpiov2_amx_inv4  sky130_fd_io__gpiov2_amx_inv4_2
timestamp 1666464484
transform -1 0 23372 0 1 -12646
box 0 10 534 616
use sky130_fd_io__gpiov2_amx_inv4  sky130_fd_io__gpiov2_amx_inv4_3
timestamp 1666464484
transform -1 0 20104 0 -1 -9588
box 0 10 534 616
use sky130_fd_io__gpiov2_amx_inv4  sky130_fd_io__gpiov2_amx_inv4_4
timestamp 1666464484
transform 1 0 22486 0 1 -12646
box 0 10 534 616
use sky130_fd_io__gpiov2_amx_inv4  sky130_fd_io__gpiov2_amx_inv4_5
timestamp 1666464484
transform -1 0 19048 0 -1 -9588
box 0 10 534 616
use sky130_fd_io__gpiov2_amx_pucsd_inv  sky130_fd_io__gpiov2_amx_pucsd_inv_0
timestamp 1666464484
transform 1 0 23189 0 1 -12655
box 1 19 1415 625
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_0
timestamp 1666464484
transform 1 0 23264 0 1 -11502
box -46 24 399 1116
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_1
timestamp 1666464484
transform -1 0 22742 0 1 -11502
box -46 24 399 1116
use sky130_fd_io__hvsbt_inv_x2  sky130_fd_io__hvsbt_inv_x2_0
timestamp 1666464484
transform 1 0 22912 0 1 -11502
box 0 24 534 1116
use sky130_fd_io__hvsbt_inv_x2  sky130_fd_io__hvsbt_inv_x2_1
timestamp 1666464484
transform 1 0 22560 0 1 -11502
box 0 24 534 1116
use sky130_fd_pr__nfet_01v8__example_55959141808576  sky130_fd_pr__nfet_01v8__example_55959141808576_0
timestamp 1666464484
transform 1 0 19943 0 1 -9509
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808577  sky130_fd_pr__nfet_01v8__example_55959141808577_0
timestamp 1666464484
transform 0 -1 17492 1 0 -10306
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808578  sky130_fd_pr__nfet_01v8__example_55959141808578_0
timestamp 1666464484
transform 0 -1 17492 1 0 -10462
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808579  sky130_fd_pr__nfet_01v8__example_55959141808579_0
timestamp 1666464484
transform 1 0 19676 0 1 -9509
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808579  sky130_fd_pr__nfet_01v8__example_55959141808579_1
timestamp 1666464484
transform -1 0 18914 0 -1 -9309
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808579  sky130_fd_pr__nfet_01v8__example_55959141808579_2
timestamp 1666464484
transform -1 0 19620 0 1 -9509
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808579  sky130_fd_pr__nfet_01v8__example_55959141808579_3
timestamp 1666464484
transform 1 0 18970 0 -1 -9309
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808572  sky130_fd_pr__pfet_01v8__example_55959141808572_0
timestamp 1666464484
transform 1 0 18313 0 1 -10530
box -1 0 401 1
use sky130_fd_pr__pfet_01v8__example_55959141808573  sky130_fd_pr__pfet_01v8__example_55959141808573_0
timestamp 1666464484
transform 1 0 17857 0 1 -10530
box -1 0 401 1
<< labels >>
flabel metal1 s 17060 -13513 17088 -13485 3 FreeSans 520 0 0 0 VSSD
port 1 nsew
flabel metal1 s 22961 -11349 22989 -11321 3 FreeSans 520 0 0 0 VSSD
port 1 nsew
flabel metal1 s 17217 -12677 17245 -12649 3 FreeSans 520 0 0 0 VDDIO_Q
port 2 nsew
flabel metal1 s 17464 -10079 17492 -10051 3 FreeSans 520 0 0 0 VSWITCH
port 3 nsew
flabel metal1 s 18501 -7072 18529 -7044 3 FreeSans 520 0 0 0 VSSA
port 4 nsew
flabel metal1 s 18925 -8000 18953 -7972 3 FreeSans 520 0 0 0 VSSA
port 4 nsew
flabel metal1 s 17759 -13207 17787 -13179 3 FreeSans 520 0 0 0 VCCD
port 5 nsew
flabel metal1 s 18158 -8801 18186 -8773 3 FreeSans 520 0 0 0 VCCD
port 5 nsew
flabel metal1 s 22906 -10546 22934 -10518 3 FreeSans 520 0 0 0 VCCD
port 5 nsew
flabel metal1 s 22462 -11144 22488 -11107 3 FreeSans 520 0 0 0 D_B
port 6 nsew
flabel metal1 s 22659 -11142 22706 -11106 3 FreeSans 520 90 0 0 D_B
port 6 nsew
flabel metal1 s 23514 -11143 23549 -11099 3 FreeSans 520 0 0 0 NMIDA_VCCD_N
port 7 nsew
flabel metal1 s 23201 -10925 23274 -10888 3 FreeSans 520 0 0 0 NMIDA_VCCD
port 8 nsew
flabel metal1 s 16798 -10755 16834 -10706 3 FreeSans 520 0 0 0 NGA_PAD_VSWITCH_H_N
port 9 nsew
flabel metal1 s 16479 -10545 16511 -10469 3 FreeSans 520 0 0 0 PD_CSD_VSWITCH_H_N
port 10 nsew
flabel metal1 s 20414 -9692 20441 -9603 3 FreeSans 520 0 0 0 NGB_PAD_VSWITCH_H_N
port 11 nsew
flabel metal1 s 19787 -9423 19815 -9395 3 FreeSans 520 0 0 0 NGA_PAD_VSWITCH_H
port 12 nsew
flabel metal1 s 18274 -10341 18302 -10313 3 FreeSans 520 0 0 0 PD_CSD_VSWITCH_H
port 13 nsew
flabel metal1 s 19121 -9835 19149 -9807 3 FreeSans 520 0 0 0 NGB_AMX_VSWITCH_H
port 14 nsew
flabel metal1 s 19481 -9423 19509 -9395 3 FreeSans 520 0 0 0 NGB_PAD_VSWITCH_H
port 15 nsew
flabel metal1 s 19777 -9256 19805 -9228 3 FreeSans 520 0 0 0 AMUX_EN_VDDIO_H_N
port 16 nsew
flabel metal1 s 18606 -9281 18634 -9253 3 FreeSans 520 90 0 0 AMUX_EN_VDDA_H_N
port 17 nsew
flabel metal1 s 23080 -10885 23108 -10857 3 FreeSans 520 0 0 0 NMIDA_ON_N
port 18 nsew
flabel metal1 s 22728 -10810 22756 -10782 3 FreeSans 520 0 0 0 D_B
port 6 nsew
flabel metal1 s 26629 -12291 26657 -12263 3 FreeSans 520 0 0 0 VCCD
port 5 nsew
flabel metal1 s 26764 -11721 26792 -11693 3 FreeSans 520 0 0 0 VDDIO_Q
port 2 nsew
flabel metal1 s 28015 -12260 28043 -12232 3 FreeSans 520 0 0 0 PU_ON_N
port 19 nsew
flabel metal1 s 27800 -12281 27828 -12253 3 FreeSans 520 0 0 0 PU_ON
port 20 nsew
flabel metal1 s 27147 -12207 27175 -12179 3 FreeSans 520 0 0 0 AMUX_EN_VDDIO_H
port 21 nsew
flabel metal1 s 16425 -13180 16453 -13152 3 FreeSans 520 0 0 0 AMUXBUSA_ON_N
port 22 nsew
flabel metal1 s 16640 -13200 16668 -13172 3 FreeSans 520 0 0 0 AMUXBUSA_ON
port 23 nsew
flabel metal1 s 16576 -9640 16604 -9612 3 FreeSans 520 0 0 0 AMUX_EN_VSWITCH_H_N
port 24 nsew
flabel metal1 s 18499 -10469 18527 -10441 3 FreeSans 520 0 0 0 VSWITCH
port 3 nsew
flabel metal1 s 20388 -7089 20416 -7061 3 FreeSans 520 0 0 0 PGB_AMX_VDDA_H_N
port 25 nsew
flabel metal1 s 18775 -9423 18803 -9395 3 FreeSans 520 0 0 0 NGA_AMX_VSWITCH_H
port 26 nsew
flabel metal1 s 18925 -9435 18953 -9407 3 FreeSans 520 0 0 0 VSSA
port 4 nsew
flabel metal1 s 19824 -8772 19852 -8744 3 FreeSans 520 0 0 0 PD_ON_N
port 27 nsew
flabel metal1 s 16434 -4653 16462 -4625 3 FreeSans 520 0 0 0 VDDA
port 28 nsew
flabel metal1 s 19419 -7347 19447 -7319 3 FreeSans 520 90 0 0 AMUX_EN_VDDA_H
port 29 nsew
flabel metal1 s 28182 -12531 28210 -12503 3 FreeSans 520 0 0 0 VSSD
port 1 nsew
flabel metal1 s 17439 -9609 17467 -9581 3 FreeSans 520 0 0 0 AMUX_EN_VSWITCH_H
port 30 nsew
flabel metal1 s 25064 -12280 25092 -12252 3 FreeSans 520 0 0 0 AMUXBUSB_ON
port 31 nsew
flabel metal1 s 23993 -12315 24065 -12272 3 FreeSans 520 180 0 0 PU_CSD_VDDIOQ_H_N
port 32 nsew
flabel metal1 s 24849 -12260 24877 -12232 3 FreeSans 520 0 0 0 AMUXBUSB_ON_N
port 33 nsew
flabel metal1 s 19609 -8792 19637 -8764 3 FreeSans 520 0 0 0 PD_ON
port 34 nsew
flabel metal1 s 23095 -12422 23123 -12394 3 FreeSans 520 180 0 0 PGB_PAD_VDDIOQ_H_N
port 35 nsew
flabel metal1 s 22734 -12422 22762 -12394 3 FreeSans 520 180 0 0 PGA_PAD_VDDIOQ_H_N
port 36 nsew
flabel metal1 s 18358 -7089 18386 -7061 3 FreeSans 520 0 0 0 PGA_AMX_VDDA_H_N
port 37 nsew
flabel comment s 18453 -8925 18453 -8925 0 FreeSans 2000 180 0 0 VSWITCH- VSSA
<< properties >>
string GDS_END 43749644
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 43606958
<< end >>
