magic
tech sky130B
magscale 1 2
timestamp 1666464484
<< obsli1 >>
rect 80 1118 214 1134
rect 80 1084 94 1118
rect 128 1084 166 1118
rect 200 1084 214 1118
rect 80 1068 214 1084
rect 44 985 78 1034
rect 44 913 78 951
rect 44 841 78 879
rect 44 769 78 807
rect 44 697 78 735
rect 44 625 78 663
rect 44 553 78 591
rect 44 481 78 519
rect 44 409 78 447
rect 44 337 78 375
rect 44 265 78 303
rect 44 193 78 231
rect 44 121 78 159
rect 44 36 78 87
rect 130 36 164 1034
rect 216 985 250 1034
rect 216 913 250 951
rect 216 841 250 879
rect 216 769 250 807
rect 216 697 250 735
rect 216 625 250 663
rect 216 553 250 591
rect 216 481 250 519
rect 216 409 250 447
rect 216 337 250 375
rect 216 265 250 303
rect 216 193 250 231
rect 216 121 250 159
rect 216 36 250 87
<< obsli1c >>
rect 94 1084 128 1118
rect 166 1084 200 1118
rect 44 951 78 985
rect 44 879 78 913
rect 44 807 78 841
rect 44 735 78 769
rect 44 663 78 697
rect 44 591 78 625
rect 44 519 78 553
rect 44 447 78 481
rect 44 375 78 409
rect 44 303 78 337
rect 44 231 78 265
rect 44 159 78 193
rect 44 87 78 121
rect 216 951 250 985
rect 216 879 250 913
rect 216 807 250 841
rect 216 735 250 769
rect 216 663 250 697
rect 216 591 250 625
rect 216 519 250 553
rect 216 447 250 481
rect 216 375 250 409
rect 216 303 250 337
rect 216 231 250 265
rect 216 159 250 193
rect 216 87 250 121
<< metal1 >>
rect 82 1118 212 1130
rect 82 1084 94 1118
rect 128 1084 166 1118
rect 200 1084 212 1118
rect 82 1072 212 1084
rect 38 985 84 1034
rect 38 951 44 985
rect 78 951 84 985
rect 38 913 84 951
rect 38 879 44 913
rect 78 879 84 913
rect 38 841 84 879
rect 38 807 44 841
rect 78 807 84 841
rect 38 769 84 807
rect 38 735 44 769
rect 78 735 84 769
rect 38 697 84 735
rect 38 663 44 697
rect 78 663 84 697
rect 38 625 84 663
rect 38 591 44 625
rect 78 591 84 625
rect 38 553 84 591
rect 38 519 44 553
rect 78 519 84 553
rect 38 481 84 519
rect 38 447 44 481
rect 78 447 84 481
rect 38 409 84 447
rect 38 375 44 409
rect 78 375 84 409
rect 38 337 84 375
rect 38 303 44 337
rect 78 303 84 337
rect 38 265 84 303
rect 38 231 44 265
rect 78 231 84 265
rect 38 193 84 231
rect 38 159 44 193
rect 78 159 84 193
rect 38 121 84 159
rect 38 87 44 121
rect 78 87 84 121
rect 38 -45 84 87
rect 210 985 256 1034
rect 210 951 216 985
rect 250 951 256 985
rect 210 913 256 951
rect 210 879 216 913
rect 250 879 256 913
rect 210 841 256 879
rect 210 807 216 841
rect 250 807 256 841
rect 210 769 256 807
rect 210 735 216 769
rect 250 735 256 769
rect 210 697 256 735
rect 210 663 216 697
rect 250 663 256 697
rect 210 625 256 663
rect 210 591 216 625
rect 250 591 256 625
rect 210 553 256 591
rect 210 519 216 553
rect 250 519 256 553
rect 210 481 256 519
rect 210 447 216 481
rect 250 447 256 481
rect 210 409 256 447
rect 210 375 216 409
rect 250 375 256 409
rect 210 337 256 375
rect 210 303 216 337
rect 250 303 256 337
rect 210 265 256 303
rect 210 231 216 265
rect 250 231 256 265
rect 210 193 256 231
rect 210 159 216 193
rect 250 159 256 193
rect 210 121 256 159
rect 210 87 216 121
rect 250 87 256 121
rect 210 -45 256 87
rect 38 -97 256 -45
<< obsm1 >>
rect 121 36 173 1034
<< metal2 >>
rect 121 904 173 1032
<< labels >>
rlabel metal2 s 121 904 173 1032 6 DRAIN
port 1 nsew
rlabel metal1 s 82 1072 212 1130 6 GATE
port 2 nsew
rlabel metal1 s 210 -45 256 1034 6 SOURCE
port 3 nsew
rlabel metal1 s 38 -45 84 1034 6 SOURCE
port 3 nsew
rlabel metal1 s 38 -97 256 -45 8 SOURCE
port 3 nsew
<< properties >>
string FIXED_BBOX 0 -97 294 1134
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 10497040
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 10488604
string device primitive
<< end >>
