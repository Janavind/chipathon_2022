magic
tech sky130A
magscale 1 2
timestamp 1666199351
<< nwell >>
rect -38 261 130 827
rect 384 261 596 827
rect 850 261 1326 827
<< pwell >>
rect 511 1050 1111 1067
rect 3 893 89 1050
rect 511 893 1245 1050
rect 511 885 1111 893
rect 601 195 1141 214
rect 3 38 89 195
rect 601 192 1245 195
rect 398 56 1245 192
rect 601 38 1245 56
rect 601 32 1141 38
<< scnmos >>
rect 590 911 620 1041
rect 676 911 706 1041
rect 762 911 792 1041
rect 848 911 878 1041
rect 1002 911 1032 1041
rect 477 82 507 166
rect 684 58 714 188
rect 770 58 800 188
rect 856 58 886 188
rect 942 58 972 188
rect 1028 58 1058 188
<< scpmoshvt >>
rect 941 618 971 776
rect 1032 618 1062 776
rect 475 297 505 497
rect 941 312 971 470
rect 1031 312 1061 470
<< ndiff >>
rect 537 1025 590 1041
rect 537 991 545 1025
rect 579 991 590 1025
rect 537 957 590 991
rect 537 923 545 957
rect 579 923 590 957
rect 537 911 590 923
rect 620 1032 676 1041
rect 620 998 631 1032
rect 665 998 676 1032
rect 620 964 676 998
rect 620 930 631 964
rect 665 930 676 964
rect 620 911 676 930
rect 706 1032 762 1041
rect 706 998 717 1032
rect 751 998 762 1032
rect 706 964 762 998
rect 706 930 717 964
rect 751 930 762 964
rect 706 911 762 930
rect 792 1032 848 1041
rect 792 998 803 1032
rect 837 998 848 1032
rect 792 964 848 998
rect 792 930 803 964
rect 837 930 848 964
rect 792 911 848 930
rect 878 1032 1002 1041
rect 878 930 889 1032
rect 991 930 1002 1032
rect 878 911 1002 930
rect 1032 1025 1085 1041
rect 1032 991 1043 1025
rect 1077 991 1085 1025
rect 1032 957 1085 991
rect 1032 923 1043 957
rect 1077 923 1085 957
rect 1032 911 1085 923
rect 627 180 684 188
rect 424 141 477 166
rect 424 107 432 141
rect 466 107 477 141
rect 424 82 477 107
rect 507 141 560 166
rect 507 107 518 141
rect 552 107 560 141
rect 507 82 560 107
rect 627 146 639 180
rect 673 146 684 180
rect 627 112 684 146
rect 627 78 639 112
rect 673 78 684 112
rect 627 58 684 78
rect 714 180 770 188
rect 714 146 725 180
rect 759 146 770 180
rect 714 112 770 146
rect 714 78 725 112
rect 759 78 770 112
rect 714 58 770 78
rect 800 112 856 188
rect 800 78 811 112
rect 845 78 856 112
rect 800 58 856 78
rect 886 180 942 188
rect 886 146 897 180
rect 931 146 942 180
rect 886 112 942 146
rect 886 78 897 112
rect 931 78 942 112
rect 886 58 942 78
rect 972 180 1028 188
rect 972 146 983 180
rect 1017 146 1028 180
rect 972 112 1028 146
rect 972 78 983 112
rect 1017 78 1028 112
rect 972 58 1028 78
rect 1058 180 1115 188
rect 1058 146 1069 180
rect 1103 146 1115 180
rect 1058 112 1115 146
rect 1058 78 1069 112
rect 1103 78 1115 112
rect 1058 58 1115 78
<< pdiff >>
rect 886 732 941 776
rect 886 698 896 732
rect 930 698 941 732
rect 886 664 941 698
rect 886 630 894 664
rect 928 630 941 664
rect 886 618 941 630
rect 971 732 1032 776
rect 971 698 984 732
rect 1018 698 1032 732
rect 971 664 1032 698
rect 971 630 984 664
rect 1018 630 1032 664
rect 971 618 1032 630
rect 1062 732 1116 776
rect 1062 698 1074 732
rect 1108 698 1116 732
rect 1062 664 1116 698
rect 1062 630 1074 664
rect 1108 630 1116 664
rect 1062 618 1116 630
rect 420 458 475 497
rect 420 424 428 458
rect 462 424 475 458
rect 420 375 475 424
rect 420 341 428 375
rect 462 341 475 375
rect 420 297 475 341
rect 505 458 560 497
rect 505 424 518 458
rect 552 424 560 458
rect 505 375 560 424
rect 886 458 941 470
rect 886 424 894 458
rect 928 424 941 458
rect 505 341 518 375
rect 552 341 560 375
rect 505 297 560 341
rect 886 375 941 424
rect 886 341 894 375
rect 928 341 941 375
rect 886 312 941 341
rect 971 458 1031 470
rect 971 424 984 458
rect 1018 424 1031 458
rect 971 375 1031 424
rect 971 341 984 375
rect 1018 341 1031 375
rect 971 312 1031 341
rect 1061 458 1116 470
rect 1061 424 1074 458
rect 1108 424 1116 458
rect 1061 375 1116 424
rect 1061 341 1074 375
rect 1108 341 1116 375
rect 1061 312 1116 341
<< ndiffc >>
rect 545 991 579 1025
rect 545 923 579 957
rect 631 998 665 1032
rect 631 930 665 964
rect 717 998 751 1032
rect 717 930 751 964
rect 803 998 837 1032
rect 803 930 837 964
rect 889 930 991 1032
rect 1043 991 1077 1025
rect 1043 923 1077 957
rect 432 107 466 141
rect 518 107 552 141
rect 639 146 673 180
rect 639 78 673 112
rect 725 146 759 180
rect 725 78 759 112
rect 811 78 845 112
rect 897 146 931 180
rect 897 78 931 112
rect 983 146 1017 180
rect 983 78 1017 112
rect 1069 146 1103 180
rect 1069 78 1103 112
<< pdiffc >>
rect 896 698 930 732
rect 894 630 928 664
rect 984 698 1018 732
rect 984 630 1018 664
rect 1074 698 1108 732
rect 1074 630 1108 664
rect 428 424 462 458
rect 428 341 462 375
rect 518 424 552 458
rect 894 424 928 458
rect 518 341 552 375
rect 894 341 928 375
rect 984 424 1018 458
rect 984 341 1018 375
rect 1074 424 1108 458
rect 1074 341 1108 375
<< psubdiff >>
rect 29 977 63 1024
rect 29 919 63 943
rect 1185 977 1219 1024
rect 1185 919 1219 943
rect 29 145 63 169
rect 29 64 63 111
rect 1185 145 1219 169
rect 1185 64 1219 111
<< nsubdiff >>
rect 29 759 63 783
rect 29 675 63 725
rect 420 715 560 743
rect 420 681 434 715
rect 468 681 512 715
rect 546 681 560 715
rect 420 654 560 681
rect 29 608 63 641
rect 1185 759 1219 783
rect 1185 675 1219 725
rect 1185 608 1219 641
<< psubdiffcont >>
rect 29 943 63 977
rect 1185 943 1219 977
rect 29 111 63 145
rect 1185 111 1219 145
<< nsubdiffcont >>
rect 29 725 63 759
rect 29 641 63 675
rect 434 681 468 715
rect 512 681 546 715
rect 1185 725 1219 759
rect 1185 641 1219 675
<< poly >>
rect 590 1041 620 1067
rect 676 1041 706 1067
rect 762 1041 792 1067
rect 848 1041 878 1067
rect 1002 1041 1032 1067
rect 590 896 620 911
rect 676 896 706 911
rect 762 896 792 911
rect 848 896 878 911
rect 590 866 878 896
rect 612 785 682 866
rect 1002 824 1032 911
rect 1142 871 1211 875
rect 1140 859 1211 871
rect 1140 825 1167 859
rect 1201 825 1211 859
rect 612 751 628 785
rect 662 751 682 785
rect 612 735 682 751
rect 788 812 1062 824
rect 788 778 804 812
rect 838 794 1062 812
rect 838 778 854 794
rect 788 644 854 778
rect 941 776 971 794
rect 1032 776 1062 794
rect 1140 803 1211 825
rect 788 610 804 644
rect 838 610 854 644
rect 788 603 854 610
rect 941 603 971 618
rect 1032 603 1062 618
rect 788 573 1062 603
rect 1140 531 1170 803
rect 475 497 505 523
rect 788 501 971 531
rect 788 499 854 501
rect 788 465 804 499
rect 838 465 854 499
rect 941 470 971 501
rect 1031 501 1170 531
rect 1031 470 1061 501
rect 788 431 854 465
rect 788 397 804 431
rect 838 397 854 431
rect 788 381 854 397
rect 475 245 505 297
rect 941 286 971 312
rect 1031 297 1061 312
rect 1140 297 1170 501
rect 592 267 658 280
rect 592 245 608 267
rect 475 233 608 245
rect 642 245 658 267
rect 642 244 726 245
rect 1031 244 1170 297
rect 642 233 972 244
rect 475 214 972 233
rect 475 202 507 214
rect 477 166 507 202
rect 684 188 714 214
rect 770 188 800 214
rect 856 188 886 214
rect 942 188 972 214
rect 1028 203 1170 244
rect 1028 188 1058 203
rect 477 21 507 82
rect 684 32 714 58
rect 770 32 800 58
rect 856 32 886 58
rect 942 32 972 58
rect 1028 32 1058 58
<< polycont >>
rect 1167 825 1201 859
rect 628 751 662 785
rect 804 778 838 812
rect 804 610 838 644
rect 804 465 838 499
rect 804 397 838 431
rect 608 233 642 267
<< locali >>
rect 0 1071 29 1105
rect 63 1071 121 1105
rect 155 1071 213 1105
rect 247 1071 305 1105
rect 339 1071 397 1105
rect 431 1071 489 1105
rect 523 1071 581 1105
rect 615 1071 673 1105
rect 707 1071 765 1105
rect 799 1071 857 1105
rect 891 1071 949 1105
rect 983 1071 1041 1105
rect 1075 1071 1133 1105
rect 1167 1071 1225 1105
rect 1259 1071 1288 1105
rect 17 977 75 1071
rect 17 943 29 977
rect 63 943 75 977
rect 17 926 75 943
rect 529 1025 581 1071
rect 529 991 545 1025
rect 579 991 581 1025
rect 529 957 581 991
rect 529 923 545 957
rect 579 923 581 957
rect 529 903 581 923
rect 615 1032 681 1037
rect 615 998 631 1032
rect 665 998 681 1032
rect 615 964 681 998
rect 615 930 631 964
rect 665 930 681 964
rect 615 865 681 930
rect 715 1032 753 1071
rect 715 998 717 1032
rect 751 998 753 1032
rect 715 964 753 998
rect 715 930 717 964
rect 751 930 753 964
rect 715 903 753 930
rect 787 1032 853 1037
rect 787 998 803 1032
rect 837 998 853 1032
rect 787 964 853 998
rect 787 930 803 964
rect 837 930 853 964
rect 787 865 853 930
rect 889 1032 991 1071
rect 889 903 991 930
rect 1027 1025 1097 1032
rect 1027 991 1043 1025
rect 1077 991 1097 1025
rect 1027 964 1097 991
rect 1173 977 1231 1071
rect 1027 957 1139 964
rect 1027 923 1043 957
rect 1077 923 1139 957
rect 1173 943 1185 977
rect 1219 943 1231 977
rect 1173 926 1231 943
rect 1027 892 1139 923
rect 1027 881 1153 892
rect 615 853 853 865
rect 1072 871 1153 881
rect 1072 859 1217 871
rect 629 831 839 853
rect 804 812 838 831
rect 17 759 75 794
rect 17 731 29 759
rect 17 697 28 731
rect 63 725 75 759
rect 612 785 678 793
rect 612 751 628 785
rect 662 751 678 785
rect 804 762 838 778
rect 1072 825 1167 859
rect 1201 825 1217 859
rect 62 697 75 725
rect 17 675 75 697
rect 17 641 29 675
rect 63 641 75 675
rect 17 597 75 641
rect 412 715 562 750
rect 412 681 434 715
rect 468 681 512 715
rect 546 681 562 715
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 378 561
rect 412 532 562 681
rect 412 467 478 532
rect 612 474 678 751
rect 882 732 944 748
rect 882 728 896 732
rect 736 698 896 728
rect 930 698 944 732
rect 736 694 944 698
rect 736 515 770 694
rect 878 664 944 694
rect 804 644 838 660
rect 878 630 894 664
rect 928 630 944 664
rect 878 617 944 630
rect 978 732 1024 748
rect 978 698 984 732
rect 1018 698 1024 732
rect 978 664 1024 698
rect 978 630 984 664
rect 1018 630 1024 664
rect 804 583 838 610
rect 804 549 928 583
rect 736 499 838 515
rect 736 481 804 499
rect 276 458 478 467
rect 276 457 428 458
rect 276 423 284 457
rect 318 423 356 457
rect 390 423 428 457
rect 462 423 478 458
rect 276 413 478 423
rect 412 375 478 413
rect 412 341 428 375
rect 462 341 478 375
rect 412 327 478 341
rect 512 458 678 474
rect 512 424 518 458
rect 552 426 678 458
rect 804 431 838 465
rect 552 424 560 426
rect 512 375 560 424
rect 512 341 518 375
rect 552 341 560 375
rect 17 145 75 162
rect 17 111 29 145
rect 63 111 75 145
rect 17 17 75 111
rect 404 141 470 179
rect 404 107 432 141
rect 466 107 470 141
rect 404 17 470 107
rect 512 141 560 341
rect 594 267 658 308
rect 594 233 608 267
rect 642 233 658 267
rect 594 214 658 233
rect 804 196 838 397
rect 894 458 928 549
rect 894 375 928 424
rect 894 325 928 341
rect 978 561 1024 630
rect 1072 732 1110 825
rect 1072 698 1074 732
rect 1108 698 1110 732
rect 1072 664 1110 698
rect 1072 630 1074 664
rect 1108 630 1110 664
rect 1072 614 1110 630
rect 1173 759 1231 791
rect 1173 725 1185 759
rect 1219 731 1231 759
rect 1173 697 1186 725
rect 1220 697 1231 731
rect 1173 675 1231 697
rect 1173 641 1185 675
rect 1219 641 1231 675
rect 1173 597 1231 641
rect 978 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 978 458 1024 527
rect 978 424 984 458
rect 1018 424 1024 458
rect 978 375 1024 424
rect 978 341 984 375
rect 1018 341 1024 375
rect 978 325 1024 341
rect 1072 458 1127 474
rect 1072 424 1074 458
rect 1108 424 1127 458
rect 1072 375 1127 424
rect 1072 341 1074 375
rect 1108 341 1127 375
rect 1072 196 1127 341
rect 723 180 933 196
rect 1067 180 1127 196
rect 512 107 518 141
rect 552 107 560 141
rect 512 75 560 107
rect 623 146 639 180
rect 673 146 689 180
rect 623 112 689 146
rect 623 78 639 112
rect 673 78 689 112
rect 623 17 689 78
rect 723 146 725 180
rect 759 146 897 180
rect 931 146 933 180
rect 723 112 761 146
rect 895 112 933 146
rect 723 78 725 112
rect 759 78 761 112
rect 723 58 761 78
rect 795 78 811 112
rect 845 78 861 112
rect 795 17 861 78
rect 895 78 897 112
rect 931 78 933 112
rect 895 58 933 78
rect 967 146 983 180
rect 1017 146 1033 180
rect 967 112 1033 146
rect 967 78 983 112
rect 1017 78 1033 112
rect 967 17 1033 78
rect 1067 146 1069 180
rect 1103 146 1127 180
rect 1067 112 1127 146
rect 1067 78 1069 112
rect 1103 78 1127 112
rect 1067 58 1127 78
rect 1173 145 1231 162
rect 1173 111 1185 145
rect 1219 111 1231 145
rect 1173 17 1231 111
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
<< viali >>
rect 29 1071 63 1105
rect 121 1071 155 1105
rect 213 1071 247 1105
rect 305 1071 339 1105
rect 397 1071 431 1105
rect 489 1071 523 1105
rect 581 1071 615 1105
rect 673 1071 707 1105
rect 765 1071 799 1105
rect 857 1071 891 1105
rect 949 1071 983 1105
rect 1041 1071 1075 1105
rect 1133 1071 1167 1105
rect 1225 1071 1259 1105
rect 28 725 29 731
rect 29 725 62 731
rect 28 697 62 725
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 284 423 318 457
rect 356 423 390 457
rect 428 424 462 457
rect 428 423 462 424
rect 1186 725 1219 731
rect 1219 725 1220 731
rect 1186 697 1220 725
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
<< metal1 >>
rect 0 1105 1288 1136
rect 0 1071 29 1105
rect 63 1071 121 1105
rect 155 1071 213 1105
rect 247 1071 305 1105
rect 339 1071 397 1105
rect 431 1071 489 1105
rect 523 1071 581 1105
rect 615 1071 673 1105
rect 707 1071 765 1105
rect 799 1071 857 1105
rect 891 1071 949 1105
rect 983 1071 1041 1105
rect 1075 1071 1133 1105
rect 1167 1071 1225 1105
rect 1259 1071 1288 1105
rect 0 1040 1288 1071
rect 16 731 74 737
rect 16 728 28 731
rect 14 700 28 728
rect 16 697 28 700
rect 62 728 74 731
rect 1174 731 1232 737
rect 1174 728 1186 731
rect 62 700 1186 728
rect 62 697 74 700
rect 16 691 74 697
rect 1174 697 1186 700
rect 1220 728 1232 731
rect 1220 700 1234 728
rect 1220 697 1232 700
rect 1174 691 1232 697
rect 0 561 1288 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 0 496 1288 527
rect 272 457 474 463
rect 272 456 284 457
rect 14 428 284 456
rect 272 423 284 428
rect 318 423 356 457
rect 390 423 428 457
rect 462 456 474 457
rect 462 428 1234 456
rect 462 423 474 428
rect 272 417 474 423
rect 0 17 1288 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
rect 0 -48 1288 -17
<< labels >>
rlabel comment s 0 0 0 0 4 lpflow_lsbuf_lh_hl_isowell_tap_1
flabel comment s 821 764 821 764 0 FreeSans 200 90 0 0 no_jumper_check
flabel metal1 s 66 1071 94 1105 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground bidirectional abutment
flabel metal1 s 98 700 125 728 0 FreeSans 200 0 0 0 VPB
port 3 nsew power bidirectional
flabel metal1 s 82 -11 116 23 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground bidirectional abutment
flabel metal1 s 87 428 99 456 0 FreeSans 200 0 0 0 VPWRIN
port 4 nsew power bidirectional abutment
flabel metal1 s 0 496 1248 544 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power bidirectional abutment
flabel locali s 607 268 641 302 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 1087 268 1121 302 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 1087 194 1121 228 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
rlabel locali s 1173 926 1231 1071 1 VGND
port 2 nsew ground bidirectional abutment
rlabel locali s 889 903 991 1071 1 VGND
port 2 nsew ground bidirectional abutment
rlabel locali s 715 903 753 1071 1 VGND
port 2 nsew ground bidirectional abutment
rlabel locali s 529 903 581 1071 1 VGND
port 2 nsew ground bidirectional abutment
rlabel locali s 17 926 75 1071 1 VGND
port 2 nsew ground bidirectional abutment
rlabel locali s 0 1071 1288 1105 1 VGND
port 2 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1288 48 1 VGND
port 2 nsew ground bidirectional abutment
rlabel metal1 s 0 1040 1288 1136 1 VGND
port 2 nsew ground bidirectional abutment
rlabel locali s 978 561 1024 748 1 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 978 527 1288 561 1 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 978 325 1024 527 1 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 496 1288 592 1 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 272 456 474 463 1 VPWRIN
port 4 nsew power bidirectional abutment
rlabel metal1 s 272 417 474 428 1 VPWRIN
port 4 nsew power bidirectional abutment
rlabel metal1 s 14 428 1234 456 1 VPWRIN
port 4 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1288 1088
string GDS_END 1544292
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1531050
string LEFclass CORE WELLTAP
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
