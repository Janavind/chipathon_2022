magic
tech sky130B
magscale 1 2
timestamp 1666464484
<< nwell >>
rect -38 261 498 582
<< pwell >>
rect 11 21 449 203
rect 29 -17 63 21
<< locali >>
rect 113 333 179 493
rect 281 337 347 493
rect 281 333 434 337
rect 113 299 434 333
rect 21 215 347 265
rect 381 181 434 299
rect 113 145 434 181
rect 113 51 179 145
rect 281 51 347 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 26 299 79 527
rect 213 367 247 527
rect 381 435 423 527
rect 26 17 79 109
rect 213 17 247 109
rect 381 17 431 110
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
rlabel locali s 21 215 347 265 6 A
port 1 nsew signal input
rlabel metal1 s 0 -48 460 48 8 VGND
port 2 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 3 nsew ground bidirectional
rlabel pwell s 11 21 449 203 6 VNB
port 3 nsew ground bidirectional
rlabel nwell s -38 261 498 582 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 496 460 592 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 281 51 347 145 6 Y
port 6 nsew signal output
rlabel locali s 113 51 179 145 6 Y
port 6 nsew signal output
rlabel locali s 113 145 434 181 6 Y
port 6 nsew signal output
rlabel locali s 381 181 434 299 6 Y
port 6 nsew signal output
rlabel locali s 113 299 434 333 6 Y
port 6 nsew signal output
rlabel locali s 281 333 434 337 6 Y
port 6 nsew signal output
rlabel locali s 281 337 347 493 6 Y
port 6 nsew signal output
rlabel locali s 113 333 179 493 6 Y
port 6 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 460 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2219812
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2214822
<< end >>
