magic
tech sky130A
magscale 1 2
timestamp 1666464484
<< nwell >>
rect -38 261 3074 582
<< pwell >>
rect 2398 201 3035 203
rect 1241 157 1695 201
rect 2016 157 3035 201
rect 1 21 3035 157
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 351 47 381 131
rect 423 47 453 131
rect 635 47 665 131
rect 734 47 764 131
rect 806 47 836 131
rect 901 47 931 119
rect 1011 47 1041 119
rect 1107 47 1137 131
rect 1221 47 1251 131
rect 1317 47 1347 175
rect 1401 47 1431 175
rect 1589 47 1619 175
rect 1684 47 1714 119
rect 1793 47 1823 119
rect 1888 47 1918 131
rect 1974 47 2004 131
rect 2092 47 2122 175
rect 2176 47 2206 175
rect 2379 47 2409 131
rect 2476 47 2506 177
rect 2560 47 2590 177
rect 2748 47 2778 131
rect 2843 47 2873 177
rect 2927 47 2957 177
<< scpmoshvt >>
rect 79 363 109 491
rect 163 363 193 491
rect 351 363 381 491
rect 423 363 453 491
rect 638 413 668 497
rect 722 413 752 497
rect 806 413 836 497
rect 903 413 933 497
rect 987 413 1017 497
rect 1107 413 1137 497
rect 1213 413 1243 497
rect 1321 329 1351 497
rect 1405 329 1435 497
rect 1542 329 1572 497
rect 1686 413 1716 497
rect 1770 413 1800 497
rect 1888 413 1918 497
rect 1996 413 2026 497
rect 2092 329 2122 497
rect 2164 329 2194 497
rect 2379 301 2409 429
rect 2476 297 2506 497
rect 2560 297 2590 497
rect 2748 353 2778 481
rect 2843 297 2873 497
rect 2927 297 2957 497
<< ndiff >>
rect 27 119 79 131
rect 27 85 35 119
rect 69 85 79 119
rect 27 47 79 85
rect 109 93 163 131
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 119 245 131
rect 193 85 203 119
rect 237 85 245 119
rect 193 47 245 85
rect 299 111 351 131
rect 299 77 307 111
rect 341 77 351 111
rect 299 47 351 77
rect 381 47 423 131
rect 453 103 505 131
rect 453 69 463 103
rect 497 69 505 103
rect 453 47 505 69
rect 583 111 635 131
rect 583 77 591 111
rect 625 77 635 111
rect 583 47 635 77
rect 665 89 734 131
rect 665 55 690 89
rect 724 55 734 89
rect 665 47 734 55
rect 764 47 806 131
rect 836 119 886 131
rect 1267 131 1317 175
rect 1056 119 1107 131
rect 836 111 901 119
rect 836 77 846 111
rect 880 77 901 111
rect 836 47 901 77
rect 931 93 1011 119
rect 931 59 956 93
rect 990 59 1011 93
rect 931 47 1011 59
rect 1041 47 1107 119
rect 1137 89 1221 131
rect 1137 55 1177 89
rect 1211 55 1221 89
rect 1137 47 1221 55
rect 1251 101 1317 131
rect 1251 67 1261 101
rect 1295 67 1317 101
rect 1251 47 1317 67
rect 1347 153 1401 175
rect 1347 119 1357 153
rect 1391 119 1401 153
rect 1347 47 1401 119
rect 1431 127 1483 175
rect 1431 93 1441 127
rect 1475 93 1483 127
rect 1431 47 1483 93
rect 1537 93 1589 175
rect 1537 59 1545 93
rect 1579 59 1589 93
rect 1537 47 1589 59
rect 1619 119 1669 175
rect 2042 131 2092 175
rect 1838 119 1888 131
rect 1619 47 1684 119
rect 1714 93 1793 119
rect 1714 59 1739 93
rect 1773 59 1793 93
rect 1714 47 1793 59
rect 1823 47 1888 119
rect 1918 89 1974 131
rect 1918 55 1930 89
rect 1964 55 1974 89
rect 1918 47 1974 55
rect 2004 109 2092 131
rect 2004 75 2032 109
rect 2066 75 2092 109
rect 2004 47 2092 75
rect 2122 153 2176 175
rect 2122 119 2132 153
rect 2166 119 2176 153
rect 2122 47 2176 119
rect 2206 101 2261 175
rect 2424 161 2476 177
rect 2424 131 2432 161
rect 2206 67 2216 101
rect 2250 67 2261 101
rect 2206 47 2261 67
rect 2327 103 2379 131
rect 2327 69 2335 103
rect 2369 69 2379 103
rect 2327 47 2379 69
rect 2409 127 2432 131
rect 2466 127 2476 161
rect 2409 93 2476 127
rect 2409 59 2432 93
rect 2466 59 2476 93
rect 2409 47 2476 59
rect 2506 127 2560 177
rect 2506 93 2516 127
rect 2550 93 2560 127
rect 2506 47 2560 93
rect 2590 161 2642 177
rect 2590 127 2600 161
rect 2634 127 2642 161
rect 2793 131 2843 177
rect 2590 93 2642 127
rect 2590 59 2600 93
rect 2634 59 2642 93
rect 2590 47 2642 59
rect 2696 119 2748 131
rect 2696 85 2704 119
rect 2738 85 2748 119
rect 2696 47 2748 85
rect 2778 93 2843 131
rect 2778 59 2799 93
rect 2833 59 2843 93
rect 2778 47 2843 59
rect 2873 129 2927 177
rect 2873 95 2883 129
rect 2917 95 2927 129
rect 2873 47 2927 95
rect 2957 161 3009 177
rect 2957 127 2967 161
rect 3001 127 3009 161
rect 2957 93 3009 127
rect 2957 59 2967 93
rect 3001 59 3009 93
rect 2957 47 3009 59
<< pdiff >>
rect 27 477 79 491
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 363 79 375
rect 109 461 163 491
rect 109 427 119 461
rect 153 427 163 461
rect 109 363 163 427
rect 193 477 245 491
rect 193 443 203 477
rect 237 443 245 477
rect 193 409 245 443
rect 193 375 203 409
rect 237 375 245 409
rect 193 363 245 375
rect 299 479 351 491
rect 299 445 307 479
rect 341 445 351 479
rect 299 411 351 445
rect 299 377 307 411
rect 341 377 351 411
rect 299 363 351 377
rect 381 363 423 491
rect 453 477 505 491
rect 453 443 463 477
rect 497 443 505 477
rect 453 409 505 443
rect 571 477 638 497
rect 571 443 579 477
rect 613 443 638 477
rect 571 413 638 443
rect 668 477 722 497
rect 668 443 678 477
rect 712 443 722 477
rect 668 413 722 443
rect 752 413 806 497
rect 836 477 903 497
rect 836 443 846 477
rect 880 443 903 477
rect 836 413 903 443
rect 933 484 987 497
rect 933 450 943 484
rect 977 450 987 484
rect 933 413 987 450
rect 1017 413 1107 497
rect 1137 475 1213 497
rect 1137 441 1157 475
rect 1191 441 1213 475
rect 1137 413 1213 441
rect 1243 459 1321 497
rect 1243 425 1277 459
rect 1311 425 1321 459
rect 1243 413 1321 425
rect 453 375 463 409
rect 497 375 505 409
rect 453 363 505 375
rect 1259 391 1321 413
rect 1259 357 1277 391
rect 1311 357 1321 391
rect 1259 329 1321 357
rect 1351 329 1405 497
rect 1435 485 1542 497
rect 1435 451 1451 485
rect 1485 451 1542 485
rect 1435 417 1542 451
rect 1435 383 1451 417
rect 1485 383 1542 417
rect 1435 329 1542 383
rect 1572 413 1686 497
rect 1716 484 1770 497
rect 1716 450 1726 484
rect 1760 450 1770 484
rect 1716 413 1770 450
rect 1800 413 1888 497
rect 1918 485 1996 497
rect 1918 451 1940 485
rect 1974 451 1996 485
rect 1918 413 1996 451
rect 2026 459 2092 497
rect 2026 425 2048 459
rect 2082 425 2092 459
rect 2026 413 2092 425
rect 1572 329 1624 413
rect 2041 329 2092 413
rect 2122 329 2164 497
rect 2194 485 2246 497
rect 2194 451 2204 485
rect 2238 451 2246 485
rect 2424 485 2476 497
rect 2194 329 2246 451
rect 2424 451 2432 485
rect 2466 451 2476 485
rect 2424 429 2476 451
rect 2327 349 2379 429
rect 2327 315 2335 349
rect 2369 315 2379 349
rect 2327 301 2379 315
rect 2409 301 2476 429
rect 2424 297 2476 301
rect 2506 448 2560 497
rect 2506 414 2516 448
rect 2550 414 2560 448
rect 2506 380 2560 414
rect 2506 346 2516 380
rect 2550 346 2560 380
rect 2506 297 2560 346
rect 2590 485 2642 497
rect 2590 451 2600 485
rect 2634 451 2642 485
rect 2793 481 2843 497
rect 2590 417 2642 451
rect 2590 383 2600 417
rect 2634 383 2642 417
rect 2590 349 2642 383
rect 2696 467 2748 481
rect 2696 433 2704 467
rect 2738 433 2748 467
rect 2696 399 2748 433
rect 2696 365 2704 399
rect 2738 365 2748 399
rect 2696 353 2748 365
rect 2778 473 2843 481
rect 2778 439 2799 473
rect 2833 439 2843 473
rect 2778 405 2843 439
rect 2778 371 2799 405
rect 2833 371 2843 405
rect 2778 353 2843 371
rect 2590 315 2600 349
rect 2634 315 2642 349
rect 2590 297 2642 315
rect 2793 297 2843 353
rect 2873 449 2927 497
rect 2873 415 2883 449
rect 2917 415 2927 449
rect 2873 381 2927 415
rect 2873 347 2883 381
rect 2917 347 2927 381
rect 2873 297 2927 347
rect 2957 485 3009 497
rect 2957 451 2967 485
rect 3001 451 3009 485
rect 2957 417 3009 451
rect 2957 383 2967 417
rect 3001 383 3009 417
rect 2957 349 3009 383
rect 2957 315 2967 349
rect 3001 315 3009 349
rect 2957 297 3009 315
<< ndiffc >>
rect 35 85 69 119
rect 119 59 153 93
rect 203 85 237 119
rect 307 77 341 111
rect 463 69 497 103
rect 591 77 625 111
rect 690 55 724 89
rect 846 77 880 111
rect 956 59 990 93
rect 1177 55 1211 89
rect 1261 67 1295 101
rect 1357 119 1391 153
rect 1441 93 1475 127
rect 1545 59 1579 93
rect 1739 59 1773 93
rect 1930 55 1964 89
rect 2032 75 2066 109
rect 2132 119 2166 153
rect 2216 67 2250 101
rect 2335 69 2369 103
rect 2432 127 2466 161
rect 2432 59 2466 93
rect 2516 93 2550 127
rect 2600 127 2634 161
rect 2600 59 2634 93
rect 2704 85 2738 119
rect 2799 59 2833 93
rect 2883 95 2917 129
rect 2967 127 3001 161
rect 2967 59 3001 93
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 119 427 153 461
rect 203 443 237 477
rect 203 375 237 409
rect 307 445 341 479
rect 307 377 341 411
rect 463 443 497 477
rect 579 443 613 477
rect 678 443 712 477
rect 846 443 880 477
rect 943 450 977 484
rect 1157 441 1191 475
rect 1277 425 1311 459
rect 463 375 497 409
rect 1277 357 1311 391
rect 1451 451 1485 485
rect 1451 383 1485 417
rect 1726 450 1760 484
rect 1940 451 1974 485
rect 2048 425 2082 459
rect 2204 451 2238 485
rect 2432 451 2466 485
rect 2335 315 2369 349
rect 2516 414 2550 448
rect 2516 346 2550 380
rect 2600 451 2634 485
rect 2600 383 2634 417
rect 2704 433 2738 467
rect 2704 365 2738 399
rect 2799 439 2833 473
rect 2799 371 2833 405
rect 2600 315 2634 349
rect 2883 415 2917 449
rect 2883 347 2917 381
rect 2967 451 3001 485
rect 2967 383 3001 417
rect 2967 315 3001 349
<< poly >>
rect 79 491 109 517
rect 163 491 193 517
rect 351 491 381 517
rect 423 491 453 517
rect 638 497 668 523
rect 722 497 752 523
rect 806 497 836 523
rect 903 497 933 523
rect 987 497 1017 523
rect 1107 497 1137 523
rect 1213 497 1243 523
rect 1321 497 1351 523
rect 1405 497 1435 523
rect 1542 497 1572 523
rect 1686 497 1716 523
rect 1770 497 1800 523
rect 1888 497 1918 523
rect 1996 497 2026 523
rect 2092 497 2122 523
rect 2164 497 2194 523
rect 2476 497 2506 523
rect 2560 497 2590 523
rect 638 397 668 413
rect 722 397 752 413
rect 539 365 596 381
rect 79 348 109 363
rect 45 318 109 348
rect 45 280 75 318
rect 21 264 75 280
rect 163 274 193 363
rect 351 331 381 363
rect 21 230 31 264
rect 65 230 75 264
rect 21 214 75 230
rect 117 264 193 274
rect 295 315 381 331
rect 423 345 453 363
rect 539 345 552 365
rect 423 331 552 345
rect 586 331 596 365
rect 423 315 596 331
rect 638 367 752 397
rect 295 281 305 315
rect 339 281 381 315
rect 295 265 381 281
rect 117 230 133 264
rect 167 230 193 264
rect 117 220 193 230
rect 45 176 75 214
rect 45 146 109 176
rect 79 131 109 146
rect 163 131 193 220
rect 351 131 381 265
rect 423 203 483 219
rect 423 169 433 203
rect 467 177 483 203
rect 638 177 668 367
rect 806 325 836 413
rect 755 315 836 325
rect 755 281 771 315
rect 805 281 836 315
rect 755 271 836 281
rect 467 169 668 177
rect 423 147 668 169
rect 710 203 764 219
rect 710 169 720 203
rect 754 169 764 203
rect 710 153 764 169
rect 423 131 453 147
rect 635 131 665 147
rect 734 131 764 153
rect 806 131 836 271
rect 903 279 933 413
rect 987 375 1017 413
rect 1107 381 1137 413
rect 975 365 1041 375
rect 975 331 991 365
rect 1025 331 1041 365
rect 975 321 1041 331
rect 1107 365 1171 381
rect 1107 331 1127 365
rect 1161 331 1171 365
rect 1107 315 1171 331
rect 903 249 1041 279
rect 1011 219 1041 249
rect 901 191 969 207
rect 901 157 925 191
rect 959 157 969 191
rect 901 141 969 157
rect 1011 203 1065 219
rect 1011 169 1021 203
rect 1055 169 1065 203
rect 1011 153 1065 169
rect 901 119 931 141
rect 1011 119 1041 153
rect 1107 131 1137 315
rect 1213 229 1243 413
rect 1686 381 1716 413
rect 1662 365 1716 381
rect 1770 375 1800 413
rect 1888 381 1918 413
rect 1662 331 1672 365
rect 1706 331 1716 365
rect 1321 297 1351 329
rect 1285 281 1351 297
rect 1285 247 1295 281
rect 1329 247 1351 281
rect 1285 231 1351 247
rect 1405 297 1435 329
rect 1405 281 1491 297
rect 1405 247 1447 281
rect 1481 247 1491 281
rect 1405 231 1491 247
rect 1542 263 1572 329
rect 1662 315 1716 331
rect 1758 365 1824 375
rect 1758 331 1774 365
rect 1808 331 1824 365
rect 1758 321 1824 331
rect 1888 365 1954 381
rect 1888 331 1910 365
rect 1944 331 1954 365
rect 1686 279 1716 315
rect 1888 315 1954 331
rect 1542 247 1619 263
rect 1686 249 1823 279
rect 1542 233 1575 247
rect 1183 213 1243 229
rect 1183 179 1193 213
rect 1227 193 1243 213
rect 1227 179 1251 193
rect 1183 163 1251 179
rect 1317 175 1347 231
rect 1405 220 1435 231
rect 1401 190 1435 220
rect 1565 213 1575 233
rect 1609 213 1619 247
rect 1565 197 1619 213
rect 1401 175 1431 190
rect 1589 175 1619 197
rect 1684 191 1751 207
rect 1221 131 1251 163
rect 1684 157 1707 191
rect 1741 157 1751 191
rect 1684 141 1751 157
rect 1684 119 1714 141
rect 1793 119 1823 249
rect 1888 131 1918 315
rect 1996 229 2026 413
rect 2379 429 2409 455
rect 2092 281 2122 329
rect 1960 213 2026 229
rect 2068 265 2122 281
rect 2164 297 2194 329
rect 2164 281 2260 297
rect 2164 267 2216 281
rect 2068 231 2078 265
rect 2112 231 2122 265
rect 2068 215 2122 231
rect 1960 179 1970 213
rect 2004 179 2026 213
rect 1960 163 2026 179
rect 2092 175 2122 215
rect 2176 247 2216 267
rect 2250 247 2260 281
rect 2379 269 2409 301
rect 2748 481 2778 507
rect 2843 497 2873 523
rect 2927 497 2957 523
rect 2748 337 2778 353
rect 2722 307 2778 337
rect 2176 231 2260 247
rect 2324 253 2409 269
rect 2476 265 2506 297
rect 2176 175 2206 231
rect 2324 219 2334 253
rect 2368 219 2409 253
rect 2324 203 2409 219
rect 1974 131 2004 163
rect 2379 131 2409 203
rect 2452 259 2506 265
rect 2560 259 2590 297
rect 2722 259 2752 307
rect 2843 265 2873 297
rect 2927 265 2957 297
rect 2452 249 2752 259
rect 2452 215 2462 249
rect 2496 215 2752 249
rect 2452 205 2752 215
rect 2452 199 2506 205
rect 2476 177 2506 199
rect 2560 177 2590 205
rect 2722 176 2752 205
rect 2814 249 2957 265
rect 2814 215 2824 249
rect 2858 215 2957 249
rect 2814 199 2957 215
rect 2843 177 2873 199
rect 2927 177 2957 199
rect 2722 146 2778 176
rect 2748 131 2778 146
rect 79 21 109 47
rect 163 21 193 47
rect 351 21 381 47
rect 423 21 453 47
rect 635 21 665 47
rect 734 21 764 47
rect 806 21 836 47
rect 901 21 931 47
rect 1011 21 1041 47
rect 1107 21 1137 47
rect 1221 21 1251 47
rect 1317 21 1347 47
rect 1401 21 1431 47
rect 1589 21 1619 47
rect 1684 21 1714 47
rect 1793 21 1823 47
rect 1888 21 1918 47
rect 1974 21 2004 47
rect 2092 21 2122 47
rect 2176 21 2206 47
rect 2379 21 2409 47
rect 2476 21 2506 47
rect 2560 21 2590 47
rect 2748 21 2778 47
rect 2843 21 2873 47
rect 2927 21 2957 47
<< polycont >>
rect 31 230 65 264
rect 552 331 586 365
rect 305 281 339 315
rect 133 230 167 264
rect 433 169 467 203
rect 771 281 805 315
rect 720 169 754 203
rect 991 331 1025 365
rect 1127 331 1161 365
rect 925 157 959 191
rect 1021 169 1055 203
rect 1672 331 1706 365
rect 1295 247 1329 281
rect 1447 247 1481 281
rect 1774 331 1808 365
rect 1910 331 1944 365
rect 1193 179 1227 213
rect 1575 213 1609 247
rect 1707 157 1741 191
rect 2078 231 2112 265
rect 1970 179 2004 213
rect 2216 247 2250 281
rect 2334 219 2368 253
rect 2462 215 2496 249
rect 2824 215 2858 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3036 561
rect 34 477 69 493
rect 34 443 35 477
rect 34 409 69 443
rect 103 461 169 527
rect 103 427 119 461
rect 153 427 169 461
rect 203 477 247 493
rect 237 443 247 477
rect 34 375 35 409
rect 203 409 247 443
rect 69 375 167 393
rect 34 359 167 375
rect 17 264 87 325
rect 17 230 31 264
rect 65 230 87 264
rect 17 195 87 230
rect 121 264 167 359
rect 121 230 133 264
rect 121 187 167 230
rect 34 153 121 161
rect 155 153 167 187
rect 34 127 167 153
rect 237 391 247 409
rect 286 479 357 527
rect 286 445 307 479
rect 341 445 357 479
rect 579 477 613 493
rect 286 411 357 445
rect 286 377 307 411
rect 341 377 357 411
rect 443 443 463 477
rect 497 443 515 477
rect 443 409 515 443
rect 443 375 463 409
rect 497 375 515 409
rect 659 477 728 527
rect 659 443 678 477
rect 712 443 728 477
rect 846 477 891 493
rect 579 381 613 443
rect 203 357 213 375
rect 34 119 69 127
rect 34 85 35 119
rect 203 119 247 357
rect 283 315 339 337
rect 283 281 305 315
rect 283 205 339 281
rect 387 219 431 339
rect 481 281 515 375
rect 549 365 613 381
rect 549 331 552 365
rect 586 349 613 365
rect 586 331 729 349
rect 549 315 729 331
rect 481 255 615 281
rect 481 250 581 255
rect 487 247 581 250
rect 512 221 581 247
rect 387 203 467 219
rect 387 169 433 203
rect 387 153 467 169
rect 512 215 615 221
rect 695 219 729 315
rect 765 315 805 475
rect 765 281 771 315
rect 765 265 805 281
rect 880 443 891 477
rect 927 450 943 484
rect 977 450 1093 484
rect 846 255 891 443
rect 846 221 857 255
rect 34 69 69 85
rect 103 59 119 93
rect 153 59 169 93
rect 237 85 247 119
rect 203 69 247 85
rect 286 111 341 127
rect 286 77 307 111
rect 103 17 169 59
rect 286 17 341 77
rect 387 69 429 153
rect 512 119 546 215
rect 695 203 754 219
rect 695 169 720 203
rect 695 159 754 169
rect 463 103 546 119
rect 497 69 546 103
rect 463 53 546 69
rect 591 153 754 159
rect 591 125 729 153
rect 591 111 625 125
rect 846 111 891 221
rect 925 357 949 391
rect 983 365 1025 391
rect 983 357 991 365
rect 925 331 991 357
rect 925 315 1025 331
rect 925 191 969 315
rect 1059 281 1093 450
rect 1141 475 1217 527
rect 1435 485 1501 527
rect 1141 441 1157 475
rect 1191 441 1217 475
rect 1277 459 1311 475
rect 1277 407 1311 425
rect 1435 451 1451 485
rect 1485 451 1501 485
rect 1924 485 2000 527
rect 1435 417 1501 451
rect 1710 450 1726 484
rect 1760 450 1876 484
rect 1924 451 1940 485
rect 1974 451 2000 485
rect 2188 485 2482 527
rect 2048 459 2082 475
rect 1127 391 1397 407
rect 1127 365 1277 391
rect 1161 357 1277 365
rect 1311 357 1397 391
rect 1435 383 1451 417
rect 1485 383 1501 417
rect 1672 391 1719 397
rect 1161 331 1177 357
rect 1127 315 1177 331
rect 1279 281 1329 297
rect 1059 247 1295 281
rect 1059 239 1143 247
rect 959 157 969 191
rect 925 141 969 157
rect 1005 169 1021 203
rect 1055 187 1075 203
rect 1005 153 1041 169
rect 1005 129 1075 153
rect 591 61 625 77
rect 674 55 690 89
rect 724 55 740 89
rect 880 77 891 111
rect 1109 93 1143 239
rect 1285 231 1329 247
rect 1363 213 1397 357
rect 1672 365 1685 391
rect 1706 331 1719 357
rect 1431 323 1632 331
rect 1431 289 1593 323
rect 1627 289 1632 323
rect 1672 315 1719 331
rect 1767 365 1808 381
rect 1767 331 1774 365
rect 1431 283 1632 289
rect 1431 281 1497 283
rect 1431 247 1447 281
rect 1481 247 1497 281
rect 1767 261 1808 331
rect 1684 255 1808 261
rect 1559 213 1575 247
rect 1609 213 1625 247
rect 1177 179 1193 213
rect 1227 193 1243 213
rect 1227 187 1259 193
rect 1177 153 1225 179
rect 1363 179 1625 213
rect 1684 221 1685 255
rect 1719 225 1808 255
rect 1842 281 1876 450
rect 2188 451 2204 485
rect 2238 451 2432 485
rect 2466 451 2482 485
rect 2048 417 2082 425
rect 2516 448 2566 493
rect 1910 383 2482 417
rect 1910 365 1960 383
rect 1944 331 1960 365
rect 1910 315 1960 331
rect 1842 265 2112 281
rect 1842 247 2078 265
rect 1719 221 1741 225
rect 1684 191 1741 221
rect 1363 153 1407 179
rect 1177 147 1259 153
rect 1341 119 1357 153
rect 1391 119 1407 153
rect 1684 157 1707 191
rect 1441 127 1475 143
rect 1684 141 1741 157
rect 846 61 891 77
rect 674 17 740 55
rect 940 59 956 93
rect 990 59 1143 93
rect 940 53 1143 59
rect 1177 89 1211 105
rect 1177 17 1211 55
rect 1245 67 1261 101
rect 1295 85 1311 101
rect 1842 93 1876 247
rect 2068 231 2078 247
rect 2068 215 2112 231
rect 1951 187 1970 213
rect 1951 153 1961 187
rect 2004 179 2026 213
rect 1995 153 2026 179
rect 2146 156 2182 383
rect 1951 147 2026 153
rect 2116 153 2182 156
rect 2116 119 2132 153
rect 2166 119 2182 153
rect 2216 323 2335 349
rect 2216 289 2237 323
rect 2271 315 2335 323
rect 2369 315 2385 349
rect 2216 281 2271 289
rect 2250 247 2271 281
rect 2448 265 2482 383
rect 2550 414 2566 448
rect 2516 380 2566 414
rect 2550 346 2566 380
rect 2516 326 2566 346
rect 2216 185 2271 247
rect 2318 253 2414 265
rect 2318 219 2334 253
rect 2368 219 2414 253
rect 2448 249 2496 265
rect 2448 215 2462 249
rect 2448 199 2496 215
rect 2216 151 2369 185
rect 1441 85 1475 93
rect 1295 67 1475 85
rect 1245 51 1475 67
rect 1529 59 1545 93
rect 1579 59 1595 93
rect 1529 17 1595 59
rect 1723 59 1739 93
rect 1773 59 1876 93
rect 1723 53 1876 59
rect 1912 89 1964 105
rect 1912 55 1930 89
rect 1912 17 1964 55
rect 2016 75 2032 109
rect 2066 85 2082 109
rect 2216 101 2250 117
rect 2066 75 2216 85
rect 2016 67 2216 75
rect 2016 51 2250 67
rect 2324 103 2369 151
rect 2324 69 2335 103
rect 2324 53 2369 69
rect 2416 127 2432 161
rect 2466 127 2482 161
rect 2532 143 2566 326
rect 2600 485 2647 527
rect 2634 451 2647 485
rect 2600 417 2647 451
rect 2634 383 2647 417
rect 2600 349 2647 383
rect 2634 315 2647 349
rect 2600 299 2647 315
rect 2691 467 2754 483
rect 2691 433 2704 467
rect 2738 433 2754 467
rect 2691 399 2754 433
rect 2691 365 2704 399
rect 2738 365 2754 399
rect 2691 265 2754 365
rect 2790 473 2849 527
rect 2790 439 2799 473
rect 2833 439 2849 473
rect 2790 405 2849 439
rect 2790 371 2799 405
rect 2833 371 2849 405
rect 2790 353 2849 371
rect 2883 449 2933 493
rect 2917 415 2933 449
rect 2883 381 2933 415
rect 2917 347 2933 381
rect 2883 289 2933 347
rect 2967 485 3015 527
rect 3001 451 3015 485
rect 2967 417 3015 451
rect 3001 383 3015 417
rect 2967 349 3015 383
rect 3001 315 3015 349
rect 2967 299 3015 315
rect 2691 249 2858 265
rect 2691 215 2824 249
rect 2691 199 2858 215
rect 2416 93 2482 127
rect 2416 59 2432 93
rect 2466 59 2482 93
rect 2416 17 2482 59
rect 2516 127 2566 143
rect 2550 93 2566 127
rect 2516 51 2566 93
rect 2600 161 2647 177
rect 2634 127 2647 161
rect 2600 93 2647 127
rect 2634 59 2647 93
rect 2600 17 2647 59
rect 2691 119 2754 199
rect 2892 165 2933 289
rect 2691 85 2704 119
rect 2738 85 2754 119
rect 2883 129 2933 165
rect 2691 51 2754 85
rect 2790 93 2849 109
rect 2790 59 2799 93
rect 2833 59 2849 93
rect 2790 17 2849 59
rect 2917 95 2933 129
rect 2883 51 2933 95
rect 2967 161 3015 177
rect 3001 127 3015 161
rect 2967 93 3015 127
rect 3001 59 3015 93
rect 2967 17 3015 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3036 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 2605 527 2639 561
rect 2697 527 2731 561
rect 2789 527 2823 561
rect 2881 527 2915 561
rect 2973 527 3007 561
rect 121 153 155 187
rect 213 375 237 391
rect 237 375 247 391
rect 213 357 247 375
rect 581 221 615 255
rect 857 221 891 255
rect 949 357 983 391
rect 1041 169 1055 187
rect 1055 169 1075 187
rect 1041 153 1075 169
rect 1685 365 1719 391
rect 1685 357 1706 365
rect 1706 357 1719 365
rect 1593 289 1627 323
rect 1225 179 1227 187
rect 1227 179 1259 187
rect 1225 153 1259 179
rect 1685 221 1719 255
rect 1961 179 1970 187
rect 1970 179 1995 187
rect 1961 153 1995 179
rect 2237 289 2271 323
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
rect 2697 -17 2731 17
rect 2789 -17 2823 17
rect 2881 -17 2915 17
rect 2973 -17 3007 17
<< metal1 >>
rect 0 561 3036 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3036 561
rect 0 496 3036 527
rect 201 391 259 397
rect 201 357 213 391
rect 247 388 259 391
rect 937 391 995 397
rect 937 388 949 391
rect 247 360 949 388
rect 247 357 259 360
rect 201 351 259 357
rect 937 357 949 360
rect 983 388 995 391
rect 1673 391 1731 397
rect 1673 388 1685 391
rect 983 360 1685 388
rect 983 357 995 360
rect 937 351 995 357
rect 1673 357 1685 360
rect 1719 357 1731 391
rect 1673 351 1731 357
rect 1581 323 1639 329
rect 1581 289 1593 323
rect 1627 320 1639 323
rect 2225 323 2283 329
rect 2225 320 2237 323
rect 1627 292 2237 320
rect 1627 289 1639 292
rect 1581 283 1639 289
rect 2225 289 2237 292
rect 2271 289 2283 323
rect 2225 283 2283 289
rect 569 255 627 261
rect 569 221 581 255
rect 615 252 627 255
rect 845 255 903 261
rect 845 252 857 255
rect 615 224 857 252
rect 615 221 627 224
rect 569 215 627 221
rect 845 221 857 224
rect 891 221 903 255
rect 1673 255 1731 261
rect 1673 252 1685 255
rect 845 215 903 221
rect 1044 224 1685 252
rect 1044 193 1087 224
rect 1673 221 1685 224
rect 1719 221 1731 255
rect 1673 215 1731 221
rect 109 187 167 193
rect 109 153 121 187
rect 155 184 167 187
rect 1029 187 1087 193
rect 1029 184 1041 187
rect 155 156 1041 184
rect 155 153 167 156
rect 109 147 167 153
rect 1029 153 1041 156
rect 1075 153 1087 187
rect 1029 147 1087 153
rect 1213 187 1271 193
rect 1213 153 1225 187
rect 1259 184 1271 187
rect 1949 187 2007 193
rect 1949 184 1961 187
rect 1259 156 1961 184
rect 1259 153 1271 156
rect 1213 147 1271 153
rect 1949 153 1961 156
rect 1995 153 2007 187
rect 1949 147 2007 153
rect 0 17 3036 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3036 17
rect 0 -48 3036 -17
<< labels >>
flabel locali s 305 289 339 323 0 FreeSans 400 0 0 0 SCD
port 4 nsew signal input
flabel locali s 305 221 339 255 0 FreeSans 400 0 0 0 SCD
port 4 nsew signal input
flabel locali s 397 289 431 323 0 FreeSans 400 0 0 0 SCE
port 5 nsew signal input
flabel locali s 397 221 431 255 0 FreeSans 400 0 0 0 SCE
port 5 nsew signal input
flabel locali s 395 85 429 119 0 FreeSans 400 0 0 0 SCE
port 5 nsew signal input
flabel locali s 2340 221 2374 255 0 FreeSans 400 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 29 -17 63 17 3 FreeSans 400 0 0 0 VGND
port 7 nsew ground bidirectional abutment
flabel locali s 29 221 63 255 0 FreeSans 400 0 0 0 CLK_N
port 1 nsew clock input
flabel locali s 29 289 63 323 0 FreeSans 400 0 0 0 CLK_N
port 1 nsew clock input
flabel locali s 1225 153 1259 187 0 FreeSans 400 0 0 0 SET_B
port 6 nsew signal input
flabel locali s 2888 85 2922 119 0 FreeSans 400 0 0 0 Q
port 11 nsew signal output
flabel locali s 2888 357 2922 391 0 FreeSans 400 0 0 0 Q
port 11 nsew signal output
flabel locali s 2888 425 2922 459 0 FreeSans 400 0 0 0 Q
port 11 nsew signal output
flabel locali s 29 527 63 561 3 FreeSans 400 0 0 0 VPWR
port 10 nsew power bidirectional abutment
flabel locali s 765 289 799 323 0 FreeSans 200 0 0 0 D
port 2 nsew signal input
flabel locali s 765 425 799 459 0 FreeSans 200 0 0 0 D
port 2 nsew signal input
flabel locali s 2524 425 2558 459 0 FreeSans 400 0 0 0 Q_N
port 12 nsew signal output
flabel locali s 2524 357 2558 391 0 FreeSans 400 0 0 0 Q_N
port 12 nsew signal output
flabel locali s 2524 85 2558 119 0 FreeSans 400 0 0 0 Q_N
port 12 nsew signal output
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 7 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 10 nsew power bidirectional abutment
flabel nwell s 29 527 63 561 3 FreeSans 400 0 0 0 VPB
port 9 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
port 9 nsew
flabel pwell s 29 -17 63 17 3 FreeSans 400 0 0 0 VNB
port 8 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
port 8 nsew
rlabel comment s 0 0 0 0 4 sdfbbn_2
rlabel locali s 1951 147 2026 213 1 SET_B
port 6 nsew signal input
rlabel metal1 s 1949 184 2007 193 1 SET_B
port 6 nsew signal input
rlabel metal1 s 1949 147 2007 156 1 SET_B
port 6 nsew signal input
rlabel metal1 s 1213 184 1271 193 1 SET_B
port 6 nsew signal input
rlabel metal1 s 1213 156 2007 184 1 SET_B
port 6 nsew signal input
rlabel metal1 s 1213 147 1271 156 1 SET_B
port 6 nsew signal input
rlabel metal1 s 0 -48 3036 48 1 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 496 3036 592 1 VPWR
port 10 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3036 544
string GDS_END 218634
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 195260
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
