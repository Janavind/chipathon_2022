magic
tech sky130A
magscale 1 2
timestamp 1666199351
<< nwell >>
rect -38 261 1050 582
<< pwell >>
rect 1 21 964 157
rect 29 -17 63 21
<< locali >>
rect 284 347 336 492
rect 456 347 508 492
rect 628 347 680 492
rect 800 347 852 492
rect 284 299 946 347
rect 17 143 80 265
rect 752 181 946 299
rect 284 147 946 181
rect 284 56 336 147
rect 456 56 508 147
rect 628 56 680 147
rect 800 56 852 147
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 19 305 78 527
rect 114 265 164 492
rect 198 305 250 527
rect 370 381 422 527
rect 542 381 594 527
rect 714 381 766 527
rect 886 381 945 527
rect 114 215 718 265
rect 29 17 78 109
rect 114 53 164 215
rect 198 17 250 122
rect 370 17 422 113
rect 542 17 594 113
rect 714 17 766 113
rect 886 17 946 113
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
<< metal1 >>
rect 0 561 1012 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 0 496 1012 527
rect 0 17 1012 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
rect 0 -48 1012 -17
<< labels >>
rlabel locali s 17 143 80 265 6 A
port 1 nsew signal input
rlabel metal1 s 0 -48 1012 48 8 VGND
port 2 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 3 nsew ground bidirectional
rlabel pwell s 1 21 964 157 6 VNB
port 3 nsew ground bidirectional
rlabel nwell s -38 261 1050 582 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 496 1012 592 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 800 56 852 147 6 X
port 6 nsew signal output
rlabel locali s 628 56 680 147 6 X
port 6 nsew signal output
rlabel locali s 456 56 508 147 6 X
port 6 nsew signal output
rlabel locali s 284 56 336 147 6 X
port 6 nsew signal output
rlabel locali s 284 147 946 181 6 X
port 6 nsew signal output
rlabel locali s 752 181 946 299 6 X
port 6 nsew signal output
rlabel locali s 284 299 946 347 6 X
port 6 nsew signal output
rlabel locali s 800 347 852 492 6 X
port 6 nsew signal output
rlabel locali s 628 347 680 492 6 X
port 6 nsew signal output
rlabel locali s 456 347 508 492 6 X
port 6 nsew signal output
rlabel locali s 284 347 336 492 6 X
port 6 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1012 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3189440
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3181698
<< end >>
